VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_openram_wrapper
  CLASS BLOCK ;
  FOREIGN wb_openram_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 300.000 ;
  PIN ram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END ram_addr0[0]
  PIN ram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END ram_addr0[1]
  PIN ram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END ram_addr0[2]
  PIN ram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END ram_addr0[3]
  PIN ram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 293.800 40.000 294.400 ;
    END
  END ram_addr0[4]
  PIN ram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 296.000 39.010 300.000 ;
    END
  END ram_addr0[5]
  PIN ram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END ram_addr0[6]
  PIN ram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 25.880 40.000 26.480 ;
    END
  END ram_addr0[7]
  PIN ram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 296.000 15.090 300.000 ;
    END
  END ram_clk0
  PIN ram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 55.800 40.000 56.400 ;
    END
  END ram_csb0
  PIN ram_din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END ram_din0[0]
  PIN ram_din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 84.360 40.000 84.960 ;
    END
  END ram_din0[10]
  PIN ram_din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END ram_din0[11]
  PIN ram_din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 224.440 40.000 225.040 ;
    END
  END ram_din0[12]
  PIN ram_din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END ram_din0[13]
  PIN ram_din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END ram_din0[14]
  PIN ram_din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END ram_din0[15]
  PIN ram_din0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END ram_din0[16]
  PIN ram_din0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 296.000 28.890 300.000 ;
    END
  END ram_din0[17]
  PIN ram_din0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END ram_din0[18]
  PIN ram_din0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 239.400 40.000 240.000 ;
    END
  END ram_din0[19]
  PIN ram_din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END ram_din0[1]
  PIN ram_din0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 145.560 40.000 146.160 ;
    END
  END ram_din0[20]
  PIN ram_din0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END ram_din0[21]
  PIN ram_din0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 165.960 40.000 166.560 ;
    END
  END ram_din0[22]
  PIN ram_din0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 28.600 40.000 29.200 ;
    END
  END ram_din0[23]
  PIN ram_din0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END ram_din0[24]
  PIN ram_din0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 285.640 40.000 286.240 ;
    END
  END ram_din0[25]
  PIN ram_din0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END ram_din0[26]
  PIN ram_din0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END ram_din0[27]
  PIN ram_din0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 270.680 40.000 271.280 ;
    END
  END ram_din0[28]
  PIN ram_din0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 114.280 40.000 114.880 ;
    END
  END ram_din0[29]
  PIN ram_din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 111.560 40.000 112.160 ;
    END
  END ram_din0[2]
  PIN ram_din0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END ram_din0[30]
  PIN ram_din0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END ram_din0[31]
  PIN ram_din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END ram_din0[3]
  PIN ram_din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END ram_din0[4]
  PIN ram_din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 141.480 40.000 142.080 ;
    END
  END ram_din0[5]
  PIN ram_din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END ram_din0[6]
  PIN ram_din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 172.760 40.000 173.360 ;
    END
  END ram_din0[7]
  PIN ram_din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 296.000 12.330 300.000 ;
    END
  END ram_din0[8]
  PIN ram_din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 296.000 10.490 300.000 ;
    END
  END ram_din0[9]
  PIN ram_dout0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 278.840 40.000 279.440 ;
    END
  END ram_dout0[0]
  PIN ram_dout0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 296.000 36.250 300.000 ;
    END
  END ram_dout0[10]
  PIN ram_dout0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END ram_dout0[11]
  PIN ram_dout0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END ram_dout0[12]
  PIN ram_dout0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 251.640 40.000 252.240 ;
    END
  END ram_dout0[13]
  PIN ram_dout0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END ram_dout0[14]
  PIN ram_dout0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 204.040 40.000 204.640 ;
    END
  END ram_dout0[15]
  PIN ram_dout0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END ram_dout0[16]
  PIN ram_dout0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 95.240 40.000 95.840 ;
    END
  END ram_dout0[17]
  PIN ram_dout0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END ram_dout0[18]
  PIN ram_dout0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END ram_dout0[19]
  PIN ram_dout0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END ram_dout0[1]
  PIN ram_dout0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 53.080 40.000 53.680 ;
    END
  END ram_dout0[20]
  PIN ram_dout0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 176.840 40.000 177.440 ;
    END
  END ram_dout0[21]
  PIN ram_dout0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 274.760 40.000 275.360 ;
    END
  END ram_dout0[22]
  PIN ram_dout0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END ram_dout0[23]
  PIN ram_dout0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 197.240 40.000 197.840 ;
    END
  END ram_dout0[24]
  PIN ram_dout0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 76.200 40.000 76.800 ;
    END
  END ram_dout0[25]
  PIN ram_dout0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END ram_dout0[26]
  PIN ram_dout0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END ram_dout0[27]
  PIN ram_dout0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END ram_dout0[28]
  PIN ram_dout0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 296.000 26.130 300.000 ;
    END
  END ram_dout0[29]
  PIN ram_dout0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 296.000 30.730 300.000 ;
    END
  END ram_dout0[2]
  PIN ram_dout0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END ram_dout0[30]
  PIN ram_dout0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 21.800 40.000 22.400 ;
    END
  END ram_dout0[31]
  PIN ram_dout0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END ram_dout0[3]
  PIN ram_dout0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 296.000 20.610 300.000 ;
    END
  END ram_dout0[4]
  PIN ram_dout0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 255.720 40.000 256.320 ;
    END
  END ram_dout0[5]
  PIN ram_dout0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END ram_dout0[6]
  PIN ram_dout0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END ram_dout0[7]
  PIN ram_dout0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END ram_dout0[8]
  PIN ram_dout0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END ram_dout0[9]
  PIN ram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END ram_web0
  PIN ram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 153.720 40.000 154.320 ;
    END
  END ram_wmask0[0]
  PIN ram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END ram_wmask0[1]
  PIN ram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END ram_wmask0[2]
  PIN ram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 262.520 40.000 263.120 ;
    END
  END ram_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.545 10.640 11.145 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.195 10.640 20.795 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.850 10.640 30.450 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.370 10.640 15.970 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.025 10.640 25.625 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 59.880 40.000 60.480 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 80.280 40.000 80.880 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 212.200 40.000 212.800 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 1.400 40.000 2.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 130.600 40.000 131.200 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 126.520 40.000 127.120 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 9.560 40.000 10.160 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 91.160 40.000 91.760 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 216.280 40.000 216.880 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 296.000 23.370 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 87.080 40.000 87.680 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 289.720 40.000 290.320 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 138.760 40.000 139.360 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 185.000 40.000 185.600 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 220.360 40.000 220.960 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 122.440 40.000 123.040 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 228.520 40.000 229.120 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 36.760 40.000 37.360 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 72.120 40.000 72.720 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 107.480 40.000 108.080 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 193.160 40.000 193.760 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 149.640 40.000 150.240 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 17.720 40.000 18.320 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 266.600 40.000 267.200 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 231.240 40.000 231.840 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 170.040 40.000 170.640 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 199.960 40.000 200.560 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 40.840 40.000 41.440 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 258.440 40.000 259.040 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 296.000 7.730 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 180.920 40.000 181.520 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 63.960 40.000 64.560 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 134.680 40.000 135.280 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 99.320 40.000 99.920 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 13.640 40.000 14.240 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 161.880 40.000 162.480 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 282.920 40.000 283.520 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 235.320 40.000 235.920 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 103.400 40.000 104.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 189.080 40.000 189.680 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 247.560 40.000 248.160 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 297.880 40.000 298.480 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 118.360 40.000 118.960 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 296.000 33.490 300.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 49.000 40.000 49.600 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 32.680 40.000 33.280 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 296.000 17.850 300.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 157.800 40.000 158.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 5.480 40.000 6.080 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 243.480 40.000 244.080 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 44.920 40.000 45.520 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 296.000 4.970 300.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 296.000 2.210 300.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 68.040 40.000 68.640 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 208.120 40.000 208.720 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 4.285 10.795 39.875 288.405 ;
      LAYER met1 ;
        RECT 0.070 10.640 39.950 288.560 ;
      LAYER met2 ;
        RECT 0.100 295.720 1.650 299.725 ;
        RECT 2.490 295.720 4.410 299.725 ;
        RECT 5.250 295.720 7.170 299.725 ;
        RECT 8.010 295.720 9.930 299.725 ;
        RECT 10.770 295.720 11.770 299.725 ;
        RECT 12.610 295.720 14.530 299.725 ;
        RECT 15.370 295.720 17.290 299.725 ;
        RECT 18.130 295.720 20.050 299.725 ;
        RECT 20.890 295.720 22.810 299.725 ;
        RECT 23.650 295.720 25.570 299.725 ;
        RECT 26.410 295.720 28.330 299.725 ;
        RECT 29.170 295.720 30.170 299.725 ;
        RECT 31.010 295.720 32.930 299.725 ;
        RECT 33.770 295.720 35.690 299.725 ;
        RECT 36.530 295.720 38.450 299.725 ;
        RECT 39.290 295.720 39.920 299.725 ;
        RECT 0.100 4.280 39.920 295.720 ;
        RECT 0.650 2.875 1.650 4.280 ;
        RECT 2.490 2.875 4.410 4.280 ;
        RECT 5.250 2.875 7.170 4.280 ;
        RECT 8.010 2.875 9.930 4.280 ;
        RECT 10.770 2.875 12.690 4.280 ;
        RECT 13.530 2.875 15.450 4.280 ;
        RECT 16.290 2.875 18.210 4.280 ;
        RECT 19.050 2.875 20.050 4.280 ;
        RECT 20.890 2.875 22.810 4.280 ;
        RECT 23.650 2.875 25.570 4.280 ;
        RECT 26.410 2.875 28.330 4.280 ;
        RECT 29.170 2.875 31.090 4.280 ;
        RECT 31.930 2.875 33.850 4.280 ;
        RECT 34.690 2.875 36.610 4.280 ;
        RECT 37.450 2.875 38.450 4.280 ;
        RECT 39.290 2.875 39.920 4.280 ;
      LAYER met3 ;
        RECT 4.400 298.880 36.490 299.705 ;
        RECT 4.400 298.840 35.600 298.880 ;
        RECT 4.000 297.480 35.600 298.840 ;
        RECT 4.000 296.160 36.490 297.480 ;
        RECT 4.400 294.800 36.490 296.160 ;
        RECT 4.400 294.760 35.600 294.800 ;
        RECT 4.000 293.400 35.600 294.760 ;
        RECT 4.000 292.080 36.490 293.400 ;
        RECT 4.400 290.720 36.490 292.080 ;
        RECT 4.400 290.680 35.600 290.720 ;
        RECT 4.000 289.320 35.600 290.680 ;
        RECT 4.000 288.000 36.490 289.320 ;
        RECT 4.400 286.640 36.490 288.000 ;
        RECT 4.400 286.600 35.600 286.640 ;
        RECT 4.000 285.280 35.600 286.600 ;
        RECT 4.400 285.240 35.600 285.280 ;
        RECT 4.400 283.920 36.490 285.240 ;
        RECT 4.400 283.880 35.600 283.920 ;
        RECT 4.000 282.520 35.600 283.880 ;
        RECT 4.000 281.200 36.490 282.520 ;
        RECT 4.400 279.840 36.490 281.200 ;
        RECT 4.400 279.800 35.600 279.840 ;
        RECT 4.000 278.440 35.600 279.800 ;
        RECT 4.000 277.120 36.490 278.440 ;
        RECT 4.400 275.760 36.490 277.120 ;
        RECT 4.400 275.720 35.600 275.760 ;
        RECT 4.000 274.360 35.600 275.720 ;
        RECT 4.000 273.040 36.490 274.360 ;
        RECT 4.400 271.680 36.490 273.040 ;
        RECT 4.400 271.640 35.600 271.680 ;
        RECT 4.000 270.280 35.600 271.640 ;
        RECT 4.000 268.960 36.490 270.280 ;
        RECT 4.400 267.600 36.490 268.960 ;
        RECT 4.400 267.560 35.600 267.600 ;
        RECT 4.000 266.200 35.600 267.560 ;
        RECT 4.000 264.880 36.490 266.200 ;
        RECT 4.400 263.520 36.490 264.880 ;
        RECT 4.400 263.480 35.600 263.520 ;
        RECT 4.000 262.120 35.600 263.480 ;
        RECT 4.000 260.800 36.490 262.120 ;
        RECT 4.400 259.440 36.490 260.800 ;
        RECT 4.400 259.400 35.600 259.440 ;
        RECT 4.000 258.080 35.600 259.400 ;
        RECT 4.400 258.040 35.600 258.080 ;
        RECT 4.400 256.720 36.490 258.040 ;
        RECT 4.400 256.680 35.600 256.720 ;
        RECT 4.000 255.320 35.600 256.680 ;
        RECT 4.000 254.000 36.490 255.320 ;
        RECT 4.400 252.640 36.490 254.000 ;
        RECT 4.400 252.600 35.600 252.640 ;
        RECT 4.000 251.240 35.600 252.600 ;
        RECT 4.000 249.920 36.490 251.240 ;
        RECT 4.400 248.560 36.490 249.920 ;
        RECT 4.400 248.520 35.600 248.560 ;
        RECT 4.000 247.160 35.600 248.520 ;
        RECT 4.000 245.840 36.490 247.160 ;
        RECT 4.400 244.480 36.490 245.840 ;
        RECT 4.400 244.440 35.600 244.480 ;
        RECT 4.000 243.080 35.600 244.440 ;
        RECT 4.000 241.760 36.490 243.080 ;
        RECT 4.400 240.400 36.490 241.760 ;
        RECT 4.400 240.360 35.600 240.400 ;
        RECT 4.000 239.000 35.600 240.360 ;
        RECT 4.000 237.680 36.490 239.000 ;
        RECT 4.400 236.320 36.490 237.680 ;
        RECT 4.400 236.280 35.600 236.320 ;
        RECT 4.000 234.920 35.600 236.280 ;
        RECT 4.000 233.600 36.490 234.920 ;
        RECT 4.400 232.240 36.490 233.600 ;
        RECT 4.400 232.200 35.600 232.240 ;
        RECT 4.000 230.880 35.600 232.200 ;
        RECT 4.400 230.840 35.600 230.880 ;
        RECT 4.400 229.520 36.490 230.840 ;
        RECT 4.400 229.480 35.600 229.520 ;
        RECT 4.000 228.120 35.600 229.480 ;
        RECT 4.000 226.800 36.490 228.120 ;
        RECT 4.400 225.440 36.490 226.800 ;
        RECT 4.400 225.400 35.600 225.440 ;
        RECT 4.000 224.040 35.600 225.400 ;
        RECT 4.000 222.720 36.490 224.040 ;
        RECT 4.400 221.360 36.490 222.720 ;
        RECT 4.400 221.320 35.600 221.360 ;
        RECT 4.000 219.960 35.600 221.320 ;
        RECT 4.000 218.640 36.490 219.960 ;
        RECT 4.400 217.280 36.490 218.640 ;
        RECT 4.400 217.240 35.600 217.280 ;
        RECT 4.000 215.880 35.600 217.240 ;
        RECT 4.000 214.560 36.490 215.880 ;
        RECT 4.400 213.200 36.490 214.560 ;
        RECT 4.400 213.160 35.600 213.200 ;
        RECT 4.000 211.800 35.600 213.160 ;
        RECT 4.000 210.480 36.490 211.800 ;
        RECT 4.400 209.120 36.490 210.480 ;
        RECT 4.400 209.080 35.600 209.120 ;
        RECT 4.000 207.720 35.600 209.080 ;
        RECT 4.000 206.400 36.490 207.720 ;
        RECT 4.400 205.040 36.490 206.400 ;
        RECT 4.400 205.000 35.600 205.040 ;
        RECT 4.000 203.640 35.600 205.000 ;
        RECT 4.000 202.320 36.490 203.640 ;
        RECT 4.400 200.960 36.490 202.320 ;
        RECT 4.400 200.920 35.600 200.960 ;
        RECT 4.000 199.600 35.600 200.920 ;
        RECT 4.400 199.560 35.600 199.600 ;
        RECT 4.400 198.240 36.490 199.560 ;
        RECT 4.400 198.200 35.600 198.240 ;
        RECT 4.000 196.840 35.600 198.200 ;
        RECT 4.000 195.520 36.490 196.840 ;
        RECT 4.400 194.160 36.490 195.520 ;
        RECT 4.400 194.120 35.600 194.160 ;
        RECT 4.000 192.760 35.600 194.120 ;
        RECT 4.000 191.440 36.490 192.760 ;
        RECT 4.400 190.080 36.490 191.440 ;
        RECT 4.400 190.040 35.600 190.080 ;
        RECT 4.000 188.680 35.600 190.040 ;
        RECT 4.000 187.360 36.490 188.680 ;
        RECT 4.400 186.000 36.490 187.360 ;
        RECT 4.400 185.960 35.600 186.000 ;
        RECT 4.000 184.600 35.600 185.960 ;
        RECT 4.000 183.280 36.490 184.600 ;
        RECT 4.400 181.920 36.490 183.280 ;
        RECT 4.400 181.880 35.600 181.920 ;
        RECT 4.000 180.520 35.600 181.880 ;
        RECT 4.000 179.200 36.490 180.520 ;
        RECT 4.400 177.840 36.490 179.200 ;
        RECT 4.400 177.800 35.600 177.840 ;
        RECT 4.000 176.440 35.600 177.800 ;
        RECT 4.000 175.120 36.490 176.440 ;
        RECT 4.400 173.760 36.490 175.120 ;
        RECT 4.400 173.720 35.600 173.760 ;
        RECT 4.000 172.400 35.600 173.720 ;
        RECT 4.400 172.360 35.600 172.400 ;
        RECT 4.400 171.040 36.490 172.360 ;
        RECT 4.400 171.000 35.600 171.040 ;
        RECT 4.000 169.640 35.600 171.000 ;
        RECT 4.000 168.320 36.490 169.640 ;
        RECT 4.400 166.960 36.490 168.320 ;
        RECT 4.400 166.920 35.600 166.960 ;
        RECT 4.000 165.560 35.600 166.920 ;
        RECT 4.000 164.240 36.490 165.560 ;
        RECT 4.400 162.880 36.490 164.240 ;
        RECT 4.400 162.840 35.600 162.880 ;
        RECT 4.000 161.480 35.600 162.840 ;
        RECT 4.000 160.160 36.490 161.480 ;
        RECT 4.400 158.800 36.490 160.160 ;
        RECT 4.400 158.760 35.600 158.800 ;
        RECT 4.000 157.400 35.600 158.760 ;
        RECT 4.000 156.080 36.490 157.400 ;
        RECT 4.400 154.720 36.490 156.080 ;
        RECT 4.400 154.680 35.600 154.720 ;
        RECT 4.000 153.320 35.600 154.680 ;
        RECT 4.000 152.000 36.490 153.320 ;
        RECT 4.400 150.640 36.490 152.000 ;
        RECT 4.400 150.600 35.600 150.640 ;
        RECT 4.000 149.240 35.600 150.600 ;
        RECT 4.000 147.920 36.490 149.240 ;
        RECT 4.400 146.560 36.490 147.920 ;
        RECT 4.400 146.520 35.600 146.560 ;
        RECT 4.000 145.160 35.600 146.520 ;
        RECT 4.000 143.840 36.490 145.160 ;
        RECT 4.400 142.480 36.490 143.840 ;
        RECT 4.400 142.440 35.600 142.480 ;
        RECT 4.000 141.120 35.600 142.440 ;
        RECT 4.400 141.080 35.600 141.120 ;
        RECT 4.400 139.760 36.490 141.080 ;
        RECT 4.400 139.720 35.600 139.760 ;
        RECT 4.000 138.360 35.600 139.720 ;
        RECT 4.000 137.040 36.490 138.360 ;
        RECT 4.400 135.680 36.490 137.040 ;
        RECT 4.400 135.640 35.600 135.680 ;
        RECT 4.000 134.280 35.600 135.640 ;
        RECT 4.000 132.960 36.490 134.280 ;
        RECT 4.400 131.600 36.490 132.960 ;
        RECT 4.400 131.560 35.600 131.600 ;
        RECT 4.000 130.200 35.600 131.560 ;
        RECT 4.000 128.880 36.490 130.200 ;
        RECT 4.400 127.520 36.490 128.880 ;
        RECT 4.400 127.480 35.600 127.520 ;
        RECT 4.000 126.120 35.600 127.480 ;
        RECT 4.000 124.800 36.490 126.120 ;
        RECT 4.400 123.440 36.490 124.800 ;
        RECT 4.400 123.400 35.600 123.440 ;
        RECT 4.000 122.040 35.600 123.400 ;
        RECT 4.000 120.720 36.490 122.040 ;
        RECT 4.400 119.360 36.490 120.720 ;
        RECT 4.400 119.320 35.600 119.360 ;
        RECT 4.000 117.960 35.600 119.320 ;
        RECT 4.000 116.640 36.490 117.960 ;
        RECT 4.400 115.280 36.490 116.640 ;
        RECT 4.400 115.240 35.600 115.280 ;
        RECT 4.000 113.920 35.600 115.240 ;
        RECT 4.400 113.880 35.600 113.920 ;
        RECT 4.400 112.560 36.490 113.880 ;
        RECT 4.400 112.520 35.600 112.560 ;
        RECT 4.000 111.160 35.600 112.520 ;
        RECT 4.000 109.840 36.490 111.160 ;
        RECT 4.400 108.480 36.490 109.840 ;
        RECT 4.400 108.440 35.600 108.480 ;
        RECT 4.000 107.080 35.600 108.440 ;
        RECT 4.000 105.760 36.490 107.080 ;
        RECT 4.400 104.400 36.490 105.760 ;
        RECT 4.400 104.360 35.600 104.400 ;
        RECT 4.000 103.000 35.600 104.360 ;
        RECT 4.000 101.680 36.490 103.000 ;
        RECT 4.400 100.320 36.490 101.680 ;
        RECT 4.400 100.280 35.600 100.320 ;
        RECT 4.000 98.920 35.600 100.280 ;
        RECT 4.000 97.600 36.490 98.920 ;
        RECT 4.400 96.240 36.490 97.600 ;
        RECT 4.400 96.200 35.600 96.240 ;
        RECT 4.000 94.840 35.600 96.200 ;
        RECT 4.000 93.520 36.490 94.840 ;
        RECT 4.400 92.160 36.490 93.520 ;
        RECT 4.400 92.120 35.600 92.160 ;
        RECT 4.000 90.760 35.600 92.120 ;
        RECT 4.000 89.440 36.490 90.760 ;
        RECT 4.400 88.080 36.490 89.440 ;
        RECT 4.400 88.040 35.600 88.080 ;
        RECT 4.000 86.720 35.600 88.040 ;
        RECT 4.400 86.680 35.600 86.720 ;
        RECT 4.400 85.360 36.490 86.680 ;
        RECT 4.400 85.320 35.600 85.360 ;
        RECT 4.000 83.960 35.600 85.320 ;
        RECT 4.000 82.640 36.490 83.960 ;
        RECT 4.400 81.280 36.490 82.640 ;
        RECT 4.400 81.240 35.600 81.280 ;
        RECT 4.000 79.880 35.600 81.240 ;
        RECT 4.000 78.560 36.490 79.880 ;
        RECT 4.400 77.200 36.490 78.560 ;
        RECT 4.400 77.160 35.600 77.200 ;
        RECT 4.000 75.800 35.600 77.160 ;
        RECT 4.000 74.480 36.490 75.800 ;
        RECT 4.400 73.120 36.490 74.480 ;
        RECT 4.400 73.080 35.600 73.120 ;
        RECT 4.000 71.720 35.600 73.080 ;
        RECT 4.000 70.400 36.490 71.720 ;
        RECT 4.400 69.040 36.490 70.400 ;
        RECT 4.400 69.000 35.600 69.040 ;
        RECT 4.000 67.640 35.600 69.000 ;
        RECT 4.000 66.320 36.490 67.640 ;
        RECT 4.400 64.960 36.490 66.320 ;
        RECT 4.400 64.920 35.600 64.960 ;
        RECT 4.000 63.560 35.600 64.920 ;
        RECT 4.000 62.240 36.490 63.560 ;
        RECT 4.400 60.880 36.490 62.240 ;
        RECT 4.400 60.840 35.600 60.880 ;
        RECT 4.000 59.480 35.600 60.840 ;
        RECT 4.000 58.160 36.490 59.480 ;
        RECT 4.400 56.800 36.490 58.160 ;
        RECT 4.400 56.760 35.600 56.800 ;
        RECT 4.000 55.440 35.600 56.760 ;
        RECT 4.400 55.400 35.600 55.440 ;
        RECT 4.400 54.080 36.490 55.400 ;
        RECT 4.400 54.040 35.600 54.080 ;
        RECT 4.000 52.680 35.600 54.040 ;
        RECT 4.000 51.360 36.490 52.680 ;
        RECT 4.400 50.000 36.490 51.360 ;
        RECT 4.400 49.960 35.600 50.000 ;
        RECT 4.000 48.600 35.600 49.960 ;
        RECT 4.000 47.280 36.490 48.600 ;
        RECT 4.400 45.920 36.490 47.280 ;
        RECT 4.400 45.880 35.600 45.920 ;
        RECT 4.000 44.520 35.600 45.880 ;
        RECT 4.000 43.200 36.490 44.520 ;
        RECT 4.400 41.840 36.490 43.200 ;
        RECT 4.400 41.800 35.600 41.840 ;
        RECT 4.000 40.440 35.600 41.800 ;
        RECT 4.000 39.120 36.490 40.440 ;
        RECT 4.400 37.760 36.490 39.120 ;
        RECT 4.400 37.720 35.600 37.760 ;
        RECT 4.000 36.360 35.600 37.720 ;
        RECT 4.000 35.040 36.490 36.360 ;
        RECT 4.400 33.680 36.490 35.040 ;
        RECT 4.400 33.640 35.600 33.680 ;
        RECT 4.000 32.280 35.600 33.640 ;
        RECT 4.000 30.960 36.490 32.280 ;
        RECT 4.400 29.600 36.490 30.960 ;
        RECT 4.400 29.560 35.600 29.600 ;
        RECT 4.000 28.240 35.600 29.560 ;
        RECT 4.400 28.200 35.600 28.240 ;
        RECT 4.400 26.880 36.490 28.200 ;
        RECT 4.400 26.840 35.600 26.880 ;
        RECT 4.000 25.480 35.600 26.840 ;
        RECT 4.000 24.160 36.490 25.480 ;
        RECT 4.400 22.800 36.490 24.160 ;
        RECT 4.400 22.760 35.600 22.800 ;
        RECT 4.000 21.400 35.600 22.760 ;
        RECT 4.000 20.080 36.490 21.400 ;
        RECT 4.400 18.720 36.490 20.080 ;
        RECT 4.400 18.680 35.600 18.720 ;
        RECT 4.000 17.320 35.600 18.680 ;
        RECT 4.000 16.000 36.490 17.320 ;
        RECT 4.400 14.640 36.490 16.000 ;
        RECT 4.400 14.600 35.600 14.640 ;
        RECT 4.000 13.240 35.600 14.600 ;
        RECT 4.000 11.920 36.490 13.240 ;
        RECT 4.400 10.560 36.490 11.920 ;
        RECT 4.400 10.520 35.600 10.560 ;
        RECT 4.000 9.160 35.600 10.520 ;
        RECT 4.000 7.840 36.490 9.160 ;
        RECT 4.400 6.480 36.490 7.840 ;
        RECT 4.400 6.440 35.600 6.480 ;
        RECT 4.000 5.080 35.600 6.440 ;
        RECT 4.000 3.760 36.490 5.080 ;
        RECT 4.400 2.400 36.490 3.760 ;
        RECT 4.400 2.360 35.600 2.400 ;
        RECT 4.000 1.550 35.600 2.360 ;
      LAYER met4 ;
        RECT 7.655 10.640 9.145 288.560 ;
        RECT 11.545 10.640 13.970 288.560 ;
        RECT 16.370 10.640 18.795 288.560 ;
        RECT 21.195 10.640 23.625 288.560 ;
        RECT 26.025 10.640 27.305 288.560 ;
  END
END wb_openram_wrapper
END LIBRARY

