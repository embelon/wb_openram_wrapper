magic
tech sky130A
magscale 1 2
timestamp 1647558821
<< viali >>
rect 27445 77673 27479 77707
rect 28181 77673 28215 77707
rect 1409 77537 1443 77571
rect 3801 77537 3835 77571
rect 1685 77469 1719 77503
rect 4077 77469 4111 77503
rect 27261 77469 27295 77503
rect 27997 77469 28031 77503
rect 28733 77469 28767 77503
rect 29837 77469 29871 77503
rect 28917 77333 28951 77367
rect 30021 77333 30055 77367
rect 28549 77129 28583 77163
rect 29285 77129 29319 77163
rect 2697 76993 2731 77027
rect 28365 76993 28399 77027
rect 29101 76993 29135 77027
rect 29837 76993 29871 77027
rect 1409 76925 1443 76959
rect 1685 76925 1719 76959
rect 2973 76925 3007 76959
rect 30021 76789 30055 76823
rect 28917 76585 28951 76619
rect 1409 76449 1443 76483
rect 1685 76381 1719 76415
rect 2881 76381 2915 76415
rect 28733 76381 28767 76415
rect 29837 76381 29871 76415
rect 2697 76245 2731 76279
rect 30021 76245 30055 76279
rect 1409 76041 1443 76075
rect 29285 76041 29319 76075
rect 14657 75973 14691 76007
rect 1593 75905 1627 75939
rect 14473 75905 14507 75939
rect 15853 75905 15887 75939
rect 16865 75905 16899 75939
rect 19073 75905 19107 75939
rect 19993 75905 20027 75939
rect 20085 75905 20119 75939
rect 20177 75905 20211 75939
rect 20361 75905 20395 75939
rect 29101 75905 29135 75939
rect 29837 75905 29871 75939
rect 14841 75769 14875 75803
rect 16037 75701 16071 75735
rect 17049 75701 17083 75735
rect 19257 75701 19291 75735
rect 19717 75701 19751 75735
rect 30021 75701 30055 75735
rect 14749 75497 14783 75531
rect 21189 75497 21223 75531
rect 15209 75361 15243 75395
rect 17141 75361 17175 75395
rect 19809 75361 19843 75395
rect 1593 75293 1627 75327
rect 14565 75293 14599 75327
rect 20065 75293 20099 75327
rect 29837 75293 29871 75327
rect 14381 75225 14415 75259
rect 15476 75225 15510 75259
rect 17386 75225 17420 75259
rect 1409 75157 1443 75191
rect 16589 75157 16623 75191
rect 18521 75157 18555 75191
rect 30021 75157 30055 75191
rect 14841 74953 14875 74987
rect 15669 74953 15703 74987
rect 14657 74885 14691 74919
rect 17233 74885 17267 74919
rect 1593 74817 1627 74851
rect 14473 74817 14507 74851
rect 15301 74817 15335 74851
rect 15485 74817 15519 74851
rect 17049 74817 17083 74851
rect 18501 74817 18535 74851
rect 20913 74817 20947 74851
rect 21005 74817 21039 74851
rect 21097 74817 21131 74851
rect 21281 74817 21315 74851
rect 22089 74817 22123 74851
rect 29837 74817 29871 74851
rect 17325 74749 17359 74783
rect 18245 74749 18279 74783
rect 21833 74749 21867 74783
rect 1409 74681 1443 74715
rect 16773 74681 16807 74715
rect 19625 74613 19659 74647
rect 20637 74613 20671 74647
rect 23213 74613 23247 74647
rect 30021 74613 30055 74647
rect 16037 74409 16071 74443
rect 17509 74409 17543 74443
rect 20637 74409 20671 74443
rect 14933 74341 14967 74375
rect 18061 74341 18095 74375
rect 19349 74341 19383 74375
rect 16497 74273 16531 74307
rect 18613 74273 18647 74307
rect 17325 74205 17359 74239
rect 20453 74205 20487 74239
rect 21189 74205 21223 74239
rect 21445 74205 21479 74239
rect 29837 74205 29871 74239
rect 14565 74137 14599 74171
rect 14749 74137 14783 74171
rect 16589 74137 16623 74171
rect 18337 74137 18371 74171
rect 19625 74137 19659 74171
rect 19901 74137 19935 74171
rect 16497 74069 16531 74103
rect 18521 74069 18555 74103
rect 19809 74069 19843 74103
rect 22569 74069 22603 74103
rect 30021 74069 30055 74103
rect 13737 73865 13771 73899
rect 16681 73865 16715 73899
rect 17969 73865 18003 73899
rect 19717 73865 19751 73899
rect 20637 73865 20671 73899
rect 19533 73797 19567 73831
rect 1593 73729 1627 73763
rect 13921 73729 13955 73763
rect 16957 73729 16991 73763
rect 17049 73729 17083 73763
rect 17141 73729 17175 73763
rect 17337 73729 17371 73763
rect 18245 73729 18279 73763
rect 18337 73729 18371 73763
rect 18429 73729 18463 73763
rect 18613 73729 18647 73763
rect 20913 73729 20947 73763
rect 21005 73729 21039 73763
rect 21097 73729 21131 73763
rect 21281 73729 21315 73763
rect 29837 73729 29871 73763
rect 19809 73661 19843 73695
rect 1409 73593 1443 73627
rect 19257 73593 19291 73627
rect 30021 73525 30055 73559
rect 15025 73321 15059 73355
rect 18613 73321 18647 73355
rect 19809 73321 19843 73355
rect 20729 73321 20763 73355
rect 1593 73117 1627 73151
rect 15669 73117 15703 73151
rect 15853 73117 15887 73151
rect 17029 73117 17063 73151
rect 17138 73114 17172 73148
rect 17233 73117 17267 73151
rect 17417 73117 17451 73151
rect 20545 73117 20579 73151
rect 29837 73117 29871 73151
rect 14657 73049 14691 73083
rect 14841 73049 14875 73083
rect 15485 73049 15519 73083
rect 16773 73049 16807 73083
rect 18521 73049 18555 73083
rect 19717 73049 19751 73083
rect 1409 72981 1443 73015
rect 30021 72981 30055 73015
rect 14841 72709 14875 72743
rect 16129 72709 16163 72743
rect 1593 72641 1627 72675
rect 14657 72641 14691 72675
rect 15945 72641 15979 72675
rect 17141 72641 17175 72675
rect 29837 72641 29871 72675
rect 15025 72505 15059 72539
rect 1409 72437 1443 72471
rect 17233 72437 17267 72471
rect 30021 72437 30055 72471
rect 13369 72233 13403 72267
rect 1409 72165 1443 72199
rect 1593 72029 1627 72063
rect 13553 72029 13587 72063
rect 14657 72029 14691 72063
rect 14841 72029 14875 72063
rect 17141 72029 17175 72063
rect 17233 72029 17267 72063
rect 17325 72029 17359 72063
rect 17509 72029 17543 72063
rect 29837 72029 29871 72063
rect 15025 71961 15059 71995
rect 16865 71893 16899 71927
rect 30021 71893 30055 71927
rect 13001 71621 13035 71655
rect 20177 71621 20211 71655
rect 12817 71553 12851 71587
rect 17555 71553 17589 71587
rect 17693 71553 17727 71587
rect 17790 71553 17824 71587
rect 17969 71553 18003 71587
rect 21005 71553 21039 71587
rect 29837 71553 29871 71587
rect 13185 71417 13219 71451
rect 17325 71349 17359 71383
rect 20269 71349 20303 71383
rect 21097 71349 21131 71383
rect 30021 71349 30055 71383
rect 15025 71145 15059 71179
rect 18245 71145 18279 71179
rect 20913 71145 20947 71179
rect 13185 71077 13219 71111
rect 16313 71009 16347 71043
rect 1409 70941 1443 70975
rect 1685 70941 1719 70975
rect 13001 70941 13035 70975
rect 14841 70941 14875 70975
rect 29837 70941 29871 70975
rect 12817 70873 12851 70907
rect 14657 70873 14691 70907
rect 16405 70873 16439 70907
rect 16957 70873 16991 70907
rect 19625 70873 19659 70907
rect 15835 70805 15869 70839
rect 16313 70805 16347 70839
rect 30021 70805 30055 70839
rect 1409 70601 1443 70635
rect 12173 70601 12207 70635
rect 15117 70601 15151 70635
rect 18245 70601 18279 70635
rect 19993 70601 20027 70635
rect 13001 70533 13035 70567
rect 13185 70533 13219 70567
rect 1593 70465 1627 70499
rect 12357 70465 12391 70499
rect 12817 70465 12851 70499
rect 13645 70465 13679 70499
rect 13829 70465 13863 70499
rect 14933 70465 14967 70499
rect 15577 70465 15611 70499
rect 16865 70465 16899 70499
rect 17121 70465 17155 70499
rect 18705 70465 18739 70499
rect 20913 70465 20947 70499
rect 22063 70465 22097 70499
rect 22198 70468 22232 70502
rect 22298 70465 22332 70499
rect 22477 70465 22511 70499
rect 29837 70465 29871 70499
rect 14013 70397 14047 70431
rect 15761 70261 15795 70295
rect 21097 70261 21131 70295
rect 21833 70261 21867 70295
rect 30021 70261 30055 70295
rect 13185 70057 13219 70091
rect 19349 70057 19383 70091
rect 21833 70057 21867 70091
rect 1593 69853 1627 69887
rect 12817 69853 12851 69887
rect 14749 69853 14783 69887
rect 20453 69853 20487 69887
rect 22293 69853 22327 69887
rect 29837 69853 29871 69887
rect 13001 69785 13035 69819
rect 14994 69785 15028 69819
rect 16681 69785 16715 69819
rect 19625 69785 19659 69819
rect 19809 69785 19843 69819
rect 19901 69785 19935 69819
rect 20720 69785 20754 69819
rect 22538 69785 22572 69819
rect 1409 69717 1443 69751
rect 16129 69717 16163 69751
rect 17969 69717 18003 69751
rect 23673 69717 23707 69751
rect 30021 69717 30055 69751
rect 21833 69513 21867 69547
rect 13001 69445 13035 69479
rect 18398 69445 18432 69479
rect 20269 69445 20303 69479
rect 1593 69377 1627 69411
rect 12817 69377 12851 69411
rect 14177 69377 14211 69411
rect 17141 69377 17175 69411
rect 20085 69377 20119 69411
rect 21097 69377 21131 69411
rect 22109 69377 22143 69411
rect 22201 69377 22235 69411
rect 22293 69377 22327 69411
rect 22477 69377 22511 69411
rect 29101 69377 29135 69411
rect 29837 69377 29871 69411
rect 13921 69309 13955 69343
rect 16865 69309 16899 69343
rect 18153 69309 18187 69343
rect 21281 69241 21315 69275
rect 29285 69241 29319 69275
rect 1409 69173 1443 69207
rect 13185 69173 13219 69207
rect 15301 69173 15335 69207
rect 19533 69173 19567 69207
rect 30021 69173 30055 69207
rect 14657 68969 14691 69003
rect 17049 68969 17083 69003
rect 19993 68969 20027 69003
rect 22017 68969 22051 69003
rect 17601 68833 17635 68867
rect 20453 68833 20487 68867
rect 21373 68833 21407 68867
rect 1593 68765 1627 68799
rect 12633 68765 12667 68799
rect 14933 68765 14967 68799
rect 15025 68765 15059 68799
rect 15117 68765 15151 68799
rect 15301 68765 15335 68799
rect 18429 68765 18463 68799
rect 21833 68765 21867 68799
rect 28733 68765 28767 68799
rect 29837 68765 29871 68799
rect 12817 68697 12851 68731
rect 17325 68697 17359 68731
rect 18613 68697 18647 68731
rect 20453 68697 20487 68731
rect 20545 68697 20579 68731
rect 21189 68697 21223 68731
rect 1409 68629 1443 68663
rect 13001 68629 13035 68663
rect 17509 68629 17543 68663
rect 28917 68629 28951 68663
rect 30021 68629 30055 68663
rect 13369 68425 13403 68459
rect 20545 68425 20579 68459
rect 26985 68425 27019 68459
rect 17325 68357 17359 68391
rect 19533 68357 19567 68391
rect 20361 68357 20395 68391
rect 13185 68289 13219 68323
rect 14085 68289 14119 68323
rect 14194 68289 14228 68323
rect 14310 68289 14344 68323
rect 14473 68289 14507 68323
rect 19349 68289 19383 68323
rect 27215 68289 27249 68323
rect 27353 68289 27387 68323
rect 27445 68289 27479 68323
rect 27629 68289 27663 68323
rect 29837 68289 29871 68323
rect 20637 68221 20671 68255
rect 13829 68153 13863 68187
rect 20085 68153 20119 68187
rect 17417 68085 17451 68119
rect 30021 68085 30055 68119
rect 18521 67881 18555 67915
rect 26249 67881 26283 67915
rect 27353 67881 27387 67915
rect 1409 67813 1443 67847
rect 21281 67813 21315 67847
rect 24869 67813 24903 67847
rect 28917 67813 28951 67847
rect 30021 67813 30055 67847
rect 1593 67677 1627 67711
rect 12909 67677 12943 67711
rect 16681 67677 16715 67711
rect 17417 67677 17451 67711
rect 18337 67677 18371 67711
rect 25053 67677 25087 67711
rect 25329 67677 25363 67711
rect 26505 67677 26539 67711
rect 26614 67677 26648 67711
rect 26709 67677 26743 67711
rect 26893 67677 26927 67711
rect 27629 67677 27663 67711
rect 27721 67677 27755 67711
rect 27813 67677 27847 67711
rect 27997 67677 28031 67711
rect 28733 67677 28767 67711
rect 29837 67677 29871 67711
rect 12725 67609 12759 67643
rect 17601 67609 17635 67643
rect 19993 67609 20027 67643
rect 25237 67609 25271 67643
rect 13093 67541 13127 67575
rect 16773 67541 16807 67575
rect 19165 67337 19199 67371
rect 24869 67337 24903 67371
rect 12817 67269 12851 67303
rect 18981 67269 19015 67303
rect 1593 67201 1627 67235
rect 12633 67201 12667 67235
rect 15071 67201 15105 67235
rect 15206 67201 15240 67235
rect 15306 67201 15340 67235
rect 15485 67201 15519 67235
rect 23305 67201 23339 67235
rect 23489 67201 23523 67235
rect 25053 67201 25087 67235
rect 25237 67201 25271 67235
rect 25329 67201 25363 67235
rect 25973 67201 26007 67235
rect 26157 67201 26191 67235
rect 26249 67201 26283 67235
rect 27261 67201 27295 67235
rect 27350 67201 27384 67235
rect 27450 67201 27484 67235
rect 27629 67201 27663 67235
rect 29101 67201 29135 67235
rect 29837 67201 29871 67235
rect 19257 67133 19291 67167
rect 25789 67133 25823 67167
rect 18705 67065 18739 67099
rect 1409 66997 1443 67031
rect 13001 66997 13035 67031
rect 14841 66997 14875 67031
rect 23673 66997 23707 67031
rect 26985 66997 27019 67031
rect 29285 66997 29319 67031
rect 30021 66997 30055 67031
rect 18429 66793 18463 66827
rect 19441 66793 19475 66827
rect 26433 66793 26467 66827
rect 16681 66725 16715 66759
rect 25329 66725 25363 66759
rect 22385 66657 22419 66691
rect 24409 66657 24443 66691
rect 27813 66657 27847 66691
rect 1593 66589 1627 66623
rect 14381 66589 14415 66623
rect 14473 66589 14507 66623
rect 14565 66589 14599 66623
rect 14749 66589 14783 66623
rect 15301 66589 15335 66623
rect 15557 66589 15591 66623
rect 17397 66589 17431 66623
rect 17509 66589 17543 66623
rect 17601 66589 17635 66623
rect 17785 66589 17819 66623
rect 18245 66589 18279 66623
rect 19257 66589 19291 66623
rect 20545 66589 20579 66623
rect 22569 66589 22603 66623
rect 23397 66589 23431 66623
rect 23489 66589 23523 66623
rect 24593 66589 24627 66623
rect 25513 66589 25547 66623
rect 25789 66589 25823 66623
rect 26709 66589 26743 66623
rect 26801 66589 26835 66623
rect 26893 66589 26927 66623
rect 27089 66589 27123 66623
rect 27537 66589 27571 66623
rect 29837 66589 29871 66623
rect 1409 66453 1443 66487
rect 14105 66453 14139 66487
rect 17141 66453 17175 66487
rect 20729 66453 20763 66487
rect 22753 66453 22787 66487
rect 23673 66453 23707 66487
rect 24777 66453 24811 66487
rect 25697 66453 25731 66487
rect 30021 66453 30055 66487
rect 25053 66249 25087 66283
rect 12817 66181 12851 66215
rect 14004 66181 14038 66215
rect 17294 66181 17328 66215
rect 23673 66181 23707 66215
rect 30113 66181 30147 66215
rect 1593 66113 1627 66147
rect 12633 66113 12667 66147
rect 15945 66113 15979 66147
rect 19533 66113 19567 66147
rect 22063 66113 22097 66147
rect 22182 66116 22216 66150
rect 22293 66113 22327 66147
rect 22477 66113 22511 66147
rect 23305 66113 23339 66147
rect 23489 66113 23523 66147
rect 25237 66113 25271 66147
rect 25421 66113 25455 66147
rect 25513 66113 25547 66147
rect 27905 66113 27939 66147
rect 28641 66113 28675 66147
rect 29377 66113 29411 66147
rect 29561 66113 29595 66147
rect 29653 66113 29687 66147
rect 29929 66113 29963 66147
rect 13737 66045 13771 66079
rect 17049 66045 17083 66079
rect 29745 66045 29779 66079
rect 16129 65977 16163 66011
rect 20821 65977 20855 66011
rect 1409 65909 1443 65943
rect 13001 65909 13035 65943
rect 15117 65909 15151 65943
rect 18429 65909 18463 65943
rect 21833 65909 21867 65943
rect 28089 65909 28123 65943
rect 28825 65909 28859 65943
rect 12725 65705 12759 65739
rect 15485 65705 15519 65739
rect 16865 65705 16899 65739
rect 18153 65705 18187 65739
rect 19441 65705 19475 65739
rect 19993 65705 20027 65739
rect 27445 65705 27479 65739
rect 28733 65705 28767 65739
rect 17325 65569 17359 65603
rect 17417 65569 17451 65603
rect 20545 65569 20579 65603
rect 21373 65569 21407 65603
rect 25237 65569 25271 65603
rect 1593 65501 1627 65535
rect 12909 65501 12943 65535
rect 15301 65501 15335 65535
rect 17969 65501 18003 65535
rect 19257 65501 19291 65535
rect 24961 65501 24995 65535
rect 27721 65501 27755 65535
rect 27813 65501 27847 65535
rect 27905 65501 27939 65535
rect 28089 65501 28123 65535
rect 29837 65501 29871 65535
rect 20269 65433 20303 65467
rect 21618 65433 21652 65467
rect 28641 65433 28675 65467
rect 1409 65365 1443 65399
rect 17325 65365 17359 65399
rect 20453 65365 20487 65399
rect 22753 65365 22787 65399
rect 30021 65365 30055 65399
rect 13921 65161 13955 65195
rect 15467 65161 15501 65195
rect 15945 65161 15979 65195
rect 18705 65161 18739 65195
rect 23213 65161 23247 65195
rect 25973 65161 26007 65195
rect 17509 65093 17543 65127
rect 19257 65093 19291 65127
rect 19441 65093 19475 65127
rect 20453 65093 20487 65127
rect 20545 65093 20579 65127
rect 22078 65093 22112 65127
rect 12909 65025 12943 65059
rect 13737 65025 13771 65059
rect 15761 65025 15795 65059
rect 17325 65025 17359 65059
rect 18521 65025 18555 65059
rect 20269 65025 20303 65059
rect 21097 65025 21131 65059
rect 26157 65025 26191 65059
rect 26341 65025 26375 65059
rect 26433 65025 26467 65059
rect 29561 65025 29595 65059
rect 16037 64957 16071 64991
rect 21833 64957 21867 64991
rect 27997 64957 28031 64991
rect 28273 64957 28307 64991
rect 29285 64957 29319 64991
rect 19993 64889 20027 64923
rect 21281 64889 21315 64923
rect 12725 64821 12759 64855
rect 19441 64617 19475 64651
rect 20085 64617 20119 64651
rect 21189 64617 21223 64651
rect 27353 64617 27387 64651
rect 28089 64481 28123 64515
rect 1593 64413 1627 64447
rect 12909 64413 12943 64447
rect 19257 64413 19291 64447
rect 21465 64413 21499 64447
rect 21557 64413 21591 64447
rect 21649 64413 21683 64447
rect 21833 64413 21867 64447
rect 23397 64413 23431 64447
rect 23581 64413 23615 64447
rect 24869 64413 24903 64447
rect 25145 64413 25179 64447
rect 25881 64413 25915 64447
rect 26157 64413 26191 64447
rect 26617 64413 26651 64447
rect 26801 64413 26835 64447
rect 26893 64413 26927 64447
rect 26985 64413 27019 64447
rect 27169 64413 27203 64447
rect 27813 64413 27847 64447
rect 12725 64345 12759 64379
rect 19993 64345 20027 64379
rect 25053 64345 25087 64379
rect 25697 64345 25731 64379
rect 29929 64345 29963 64379
rect 1409 64277 1443 64311
rect 13093 64277 13127 64311
rect 23765 64277 23799 64311
rect 24685 64277 24719 64311
rect 26065 64277 26099 64311
rect 30021 64277 30055 64311
rect 26985 64073 27019 64107
rect 28917 64073 28951 64107
rect 30113 64073 30147 64107
rect 12173 64005 12207 64039
rect 13001 64005 13035 64039
rect 14473 64005 14507 64039
rect 19809 64005 19843 64039
rect 19993 64005 20027 64039
rect 20729 64005 20763 64039
rect 1593 63937 1627 63971
rect 11989 63937 12023 63971
rect 12817 63937 12851 63971
rect 14289 63937 14323 63971
rect 17141 63937 17175 63971
rect 20545 63937 20579 63971
rect 23397 63937 23431 63971
rect 23581 63937 23615 63971
rect 25237 63937 25271 63971
rect 27261 63937 27295 63971
rect 27350 63937 27384 63971
rect 27445 63937 27479 63971
rect 27629 63937 27663 63971
rect 28181 63937 28215 63971
rect 28365 63937 28399 63971
rect 28733 63937 28767 63971
rect 29377 63937 29411 63971
rect 29561 63937 29595 63971
rect 29653 63937 29687 63971
rect 29929 63937 29963 63971
rect 12357 63869 12391 63903
rect 14565 63869 14599 63903
rect 17325 63869 17359 63903
rect 24961 63869 24995 63903
rect 28457 63869 28491 63903
rect 28549 63869 28583 63903
rect 29745 63869 29779 63903
rect 14013 63801 14047 63835
rect 23765 63801 23799 63835
rect 1409 63733 1443 63767
rect 13185 63733 13219 63767
rect 14197 63461 14231 63495
rect 15577 63461 15611 63495
rect 16773 63461 16807 63495
rect 19901 63461 19935 63495
rect 23305 63461 23339 63495
rect 27537 63461 27571 63495
rect 29009 63461 29043 63495
rect 13185 63393 13219 63427
rect 14657 63393 14691 63427
rect 20269 63393 20303 63427
rect 20453 63393 20487 63427
rect 24593 63393 24627 63427
rect 28543 63393 28577 63427
rect 1593 63325 1627 63359
rect 13001 63325 13035 63359
rect 23489 63325 23523 63359
rect 24869 63325 24903 63359
rect 25973 63325 26007 63359
rect 26801 63325 26835 63359
rect 27353 63325 27387 63359
rect 28273 63325 28307 63359
rect 28457 63325 28491 63359
rect 28641 63325 28675 63359
rect 28825 63325 28859 63359
rect 29837 63325 29871 63359
rect 12817 63257 12851 63291
rect 14749 63257 14783 63291
rect 15393 63257 15427 63291
rect 16589 63257 16623 63291
rect 27997 63257 28031 63291
rect 1409 63189 1443 63223
rect 14657 63189 14691 63223
rect 20361 63189 20395 63223
rect 26065 63189 26099 63223
rect 26985 63189 27019 63223
rect 30021 63189 30055 63223
rect 27721 62985 27755 63019
rect 30113 62985 30147 63019
rect 12817 62917 12851 62951
rect 13001 62917 13035 62951
rect 1593 62849 1627 62883
rect 12633 62849 12667 62883
rect 17463 62849 17497 62883
rect 17582 62852 17616 62886
rect 17714 62852 17748 62886
rect 17877 62849 17911 62883
rect 19349 62849 19383 62883
rect 20361 62849 20395 62883
rect 23581 62849 23615 62883
rect 26985 62849 27019 62883
rect 27951 62849 27985 62883
rect 28070 62849 28104 62883
rect 28202 62849 28236 62883
rect 28365 62849 28399 62883
rect 29377 62849 29411 62883
rect 29561 62849 29595 62883
rect 29929 62849 29963 62883
rect 29653 62781 29687 62815
rect 29745 62781 29779 62815
rect 1409 62645 1443 62679
rect 17233 62645 17267 62679
rect 19533 62645 19567 62679
rect 20545 62645 20579 62679
rect 23765 62645 23799 62679
rect 27169 62645 27203 62679
rect 23673 62441 23707 62475
rect 26893 62441 26927 62475
rect 29561 62441 29595 62475
rect 22477 62373 22511 62407
rect 21097 62305 21131 62339
rect 23305 62305 23339 62339
rect 16083 62237 16117 62271
rect 16221 62237 16255 62271
rect 16313 62237 16347 62271
rect 16497 62237 16531 62271
rect 17325 62237 17359 62271
rect 17581 62237 17615 62271
rect 23489 62237 23523 62271
rect 24685 62237 24719 62271
rect 24869 62237 24903 62271
rect 24961 62237 24995 62271
rect 27123 62237 27157 62271
rect 27261 62237 27295 62271
rect 27353 62237 27387 62271
rect 27537 62237 27571 62271
rect 29745 62237 29779 62271
rect 30021 62237 30055 62271
rect 14841 62169 14875 62203
rect 21364 62169 21398 62203
rect 28641 62169 28675 62203
rect 29929 62169 29963 62203
rect 14933 62101 14967 62135
rect 15853 62101 15887 62135
rect 18705 62101 18739 62135
rect 24501 62101 24535 62135
rect 28733 62101 28767 62135
rect 21833 61897 21867 61931
rect 24685 61897 24719 61931
rect 25053 61897 25087 61931
rect 25697 61897 25731 61931
rect 26985 61897 27019 61931
rect 12725 61829 12759 61863
rect 1593 61761 1627 61795
rect 12541 61761 12575 61795
rect 15209 61761 15243 61795
rect 15298 61761 15332 61795
rect 15393 61761 15427 61795
rect 15577 61761 15611 61795
rect 16681 61761 16715 61795
rect 18788 61761 18822 61795
rect 22109 61761 22143 61795
rect 22198 61761 22232 61795
rect 22298 61761 22332 61795
rect 22477 61761 22511 61795
rect 23305 61761 23339 61795
rect 23949 61761 23983 61795
rect 24133 61761 24167 61795
rect 24225 61761 24259 61795
rect 24869 61761 24903 61795
rect 25145 61761 25179 61795
rect 25881 61761 25915 61795
rect 26065 61761 26099 61795
rect 26157 61761 26191 61795
rect 27261 61761 27295 61795
rect 27353 61761 27387 61795
rect 27445 61761 27479 61795
rect 27629 61761 27663 61795
rect 28181 61761 28215 61795
rect 29193 61761 29227 61795
rect 16957 61693 16991 61727
rect 18521 61693 18555 61727
rect 28917 61693 28951 61727
rect 23765 61625 23799 61659
rect 1409 61557 1443 61591
rect 12909 61557 12943 61591
rect 14933 61557 14967 61591
rect 19901 61557 19935 61591
rect 23121 61557 23155 61591
rect 28365 61557 28399 61591
rect 16405 61353 16439 61387
rect 18705 61353 18739 61387
rect 27261 61353 27295 61387
rect 28549 61353 28583 61387
rect 29561 61353 29595 61387
rect 14473 61285 14507 61319
rect 25881 61217 25915 61251
rect 1593 61149 1627 61183
rect 12909 61149 12943 61183
rect 14289 61149 14323 61183
rect 17601 61149 17635 61183
rect 17706 61149 17740 61183
rect 17806 61146 17840 61180
rect 17969 61149 18003 61183
rect 18521 61149 18555 61183
rect 19717 61149 19751 61183
rect 23305 61149 23339 61183
rect 23489 61149 23523 61183
rect 24409 61149 24443 61183
rect 24685 61149 24719 61183
rect 26065 61149 26099 61183
rect 26341 61149 26375 61183
rect 27537 61149 27571 61183
rect 27629 61149 27663 61183
rect 27721 61149 27755 61183
rect 27905 61149 27939 61183
rect 28733 61149 28767 61183
rect 28917 61149 28951 61183
rect 29009 61149 29043 61183
rect 29745 61149 29779 61183
rect 30021 61149 30055 61183
rect 14105 61081 14139 61115
rect 15117 61081 15151 61115
rect 29929 61081 29963 61115
rect 1409 61013 1443 61047
rect 12725 61013 12759 61047
rect 17325 61013 17359 61047
rect 19809 61013 19843 61047
rect 23673 61013 23707 61047
rect 26249 61013 26283 61047
rect 18337 60809 18371 60843
rect 18889 60809 18923 60843
rect 26985 60809 27019 60843
rect 12541 60741 12575 60775
rect 25053 60741 25087 60775
rect 27353 60741 27387 60775
rect 29745 60741 29779 60775
rect 1593 60673 1627 60707
rect 12725 60673 12759 60707
rect 13645 60673 13679 60707
rect 13737 60673 13771 60707
rect 13829 60673 13863 60707
rect 14013 60673 14047 60707
rect 14729 60673 14763 60707
rect 17213 60673 17247 60707
rect 19165 60673 19199 60707
rect 19257 60673 19291 60707
rect 19349 60673 19383 60707
rect 19527 60673 19561 60707
rect 20867 60673 20901 60707
rect 21005 60673 21039 60707
rect 21097 60673 21131 60707
rect 21293 60673 21327 60707
rect 22845 60673 22879 60707
rect 23029 60673 23063 60707
rect 23949 60673 23983 60707
rect 24869 60673 24903 60707
rect 25145 60673 25179 60707
rect 25973 60673 26007 60707
rect 26157 60673 26191 60707
rect 26341 60673 26375 60707
rect 26433 60673 26467 60707
rect 27169 60673 27203 60707
rect 27445 60673 27479 60707
rect 28089 60673 28123 60707
rect 28917 60673 28951 60707
rect 14473 60605 14507 60639
rect 16957 60605 16991 60639
rect 23765 60605 23799 60639
rect 1409 60469 1443 60503
rect 12909 60469 12943 60503
rect 13369 60469 13403 60503
rect 15853 60469 15887 60503
rect 20637 60469 20671 60503
rect 23213 60469 23247 60503
rect 24133 60469 24167 60503
rect 24685 60469 24719 60503
rect 28181 60469 28215 60503
rect 29101 60469 29135 60503
rect 29837 60469 29871 60503
rect 17877 60265 17911 60299
rect 22385 60265 22419 60299
rect 25605 60265 25639 60299
rect 28549 60265 28583 60299
rect 14197 60197 14231 60231
rect 27445 60197 27479 60231
rect 12909 60129 12943 60163
rect 22937 60129 22971 60163
rect 28089 60129 28123 60163
rect 1593 60061 1627 60095
rect 12541 60061 12575 60095
rect 17693 60061 17727 60095
rect 19487 60061 19521 60095
rect 19625 60061 19659 60095
rect 19717 60061 19751 60095
rect 19901 60061 19935 60095
rect 21005 60061 21039 60095
rect 23121 60061 23155 60095
rect 25789 60061 25823 60095
rect 26065 60061 26099 60095
rect 26893 60061 26927 60095
rect 27813 60061 27847 60095
rect 27997 60061 28031 60095
rect 28181 60061 28215 60095
rect 28365 60061 28399 60095
rect 29837 60061 29871 60095
rect 12725 59993 12759 60027
rect 14473 59993 14507 60027
rect 14657 59993 14691 60027
rect 14749 59993 14783 60027
rect 15485 59993 15519 60027
rect 21250 59993 21284 60027
rect 25973 59993 26007 60027
rect 1409 59925 1443 59959
rect 16773 59925 16807 59959
rect 19257 59925 19291 59959
rect 23305 59925 23339 59959
rect 27077 59925 27111 59959
rect 30021 59925 30055 59959
rect 13553 59721 13587 59755
rect 14289 59721 14323 59755
rect 16865 59721 16899 59755
rect 23857 59721 23891 59755
rect 25789 59721 25823 59755
rect 27445 59721 27479 59755
rect 12541 59653 12575 59687
rect 12725 59653 12759 59687
rect 19524 59653 19558 59687
rect 1593 59585 1627 59619
rect 13461 59585 13495 59619
rect 14105 59585 14139 59619
rect 16681 59585 16715 59619
rect 19257 59585 19291 59619
rect 22937 59585 22971 59619
rect 23121 59585 23155 59619
rect 24041 59585 24075 59619
rect 25605 59585 25639 59619
rect 25881 59585 25915 59619
rect 27721 59585 27755 59619
rect 27813 59585 27847 59619
rect 27905 59585 27939 59619
rect 28089 59585 28123 59619
rect 28917 59585 28951 59619
rect 29745 59585 29779 59619
rect 20637 59449 20671 59483
rect 29101 59449 29135 59483
rect 1409 59381 1443 59415
rect 12909 59381 12943 59415
rect 23305 59381 23339 59415
rect 25421 59381 25455 59415
rect 29837 59381 29871 59415
rect 19809 59177 19843 59211
rect 20821 59177 20855 59211
rect 28733 59177 28767 59211
rect 13553 59109 13587 59143
rect 27169 59041 27203 59075
rect 13369 58973 13403 59007
rect 14657 58973 14691 59007
rect 20637 58973 20671 59007
rect 26893 58973 26927 59007
rect 13185 58905 13219 58939
rect 17877 58905 17911 58939
rect 19717 58905 19751 58939
rect 28641 58905 28675 58939
rect 29745 58905 29779 58939
rect 30113 58905 30147 58939
rect 14749 58837 14783 58871
rect 17969 58837 18003 58871
rect 19717 58633 19751 58667
rect 27445 58633 27479 58667
rect 30113 58633 30147 58667
rect 13369 58565 13403 58599
rect 15945 58565 15979 58599
rect 17233 58565 17267 58599
rect 19073 58565 19107 58599
rect 20821 58565 20855 58599
rect 26249 58565 26283 58599
rect 1409 58497 1443 58531
rect 13185 58497 13219 58531
rect 18889 58497 18923 58531
rect 19533 58497 19567 58531
rect 20637 58497 20671 58531
rect 26065 58497 26099 58531
rect 27721 58497 27755 58531
rect 27813 58503 27847 58537
rect 27905 58497 27939 58531
rect 28089 58497 28123 58531
rect 28641 58497 28675 58531
rect 29377 58497 29411 58531
rect 29561 58497 29595 58531
rect 29653 58497 29687 58531
rect 29929 58497 29963 58531
rect 17233 58429 17267 58463
rect 17325 58429 17359 58463
rect 29745 58429 29779 58463
rect 1593 58361 1627 58395
rect 16129 58361 16163 58395
rect 16773 58361 16807 58395
rect 28825 58361 28859 58395
rect 13553 58293 13587 58327
rect 17233 58089 17267 58123
rect 29561 58089 29595 58123
rect 26525 58021 26559 58055
rect 1409 57885 1443 57919
rect 15485 57885 15519 57919
rect 17509 57885 17543 57919
rect 20729 57885 20763 57919
rect 27077 57885 27111 57919
rect 28733 57885 28767 57919
rect 28917 57885 28951 57919
rect 29009 57885 29043 57919
rect 29745 57885 29779 57919
rect 30021 57885 30055 57919
rect 15301 57817 15335 57851
rect 16313 57817 16347 57851
rect 16589 57817 16623 57851
rect 17785 57817 17819 57851
rect 18429 57817 18463 57851
rect 26341 57817 26375 57851
rect 27905 57817 27939 57851
rect 1593 57749 1627 57783
rect 16019 57749 16053 57783
rect 16497 57749 16531 57783
rect 17693 57749 17727 57783
rect 18521 57749 18555 57783
rect 20913 57749 20947 57783
rect 27169 57749 27203 57783
rect 27997 57749 28031 57783
rect 28549 57749 28583 57783
rect 29929 57749 29963 57783
rect 2145 57545 2179 57579
rect 25881 57545 25915 57579
rect 29837 57545 29871 57579
rect 14924 57477 14958 57511
rect 26249 57477 26283 57511
rect 1409 57409 1443 57443
rect 2329 57409 2363 57443
rect 13783 57409 13817 57443
rect 13918 57412 13952 57446
rect 14013 57409 14047 57443
rect 14197 57409 14231 57443
rect 17049 57409 17083 57443
rect 19487 57409 19521 57443
rect 19625 57409 19659 57443
rect 19717 57409 19751 57443
rect 19901 57409 19935 57443
rect 20637 57409 20671 57443
rect 20729 57409 20763 57443
rect 20821 57409 20855 57443
rect 21005 57409 21039 57443
rect 22845 57409 22879 57443
rect 23029 57409 23063 57443
rect 23949 57409 23983 57443
rect 26065 57409 26099 57443
rect 26341 57409 26375 57443
rect 26985 57409 27019 57443
rect 29745 57409 29779 57443
rect 14657 57341 14691 57375
rect 28365 57341 28399 57375
rect 28641 57341 28675 57375
rect 23213 57273 23247 57307
rect 1593 57205 1627 57239
rect 13553 57205 13587 57239
rect 16037 57205 16071 57239
rect 18337 57205 18371 57239
rect 19257 57205 19291 57239
rect 20361 57205 20395 57239
rect 23765 57205 23799 57239
rect 27169 57205 27203 57239
rect 2145 57001 2179 57035
rect 16221 57001 16255 57035
rect 16773 57001 16807 57035
rect 25697 57001 25731 57035
rect 27721 57001 27755 57035
rect 28411 57001 28445 57035
rect 29745 57001 29779 57035
rect 13553 56933 13587 56967
rect 15485 56933 15519 56967
rect 14105 56865 14139 56899
rect 17233 56865 17267 56899
rect 17877 56865 17911 56899
rect 28181 56865 28215 56899
rect 1409 56797 1443 56831
rect 2329 56797 2363 56831
rect 13369 56797 13403 56831
rect 14361 56797 14395 56831
rect 16037 56797 16071 56831
rect 18153 56797 18187 56831
rect 19257 56797 19291 56831
rect 19524 56797 19558 56831
rect 21327 56797 21361 56831
rect 21465 56797 21499 56831
rect 21557 56797 21591 56831
rect 21741 56797 21775 56831
rect 22477 56797 22511 56831
rect 22566 56797 22600 56831
rect 22661 56797 22695 56831
rect 22857 56797 22891 56831
rect 24593 56797 24627 56831
rect 25881 56797 25915 56831
rect 26065 56797 26099 56831
rect 26157 56797 26191 56831
rect 26985 56797 27019 56831
rect 27169 56797 27203 56831
rect 27261 56797 27295 56831
rect 27353 56797 27387 56831
rect 27537 56797 27571 56831
rect 29745 56797 29779 56831
rect 17325 56729 17359 56763
rect 23397 56729 23431 56763
rect 24409 56729 24443 56763
rect 24961 56729 24995 56763
rect 1593 56661 1627 56695
rect 17233 56661 17267 56695
rect 20637 56661 20671 56695
rect 21097 56661 21131 56695
rect 22201 56661 22235 56695
rect 23489 56661 23523 56695
rect 24685 56661 24719 56695
rect 24777 56661 24811 56695
rect 2145 56457 2179 56491
rect 15393 56457 15427 56491
rect 23213 56457 23247 56491
rect 24409 56457 24443 56491
rect 24501 56457 24535 56491
rect 25789 56457 25823 56491
rect 28365 56457 28399 56491
rect 14473 56389 14507 56423
rect 17316 56389 17350 56423
rect 1409 56321 1443 56355
rect 2329 56321 2363 56355
rect 14565 56321 14599 56355
rect 15209 56321 15243 56355
rect 15945 56321 15979 56355
rect 18889 56321 18923 56355
rect 21833 56321 21867 56355
rect 22100 56321 22134 56355
rect 24317 56321 24351 56355
rect 24685 56321 24719 56355
rect 25973 56321 26007 56355
rect 26157 56321 26191 56355
rect 26249 56321 26283 56355
rect 27261 56321 27295 56355
rect 28549 56321 28583 56355
rect 28733 56321 28767 56355
rect 28825 56321 28859 56355
rect 29285 56321 29319 56355
rect 29561 56321 29595 56355
rect 14473 56253 14507 56287
rect 17049 56253 17083 56287
rect 26985 56253 27019 56287
rect 14013 56185 14047 56219
rect 24133 56185 24167 56219
rect 1593 56117 1627 56151
rect 16037 56117 16071 56151
rect 18429 56117 18463 56151
rect 20177 56117 20211 56151
rect 1685 55913 1719 55947
rect 21097 55913 21131 55947
rect 23213 55913 23247 55947
rect 24409 55913 24443 55947
rect 15853 55845 15887 55879
rect 16221 55777 16255 55811
rect 25053 55777 25087 55811
rect 27169 55777 27203 55811
rect 28181 55777 28215 55811
rect 1869 55709 1903 55743
rect 21833 55709 21867 55743
rect 22089 55709 22123 55743
rect 24593 55709 24627 55743
rect 24685 55709 24719 55743
rect 26893 55709 26927 55743
rect 28457 55709 28491 55743
rect 16405 55641 16439 55675
rect 16957 55641 16991 55675
rect 19625 55641 19659 55675
rect 25513 55641 25547 55675
rect 25697 55641 25731 55675
rect 26065 55641 26099 55675
rect 29745 55641 29779 55675
rect 30113 55641 30147 55675
rect 16313 55573 16347 55607
rect 18245 55573 18279 55607
rect 24777 55573 24811 55607
rect 24961 55573 24995 55607
rect 25789 55573 25823 55607
rect 25881 55573 25915 55607
rect 2145 55369 2179 55403
rect 17325 55369 17359 55403
rect 18061 55369 18095 55403
rect 20821 55369 20855 55403
rect 24593 55369 24627 55403
rect 25329 55369 25363 55403
rect 25789 55369 25823 55403
rect 26985 55369 27019 55403
rect 30113 55369 30147 55403
rect 16129 55301 16163 55335
rect 25881 55301 25915 55335
rect 27353 55301 27387 55335
rect 1409 55233 1443 55267
rect 2329 55233 2363 55267
rect 15945 55233 15979 55267
rect 17233 55233 17267 55267
rect 17877 55233 17911 55267
rect 19809 55233 19843 55267
rect 19901 55233 19935 55267
rect 19993 55233 20027 55267
rect 20177 55233 20211 55267
rect 20729 55233 20763 55267
rect 22477 55233 22511 55267
rect 23581 55233 23615 55267
rect 23673 55233 23707 55267
rect 24225 55233 24259 55267
rect 24409 55233 24443 55267
rect 25513 55233 25547 55267
rect 27169 55233 27203 55267
rect 27445 55233 27479 55267
rect 28181 55233 28215 55267
rect 28365 55233 28399 55267
rect 28733 55233 28767 55267
rect 29377 55233 29411 55267
rect 29561 55233 29595 55267
rect 29653 55233 29687 55267
rect 29929 55233 29963 55267
rect 22293 55165 22327 55199
rect 22661 55165 22695 55199
rect 23397 55165 23431 55199
rect 23489 55165 23523 55199
rect 24501 55165 24535 55199
rect 24777 55165 24811 55199
rect 24869 55165 24903 55199
rect 25605 55165 25639 55199
rect 25973 55165 26007 55199
rect 28457 55165 28491 55199
rect 28549 55165 28583 55199
rect 29745 55165 29779 55199
rect 1593 55097 1627 55131
rect 28917 55097 28951 55131
rect 19533 55029 19567 55063
rect 23213 55029 23247 55063
rect 15853 54825 15887 54859
rect 24639 54825 24673 54859
rect 25973 54825 26007 54859
rect 27905 54825 27939 54859
rect 28825 54757 28859 54791
rect 24409 54689 24443 54723
rect 30021 54689 30055 54723
rect 1409 54621 1443 54655
rect 15669 54621 15703 54655
rect 16313 54621 16347 54655
rect 26157 54621 26191 54655
rect 26433 54621 26467 54655
rect 27537 54621 27571 54655
rect 29745 54621 29779 54655
rect 22109 54553 22143 54587
rect 27721 54553 27755 54587
rect 28641 54553 28675 54587
rect 1593 54485 1627 54519
rect 16497 54485 16531 54519
rect 23397 54485 23431 54519
rect 26341 54485 26375 54519
rect 2145 54281 2179 54315
rect 18061 54281 18095 54315
rect 21097 54281 21131 54315
rect 30113 54281 30147 54315
rect 16926 54213 16960 54247
rect 28457 54213 28491 54247
rect 1409 54145 1443 54179
rect 2329 54145 2363 54179
rect 16681 54145 16715 54179
rect 19973 54145 20007 54179
rect 23121 54145 23155 54179
rect 23305 54145 23339 54179
rect 25237 54145 25271 54179
rect 27537 54145 27571 54179
rect 27721 54145 27755 54179
rect 29377 54145 29411 54179
rect 29561 54145 29595 54179
rect 29745 54145 29779 54179
rect 29929 54145 29963 54179
rect 19717 54077 19751 54111
rect 29653 54077 29687 54111
rect 28641 54009 28675 54043
rect 1593 53941 1627 53975
rect 23489 53941 23523 53975
rect 25329 53941 25363 53975
rect 27629 53941 27663 53975
rect 2145 53737 2179 53771
rect 18061 53737 18095 53771
rect 18705 53737 18739 53771
rect 19441 53737 19475 53771
rect 30021 53737 30055 53771
rect 1409 53533 1443 53567
rect 2329 53533 2363 53567
rect 17877 53533 17911 53567
rect 18521 53533 18555 53567
rect 19993 53533 20027 53567
rect 22385 53533 22419 53567
rect 25789 53533 25823 53567
rect 26709 53533 26743 53567
rect 26893 53533 26927 53567
rect 26985 53533 27019 53567
rect 27997 53533 28031 53567
rect 28733 53533 28767 53567
rect 29745 53533 29779 53567
rect 19349 53465 19383 53499
rect 1593 53397 1627 53431
rect 21281 53397 21315 53431
rect 22477 53397 22511 53431
rect 25973 53397 26007 53431
rect 26525 53397 26559 53431
rect 28181 53397 28215 53431
rect 28917 53397 28951 53431
rect 1685 53193 1719 53227
rect 17785 53193 17819 53227
rect 18521 53193 18555 53227
rect 19901 53193 19935 53227
rect 21281 53193 21315 53227
rect 27445 53193 27479 53227
rect 29285 53193 29319 53227
rect 17693 53125 17727 53159
rect 19073 53125 19107 53159
rect 21925 53125 21959 53159
rect 26341 53125 26375 53159
rect 1869 53057 1903 53091
rect 14188 53057 14222 53091
rect 18337 53057 18371 53091
rect 19717 53057 19751 53091
rect 21097 53057 21131 53091
rect 22569 53057 22603 53091
rect 23581 53057 23615 53091
rect 26157 53057 26191 53091
rect 26433 53057 26467 53091
rect 27721 53057 27755 53091
rect 27813 53057 27847 53091
rect 27905 53057 27939 53091
rect 28089 53057 28123 53091
rect 28549 53057 28583 53091
rect 28733 53057 28767 53091
rect 28917 53057 28951 53091
rect 29101 53057 29135 53091
rect 29837 53057 29871 53091
rect 13921 52989 13955 53023
rect 28825 52989 28859 53023
rect 19257 52921 19291 52955
rect 22661 52921 22695 52955
rect 25973 52921 26007 52955
rect 15301 52853 15335 52887
rect 22017 52853 22051 52887
rect 23673 52853 23707 52887
rect 30021 52853 30055 52887
rect 13369 52649 13403 52683
rect 15393 52649 15427 52683
rect 17693 52649 17727 52683
rect 19349 52649 19383 52683
rect 20729 52649 20763 52683
rect 23305 52649 23339 52683
rect 27169 52649 27203 52683
rect 29837 52649 29871 52683
rect 1409 52581 1443 52615
rect 2053 52581 2087 52615
rect 14105 52581 14139 52615
rect 19809 52513 19843 52547
rect 21925 52513 21959 52547
rect 26249 52513 26283 52547
rect 28549 52513 28583 52547
rect 1593 52445 1627 52479
rect 2237 52445 2271 52479
rect 11805 52445 11839 52479
rect 12081 52445 12115 52479
rect 14381 52445 14415 52479
rect 14473 52445 14507 52479
rect 14565 52445 14599 52479
rect 14749 52445 14783 52479
rect 15209 52445 15243 52479
rect 17141 52445 17175 52479
rect 17969 52445 18003 52479
rect 18245 52445 18279 52479
rect 26433 52445 26467 52479
rect 26709 52445 26743 52479
rect 27445 52445 27479 52479
rect 27537 52442 27571 52476
rect 27629 52445 27663 52479
rect 27813 52445 27847 52479
rect 28273 52445 28307 52479
rect 28457 52445 28491 52479
rect 28641 52445 28675 52479
rect 28825 52445 28859 52479
rect 16957 52377 16991 52411
rect 18153 52377 18187 52411
rect 19901 52377 19935 52411
rect 20637 52377 20671 52411
rect 22192 52377 22226 52411
rect 26617 52377 26651 52411
rect 29745 52377 29779 52411
rect 19809 52309 19843 52343
rect 29009 52309 29043 52343
rect 1869 52105 1903 52139
rect 11713 52105 11747 52139
rect 17233 52105 17267 52139
rect 18245 52105 18279 52139
rect 22385 52105 22419 52139
rect 25881 52105 25915 52139
rect 25973 52105 26007 52139
rect 27077 52105 27111 52139
rect 30113 52105 30147 52139
rect 14289 52037 14323 52071
rect 18061 52037 18095 52071
rect 21907 52037 21941 52071
rect 26157 52037 26191 52071
rect 1685 51969 1719 52003
rect 11529 51969 11563 52003
rect 15005 51969 15039 52003
rect 17049 51969 17083 52003
rect 18889 51969 18923 52003
rect 20637 51969 20671 52003
rect 23305 51969 23339 52003
rect 25789 51969 25823 52003
rect 27353 51969 27387 52003
rect 27445 51969 27479 52003
rect 27537 51969 27571 52003
rect 27721 51969 27755 52003
rect 28181 51969 28215 52003
rect 28365 51969 28399 52003
rect 28733 51969 28767 52003
rect 29377 51969 29411 52003
rect 29561 51969 29595 52003
rect 29929 51969 29963 52003
rect 12633 51901 12667 51935
rect 12909 51901 12943 51935
rect 14749 51901 14783 51935
rect 18337 51901 18371 51935
rect 22293 51901 22327 51935
rect 22477 51901 22511 51935
rect 23581 51901 23615 51935
rect 28457 51901 28491 51935
rect 28549 51901 28583 51935
rect 29653 51901 29687 51935
rect 29745 51901 29779 51935
rect 17785 51833 17819 51867
rect 25605 51833 25639 51867
rect 16129 51765 16163 51799
rect 28917 51765 28951 51799
rect 13001 51561 13035 51595
rect 14473 51561 14507 51595
rect 15761 51561 15795 51595
rect 17969 51561 18003 51595
rect 19349 51561 19383 51595
rect 20545 51561 20579 51595
rect 22293 51561 22327 51595
rect 18705 51425 18739 51459
rect 19901 51425 19935 51459
rect 21097 51425 21131 51459
rect 25605 51425 25639 51459
rect 1593 51357 1627 51391
rect 2237 51357 2271 51391
rect 12817 51357 12851 51391
rect 14749 51357 14783 51391
rect 14841 51357 14875 51391
rect 14933 51357 14967 51391
rect 15117 51357 15151 51391
rect 15577 51357 15611 51391
rect 17785 51357 17819 51391
rect 19625 51357 19659 51391
rect 20821 51357 20855 51391
rect 22477 51357 22511 51391
rect 22569 51357 22603 51391
rect 22753 51357 22787 51391
rect 22845 51357 22879 51391
rect 24593 51357 24627 51391
rect 28733 51357 28767 51391
rect 18521 51289 18555 51323
rect 19809 51289 19843 51323
rect 24409 51289 24443 51323
rect 24961 51289 24995 51323
rect 25789 51289 25823 51323
rect 26157 51289 26191 51323
rect 29745 51289 29779 51323
rect 1409 51221 1443 51255
rect 2053 51221 2087 51255
rect 21005 51221 21039 51255
rect 24685 51221 24719 51255
rect 24777 51221 24811 51255
rect 25881 51221 25915 51255
rect 25973 51221 26007 51255
rect 28917 51221 28951 51255
rect 29837 51221 29871 51255
rect 17509 51017 17543 51051
rect 22661 51017 22695 51051
rect 24501 51017 24535 51051
rect 24685 51017 24719 51051
rect 25513 51017 25547 51051
rect 25605 51017 25639 51051
rect 20085 50949 20119 50983
rect 22109 50949 22143 50983
rect 1593 50881 1627 50915
rect 14933 50881 14967 50915
rect 15025 50881 15059 50915
rect 15117 50881 15151 50915
rect 15301 50881 15335 50915
rect 17325 50881 17359 50915
rect 21925 50881 21959 50915
rect 22569 50881 22603 50915
rect 24317 50881 24351 50915
rect 25421 50881 25455 50915
rect 25789 50881 25823 50915
rect 28917 50881 28951 50915
rect 29745 50881 29779 50915
rect 24409 50813 24443 50847
rect 24777 50813 24811 50847
rect 25237 50745 25271 50779
rect 1409 50677 1443 50711
rect 14657 50677 14691 50711
rect 20177 50677 20211 50711
rect 24133 50677 24167 50711
rect 29101 50677 29135 50711
rect 29837 50677 29871 50711
rect 2697 50473 2731 50507
rect 19901 50473 19935 50507
rect 21741 50473 21775 50507
rect 24409 50405 24443 50439
rect 1777 50269 1811 50303
rect 2605 50269 2639 50303
rect 11805 50269 11839 50303
rect 15577 50269 15611 50303
rect 15844 50269 15878 50303
rect 19717 50269 19751 50303
rect 20361 50269 20395 50303
rect 22477 50269 22511 50303
rect 22569 50269 22603 50303
rect 22661 50269 22695 50303
rect 22845 50269 22879 50303
rect 23489 50269 23523 50303
rect 23857 50269 23891 50303
rect 24593 50269 24627 50303
rect 24817 50269 24851 50303
rect 27997 50269 28031 50303
rect 1593 50201 1627 50235
rect 1961 50201 1995 50235
rect 2421 50201 2455 50235
rect 12072 50201 12106 50235
rect 20628 50201 20662 50235
rect 22201 50201 22235 50235
rect 24961 50201 24995 50235
rect 28825 50201 28859 50235
rect 29009 50201 29043 50235
rect 29745 50201 29779 50235
rect 13185 50133 13219 50167
rect 16957 50133 16991 50167
rect 23397 50133 23431 50167
rect 23581 50133 23615 50167
rect 23673 50133 23707 50167
rect 24685 50133 24719 50167
rect 28181 50133 28215 50167
rect 29837 50133 29871 50167
rect 11897 49929 11931 49963
rect 15669 49929 15703 49963
rect 19993 49929 20027 49963
rect 23029 49929 23063 49963
rect 23765 49929 23799 49963
rect 24225 49929 24259 49963
rect 24869 49929 24903 49963
rect 25329 49929 25363 49963
rect 1593 49861 1627 49895
rect 1777 49861 1811 49895
rect 28733 49861 28767 49895
rect 29745 49861 29779 49895
rect 29929 49861 29963 49895
rect 2605 49793 2639 49827
rect 11713 49793 11747 49827
rect 13001 49793 13035 49827
rect 15485 49793 15519 49827
rect 19809 49793 19843 49827
rect 20453 49793 20487 49827
rect 22385 49793 22419 49827
rect 24409 49793 24443 49827
rect 25421 49793 25455 49827
rect 28825 49793 28859 49827
rect 1961 49725 1995 49759
rect 13277 49725 13311 49759
rect 14381 49725 14415 49759
rect 23949 49725 23983 49759
rect 24041 49725 24075 49759
rect 24317 49725 24351 49759
rect 25053 49725 25087 49759
rect 25145 49725 25179 49759
rect 25513 49725 25547 49759
rect 28733 49725 28767 49759
rect 30021 49725 30055 49759
rect 28273 49657 28307 49691
rect 29469 49657 29503 49691
rect 2421 49589 2455 49623
rect 20637 49589 20671 49623
rect 1961 49385 1995 49419
rect 14289 49385 14323 49419
rect 19625 49385 19659 49419
rect 21833 49385 21867 49419
rect 25421 49385 25455 49419
rect 26709 49385 26743 49419
rect 27629 49385 27663 49419
rect 23213 49317 23247 49351
rect 2789 49249 2823 49283
rect 12449 49249 12483 49283
rect 13369 49249 13403 49283
rect 20085 49249 20119 49283
rect 21005 49249 21039 49283
rect 25605 49249 25639 49283
rect 26065 49249 26099 49283
rect 1593 49181 1627 49215
rect 1777 49181 1811 49215
rect 9965 49181 9999 49215
rect 14105 49181 14139 49215
rect 22017 49181 22051 49215
rect 22293 49181 22327 49215
rect 23029 49181 23063 49215
rect 25697 49181 25731 49215
rect 26893 49181 26927 49215
rect 27169 49181 27203 49215
rect 27813 49181 27847 49215
rect 28089 49181 28123 49215
rect 28641 49181 28675 49215
rect 2421 49113 2455 49147
rect 2605 49113 2639 49147
rect 10210 49113 10244 49147
rect 12541 49113 12575 49147
rect 13185 49113 13219 49147
rect 20177 49113 20211 49147
rect 20821 49113 20855 49147
rect 22201 49113 22235 49147
rect 27077 49113 27111 49147
rect 29745 49113 29779 49147
rect 30113 49113 30147 49147
rect 11345 49045 11379 49079
rect 11971 49045 12005 49079
rect 12449 49045 12483 49079
rect 20085 49045 20119 49079
rect 25789 49045 25823 49079
rect 25973 49045 26007 49079
rect 27997 49045 28031 49079
rect 28917 49045 28951 49079
rect 3249 48841 3283 48875
rect 10425 48841 10459 48875
rect 23581 48841 23615 48875
rect 24317 48841 24351 48875
rect 25145 48841 25179 48875
rect 25697 48841 25731 48875
rect 26065 48841 26099 48875
rect 27169 48841 27203 48875
rect 27537 48841 27571 48875
rect 28641 48841 28675 48875
rect 1593 48773 1627 48807
rect 1777 48773 1811 48807
rect 2789 48773 2823 48807
rect 12081 48773 12115 48807
rect 19809 48773 19843 48807
rect 19993 48773 20027 48807
rect 20729 48773 20763 48807
rect 29929 48773 29963 48807
rect 2421 48705 2455 48739
rect 2605 48705 2639 48739
rect 3433 48705 3467 48739
rect 10241 48705 10275 48739
rect 14565 48705 14599 48739
rect 17397 48705 17431 48739
rect 17506 48705 17540 48739
rect 17601 48705 17635 48739
rect 17785 48705 17819 48739
rect 22569 48705 22603 48739
rect 22845 48705 22879 48739
rect 23397 48705 23431 48739
rect 24225 48705 24259 48739
rect 25053 48705 25087 48739
rect 25973 48705 26007 48739
rect 27353 48705 27387 48739
rect 27629 48705 27663 48739
rect 28549 48705 28583 48739
rect 29745 48705 29779 48739
rect 12081 48637 12115 48671
rect 12173 48637 12207 48671
rect 20085 48637 20119 48671
rect 25881 48637 25915 48671
rect 26249 48637 26283 48671
rect 26341 48637 26375 48671
rect 28825 48637 28859 48671
rect 30021 48637 30055 48671
rect 11621 48569 11655 48603
rect 14749 48569 14783 48603
rect 19533 48569 19567 48603
rect 22661 48569 22695 48603
rect 22753 48569 22787 48603
rect 1961 48501 1995 48535
rect 17141 48501 17175 48535
rect 20821 48501 20855 48535
rect 22385 48501 22419 48535
rect 28181 48501 28215 48535
rect 29469 48501 29503 48535
rect 1685 48297 1719 48331
rect 18521 48297 18555 48331
rect 2697 48229 2731 48263
rect 11897 48229 11931 48263
rect 20545 48229 20579 48263
rect 21925 48229 21959 48263
rect 25697 48229 25731 48263
rect 27077 48229 27111 48263
rect 28549 48229 28583 48263
rect 29561 48229 29595 48263
rect 26249 48161 26283 48195
rect 1869 48093 1903 48127
rect 12173 48093 12207 48127
rect 14565 48093 14599 48127
rect 14657 48093 14691 48127
rect 14749 48093 14783 48127
rect 14933 48093 14967 48127
rect 17141 48093 17175 48127
rect 19257 48093 19291 48127
rect 20361 48093 20395 48127
rect 21189 48093 21223 48127
rect 21833 48093 21867 48127
rect 25881 48093 25915 48127
rect 25973 48093 26007 48127
rect 26111 48093 26145 48127
rect 26341 48093 26375 48127
rect 27261 48093 27295 48127
rect 27537 48093 27571 48127
rect 28733 48093 28767 48127
rect 29009 48093 29043 48127
rect 29745 48093 29779 48127
rect 30021 48093 30055 48127
rect 2329 48025 2363 48059
rect 2513 48025 2547 48059
rect 12449 48025 12483 48059
rect 13369 48025 13403 48059
rect 16129 48025 16163 48059
rect 17408 48025 17442 48059
rect 21373 48025 21407 48059
rect 27445 48025 27479 48059
rect 12357 47957 12391 47991
rect 13461 47957 13495 47991
rect 14289 47957 14323 47991
rect 16221 47957 16255 47991
rect 19441 47957 19475 47991
rect 28917 47957 28951 47991
rect 29929 47957 29963 47991
rect 1409 47753 1443 47787
rect 2053 47753 2087 47787
rect 13921 47753 13955 47787
rect 15117 47753 15151 47787
rect 16037 47753 16071 47787
rect 18521 47753 18555 47787
rect 25973 47753 26007 47787
rect 14933 47685 14967 47719
rect 29929 47685 29963 47719
rect 30021 47685 30055 47719
rect 1593 47617 1627 47651
rect 2237 47617 2271 47651
rect 15945 47617 15979 47651
rect 17509 47617 17543 47651
rect 17601 47617 17635 47651
rect 17714 47623 17748 47657
rect 17877 47617 17911 47651
rect 18337 47617 18371 47651
rect 18981 47617 19015 47651
rect 20269 47617 20303 47651
rect 26157 47617 26191 47651
rect 26341 47617 26375 47651
rect 26433 47617 26467 47651
rect 13921 47549 13955 47583
rect 14013 47549 14047 47583
rect 15209 47549 15243 47583
rect 17233 47549 17267 47583
rect 27445 47549 27479 47583
rect 27721 47549 27755 47583
rect 29837 47549 29871 47583
rect 13461 47481 13495 47515
rect 14657 47481 14691 47515
rect 29469 47481 29503 47515
rect 19165 47413 19199 47447
rect 20453 47413 20487 47447
rect 18705 47209 18739 47243
rect 23489 47209 23523 47243
rect 24961 47209 24995 47243
rect 26525 47209 26559 47243
rect 16865 47141 16899 47175
rect 19441 47141 19475 47175
rect 22937 47141 22971 47175
rect 17325 47073 17359 47107
rect 27445 47073 27479 47107
rect 27721 47073 27755 47107
rect 1593 47005 1627 47039
rect 2605 47005 2639 47039
rect 13369 47005 13403 47039
rect 14657 47005 14691 47039
rect 14924 47005 14958 47039
rect 16681 47005 16715 47039
rect 19257 47005 19291 47039
rect 19901 47005 19935 47039
rect 22293 47005 22327 47039
rect 22477 47005 22511 47039
rect 23213 47005 23247 47039
rect 26709 47005 26743 47039
rect 26985 47005 27019 47039
rect 28733 47005 28767 47039
rect 13553 46937 13587 46971
rect 17570 46937 17604 46971
rect 20637 46937 20671 46971
rect 20821 46937 20855 46971
rect 24869 46937 24903 46971
rect 26893 46937 26927 46971
rect 29745 46937 29779 46971
rect 30113 46937 30147 46971
rect 1409 46869 1443 46903
rect 2421 46869 2455 46903
rect 16037 46869 16071 46903
rect 20085 46869 20119 46903
rect 22385 46869 22419 46903
rect 23121 46869 23155 46903
rect 23305 46869 23339 46903
rect 28917 46869 28951 46903
rect 13185 46665 13219 46699
rect 19073 46665 19107 46699
rect 25237 46665 25271 46699
rect 25697 46665 25731 46699
rect 14473 46597 14507 46631
rect 14657 46597 14691 46631
rect 15945 46597 15979 46631
rect 17233 46597 17267 46631
rect 18153 46597 18187 46631
rect 19533 46597 19567 46631
rect 21281 46597 21315 46631
rect 1593 46529 1627 46563
rect 11897 46529 11931 46563
rect 15761 46529 15795 46563
rect 17049 46529 17083 46563
rect 17969 46529 18003 46563
rect 18889 46529 18923 46563
rect 22017 46529 22051 46563
rect 22109 46529 22143 46563
rect 23305 46529 23339 46563
rect 23489 46529 23523 46563
rect 28917 46529 28951 46563
rect 29745 46529 29779 46563
rect 14749 46461 14783 46495
rect 16037 46461 16071 46495
rect 17325 46461 17359 46495
rect 22293 46461 22327 46495
rect 25421 46461 25455 46495
rect 25513 46461 25547 46495
rect 25789 46461 25823 46495
rect 25881 46461 25915 46495
rect 14197 46393 14231 46427
rect 15485 46393 15519 46427
rect 16773 46393 16807 46427
rect 1409 46325 1443 46359
rect 22201 46325 22235 46359
rect 23397 46325 23431 46359
rect 29101 46325 29135 46359
rect 30021 46325 30055 46359
rect 12725 46121 12759 46155
rect 14657 46121 14691 46155
rect 19993 46121 20027 46155
rect 22293 46121 22327 46155
rect 29561 46121 29595 46155
rect 11621 46053 11655 46087
rect 17049 46053 17083 46087
rect 22753 46053 22787 46087
rect 12081 45985 12115 46019
rect 18245 45985 18279 46019
rect 20913 45985 20947 46019
rect 23305 45985 23339 46019
rect 25789 45985 25823 46019
rect 1593 45917 1627 45951
rect 2513 45917 2547 45951
rect 10333 45917 10367 45951
rect 13001 45917 13035 45951
rect 13093 45917 13127 45951
rect 13185 45917 13219 45951
rect 13369 45917 13403 45951
rect 14473 45917 14507 45951
rect 15117 45917 15151 45951
rect 21180 45917 21214 45951
rect 23029 45917 23063 45951
rect 25513 45917 25547 45951
rect 29745 45917 29779 45951
rect 30021 45917 30055 45951
rect 2329 45849 2363 45883
rect 12173 45849 12207 45883
rect 15761 45849 15795 45883
rect 18061 45849 18095 45883
rect 19901 45849 19935 45883
rect 24869 45849 24903 45883
rect 1409 45781 1443 45815
rect 2697 45781 2731 45815
rect 10517 45781 10551 45815
rect 12081 45781 12115 45815
rect 15301 45781 15335 45815
rect 22937 45781 22971 45815
rect 23121 45781 23155 45815
rect 24961 45781 24995 45815
rect 29929 45781 29963 45815
rect 16129 45577 16163 45611
rect 24317 45577 24351 45611
rect 25421 45577 25455 45611
rect 29193 45577 29227 45611
rect 2329 45509 2363 45543
rect 2513 45509 2547 45543
rect 12541 45509 12575 45543
rect 17049 45509 17083 45543
rect 18613 45509 18647 45543
rect 20453 45509 20487 45543
rect 24409 45509 24443 45543
rect 28641 45509 28675 45543
rect 1593 45441 1627 45475
rect 12771 45441 12805 45475
rect 12909 45441 12943 45475
rect 13022 45441 13056 45475
rect 13185 45441 13219 45475
rect 13737 45441 13771 45475
rect 15945 45441 15979 45475
rect 19257 45441 19291 45475
rect 20269 45441 20303 45475
rect 21097 45441 21131 45475
rect 21925 45441 21959 45475
rect 24133 45441 24167 45475
rect 25605 45441 25639 45475
rect 28457 45441 28491 45475
rect 28733 45441 28767 45475
rect 29377 45441 29411 45475
rect 29561 45441 29595 45475
rect 29653 45441 29687 45475
rect 20545 45373 20579 45407
rect 22109 45373 22143 45407
rect 24041 45373 24075 45407
rect 24501 45373 24535 45407
rect 25145 45373 25179 45407
rect 25237 45373 25271 45407
rect 25513 45373 25547 45407
rect 15025 45305 15059 45339
rect 19993 45305 20027 45339
rect 1409 45237 1443 45271
rect 2697 45237 2731 45271
rect 19441 45237 19475 45271
rect 21189 45237 21223 45271
rect 23857 45237 23891 45271
rect 24961 45237 24995 45271
rect 28273 45237 28307 45271
rect 1961 45033 1995 45067
rect 11989 45033 12023 45067
rect 18245 45033 18279 45067
rect 20545 45033 20579 45067
rect 29561 45033 29595 45067
rect 19349 44965 19383 44999
rect 28089 44965 28123 44999
rect 10057 44897 10091 44931
rect 19809 44897 19843 44931
rect 21005 44897 21039 44931
rect 21097 44897 21131 44931
rect 25053 44897 25087 44931
rect 25421 44897 25455 44931
rect 1777 44829 1811 44863
rect 12219 44829 12253 44863
rect 12357 44829 12391 44863
rect 12449 44829 12483 44863
rect 12645 44829 12679 44863
rect 13369 44829 13403 44863
rect 21925 44829 21959 44863
rect 22192 44829 22226 44863
rect 25145 44829 25179 44863
rect 25513 44829 25547 44863
rect 27169 44829 27203 44863
rect 28273 44829 28307 44863
rect 28733 44829 28767 44863
rect 29745 44829 29779 44863
rect 30021 44829 30055 44863
rect 1593 44761 1627 44795
rect 10302 44761 10336 44795
rect 14473 44761 14507 44795
rect 16957 44761 16991 44795
rect 19901 44761 19935 44795
rect 11437 44693 11471 44727
rect 13461 44693 13495 44727
rect 15761 44693 15795 44727
rect 19809 44693 19843 44727
rect 21005 44693 21039 44727
rect 23305 44693 23339 44727
rect 24869 44693 24903 44727
rect 25237 44693 25271 44727
rect 27353 44693 27387 44727
rect 28917 44693 28951 44727
rect 29929 44693 29963 44727
rect 2421 44489 2455 44523
rect 13093 44489 13127 44523
rect 15945 44489 15979 44523
rect 16763 44489 16797 44523
rect 20821 44489 20855 44523
rect 24501 44489 24535 44523
rect 29285 44489 29319 44523
rect 1593 44421 1627 44455
rect 1777 44421 1811 44455
rect 10793 44421 10827 44455
rect 10977 44421 11011 44455
rect 13001 44421 13035 44455
rect 14197 44421 14231 44455
rect 15761 44421 15795 44455
rect 16037 44421 16071 44455
rect 17233 44421 17267 44455
rect 19533 44421 19567 44455
rect 21925 44421 21959 44455
rect 24409 44421 24443 44455
rect 27629 44421 27663 44455
rect 2605 44353 2639 44387
rect 12081 44353 12115 44387
rect 12170 44353 12204 44387
rect 12265 44353 12299 44387
rect 12449 44353 12483 44387
rect 14013 44353 14047 44387
rect 14749 44353 14783 44387
rect 14933 44353 14967 44387
rect 17325 44353 17359 44387
rect 18153 44353 18187 44387
rect 18245 44353 18279 44387
rect 18337 44353 18371 44387
rect 18521 44353 18555 44387
rect 22661 44353 22695 44387
rect 23489 44353 23523 44387
rect 23673 44353 23707 44387
rect 25605 44353 25639 44387
rect 27813 44353 27847 44387
rect 27997 44353 28031 44387
rect 28089 44353 28123 44387
rect 29101 44353 29135 44387
rect 29837 44353 29871 44387
rect 11805 44285 11839 44319
rect 17141 44285 17175 44319
rect 23857 44285 23891 44319
rect 25881 44285 25915 44319
rect 1961 44217 1995 44251
rect 15485 44217 15519 44251
rect 30021 44217 30055 44251
rect 17877 44149 17911 44183
rect 22017 44149 22051 44183
rect 22845 44149 22879 44183
rect 2789 43945 2823 43979
rect 13553 43945 13587 43979
rect 15393 43945 15427 43979
rect 17877 43945 17911 43979
rect 22661 43945 22695 43979
rect 23397 43945 23431 43979
rect 26893 43945 26927 43979
rect 10885 43877 10919 43911
rect 14197 43877 14231 43911
rect 19349 43877 19383 43911
rect 20545 43877 20579 43911
rect 11345 43809 11379 43843
rect 14749 43809 14783 43843
rect 15853 43809 15887 43843
rect 19809 43809 19843 43843
rect 21005 43809 21039 43843
rect 23581 43809 23615 43843
rect 24685 43809 24719 43843
rect 28273 43809 28307 43843
rect 1777 43741 1811 43775
rect 9945 43741 9979 43775
rect 10054 43738 10088 43772
rect 10149 43738 10183 43772
rect 10333 43741 10367 43775
rect 12521 43741 12555 43775
rect 12614 43741 12648 43775
rect 12725 43741 12759 43775
rect 12909 43741 12943 43775
rect 13369 43741 13403 43775
rect 15945 43741 15979 43775
rect 19901 43741 19935 43775
rect 21097 43741 21131 43775
rect 22017 43741 22051 43775
rect 22477 43741 22511 43775
rect 23765 43741 23799 43775
rect 23857 43741 23891 43775
rect 24593 43741 24627 43775
rect 25053 43741 25087 43775
rect 27077 43741 27111 43775
rect 27353 43741 27387 43775
rect 27997 43741 28031 43775
rect 29837 43741 29871 43775
rect 1593 43673 1627 43707
rect 2421 43673 2455 43707
rect 2605 43673 2639 43707
rect 9689 43673 9723 43707
rect 11437 43673 11471 43707
rect 14473 43673 14507 43707
rect 14657 43673 14691 43707
rect 15853 43673 15887 43707
rect 16589 43673 16623 43707
rect 1961 43605 1995 43639
rect 11345 43605 11379 43639
rect 12265 43605 12299 43639
rect 19809 43605 19843 43639
rect 21005 43605 21039 43639
rect 21833 43605 21867 43639
rect 24409 43605 24443 43639
rect 24777 43605 24811 43639
rect 24961 43605 24995 43639
rect 27261 43605 27295 43639
rect 30021 43605 30055 43639
rect 2421 43401 2455 43435
rect 9597 43401 9631 43435
rect 18337 43401 18371 43435
rect 20821 43401 20855 43435
rect 23673 43401 23707 43435
rect 1593 43333 1627 43367
rect 15945 43333 15979 43367
rect 19533 43333 19567 43367
rect 22293 43333 22327 43367
rect 23765 43333 23799 43367
rect 30113 43333 30147 43367
rect 1777 43265 1811 43299
rect 2605 43265 2639 43299
rect 9853 43265 9887 43299
rect 9962 43271 9996 43305
rect 10057 43265 10091 43299
rect 10241 43265 10275 43299
rect 11805 43265 11839 43299
rect 13093 43265 13127 43299
rect 15025 43265 15059 43299
rect 15761 43265 15795 43299
rect 17049 43265 17083 43299
rect 23489 43265 23523 43299
rect 23857 43265 23891 43299
rect 24593 43265 24627 43299
rect 25789 43265 25823 43299
rect 27997 43265 28031 43299
rect 28641 43265 28675 43299
rect 29101 43265 29135 43299
rect 29929 43265 29963 43299
rect 11529 43197 11563 43231
rect 12817 43197 12851 43231
rect 23397 43197 23431 43231
rect 24317 43197 24351 43231
rect 25973 43197 26007 43231
rect 1961 43129 1995 43163
rect 15209 43129 15243 43163
rect 14381 43061 14415 43095
rect 22385 43061 22419 43095
rect 23213 43061 23247 43095
rect 27813 43061 27847 43095
rect 28457 43061 28491 43095
rect 29285 43061 29319 43095
rect 1409 42857 1443 42891
rect 2053 42857 2087 42891
rect 12541 42857 12575 42891
rect 27537 42857 27571 42891
rect 13277 42721 13311 42755
rect 14105 42721 14139 42755
rect 19533 42721 19567 42755
rect 21925 42721 21959 42755
rect 24593 42721 24627 42755
rect 1593 42653 1627 42687
rect 2237 42653 2271 42687
rect 9505 42653 9539 42687
rect 10149 42653 10183 42687
rect 10425 42653 10459 42687
rect 12357 42653 12391 42687
rect 14381 42653 14415 42687
rect 15669 42653 15703 42687
rect 15761 42653 15795 42687
rect 15853 42653 15887 42687
rect 16037 42653 16071 42687
rect 19349 42653 19383 42687
rect 20269 42653 20303 42687
rect 22477 42653 22511 42687
rect 24685 42653 24719 42687
rect 25053 42653 25087 42687
rect 26801 42653 26835 42687
rect 28733 42653 28767 42687
rect 29009 42653 29043 42687
rect 29745 42653 29779 42687
rect 30021 42653 30055 42687
rect 11805 42585 11839 42619
rect 13093 42585 13127 42619
rect 16957 42585 16991 42619
rect 24409 42585 24443 42619
rect 25881 42585 25915 42619
rect 26617 42585 26651 42619
rect 27445 42585 27479 42619
rect 9689 42517 9723 42551
rect 15393 42517 15427 42551
rect 18245 42517 18279 42551
rect 22661 42517 22695 42551
rect 24777 42517 24811 42551
rect 24961 42517 24995 42551
rect 25973 42517 26007 42551
rect 28549 42517 28583 42551
rect 28917 42517 28951 42551
rect 29561 42517 29595 42551
rect 29929 42517 29963 42551
rect 1409 42313 1443 42347
rect 9689 42313 9723 42347
rect 12173 42313 12207 42347
rect 14565 42313 14599 42347
rect 15393 42313 15427 42347
rect 16129 42313 16163 42347
rect 20085 42313 20119 42347
rect 23489 42313 23523 42347
rect 27195 42313 27229 42347
rect 8585 42245 8619 42279
rect 8769 42245 8803 42279
rect 13553 42245 13587 42279
rect 14381 42245 14415 42279
rect 16773 42245 16807 42279
rect 22354 42245 22388 42279
rect 26985 42245 27019 42279
rect 1593 42177 1627 42211
rect 8401 42177 8435 42211
rect 9945 42177 9979 42211
rect 10038 42177 10072 42211
rect 10149 42177 10183 42211
rect 10333 42177 10367 42211
rect 11989 42177 12023 42211
rect 13369 42177 13403 42211
rect 15301 42177 15335 42211
rect 15945 42177 15979 42211
rect 17684 42177 17718 42211
rect 19257 42177 19291 42211
rect 19349 42177 19383 42211
rect 19901 42177 19935 42211
rect 20545 42177 20579 42211
rect 24869 42177 24903 42211
rect 26065 42177 26099 42211
rect 28181 42177 28215 42211
rect 28457 42177 28491 42211
rect 29745 42177 29779 42211
rect 29837 42177 29871 42211
rect 29929 42177 29963 42211
rect 30113 42177 30147 42211
rect 14657 42109 14691 42143
rect 17417 42109 17451 42143
rect 22109 42109 22143 42143
rect 16957 42041 16991 42075
rect 18797 42041 18831 42075
rect 20729 42041 20763 42075
rect 26249 42041 26283 42075
rect 14105 41973 14139 42007
rect 24961 41973 24995 42007
rect 27169 41973 27203 42007
rect 27353 41973 27387 42007
rect 29469 41973 29503 42007
rect 9321 41769 9355 41803
rect 13001 41769 13035 41803
rect 17693 41769 17727 41803
rect 19441 41769 19475 41803
rect 21833 41769 21867 41803
rect 26801 41769 26835 41803
rect 14289 41701 14323 41735
rect 16129 41701 16163 41735
rect 18521 41701 18555 41735
rect 24685 41701 24719 41735
rect 26433 41701 26467 41735
rect 26985 41701 27019 41735
rect 27445 41701 27479 41735
rect 10425 41633 10459 41667
rect 14749 41633 14783 41667
rect 19993 41633 20027 41667
rect 22293 41633 22327 41667
rect 23673 41633 23707 41667
rect 25421 41633 25455 41667
rect 25513 41633 25547 41667
rect 25605 41633 25639 41667
rect 25697 41633 25731 41667
rect 1593 41565 1627 41599
rect 8953 41565 8987 41599
rect 10701 41565 10735 41599
rect 14105 41565 14139 41599
rect 15016 41565 15050 41599
rect 16865 41565 16899 41599
rect 18337 41565 18371 41599
rect 20637 41565 20671 41599
rect 22937 41565 22971 41599
rect 23581 41565 23615 41599
rect 24501 41565 24535 41599
rect 27629 41565 27663 41599
rect 27905 41565 27939 41599
rect 28641 41565 28675 41599
rect 28733 41559 28767 41593
rect 28825 41562 28859 41596
rect 29021 41565 29055 41599
rect 29745 41565 29779 41599
rect 29929 41565 29963 41599
rect 30021 41565 30055 41599
rect 9137 41497 9171 41531
rect 11713 41497 11747 41531
rect 17601 41497 17635 41531
rect 19717 41497 19751 41531
rect 22385 41497 22419 41531
rect 26801 41497 26835 41531
rect 27813 41497 27847 41531
rect 1409 41429 1443 41463
rect 16957 41429 16991 41463
rect 19901 41429 19935 41463
rect 20821 41429 20855 41463
rect 22293 41429 22327 41463
rect 23029 41429 23063 41463
rect 25237 41429 25271 41463
rect 28365 41429 28399 41463
rect 29561 41429 29595 41463
rect 15393 41225 15427 41259
rect 18613 41225 18647 41259
rect 19257 41225 19291 41259
rect 20361 41225 20395 41259
rect 21189 41225 21223 41259
rect 25789 41225 25823 41259
rect 27721 41225 27755 41259
rect 15945 41157 15979 41191
rect 19165 41157 19199 41191
rect 20177 41157 20211 41191
rect 21097 41157 21131 41191
rect 25237 41157 25271 41191
rect 1593 41089 1627 41123
rect 15209 41089 15243 41123
rect 16681 41089 16715 41123
rect 17601 41089 17635 41123
rect 17690 41092 17724 41126
rect 17806 41089 17840 41123
rect 17969 41089 18003 41123
rect 18429 41089 18463 41123
rect 22477 41089 22511 41123
rect 23121 41089 23155 41123
rect 23305 41089 23339 41123
rect 25137 41089 25171 41123
rect 25973 41089 26007 41123
rect 27537 41089 27571 41123
rect 27813 41089 27847 41123
rect 28503 41089 28537 41123
rect 28622 41095 28656 41129
rect 28722 41089 28756 41123
rect 28929 41089 28963 41123
rect 29699 41089 29733 41123
rect 29834 41092 29868 41126
rect 29934 41089 29968 41123
rect 30113 41089 30147 41123
rect 16129 41021 16163 41055
rect 20453 41021 20487 41055
rect 26249 41021 26283 41055
rect 27353 41021 27387 41055
rect 19901 40953 19935 40987
rect 26157 40953 26191 40987
rect 1409 40885 1443 40919
rect 16865 40885 16899 40919
rect 17325 40885 17359 40919
rect 22569 40885 22603 40919
rect 23121 40885 23155 40919
rect 28273 40885 28307 40919
rect 29469 40885 29503 40919
rect 17233 40681 17267 40715
rect 17877 40681 17911 40715
rect 19349 40681 19383 40715
rect 21373 40613 21407 40647
rect 25329 40613 25363 40647
rect 22937 40545 22971 40579
rect 28273 40545 28307 40579
rect 30113 40545 30147 40579
rect 8033 40477 8067 40511
rect 8217 40477 8251 40511
rect 9853 40477 9887 40511
rect 9946 40477 9980 40511
rect 10057 40477 10091 40511
rect 10241 40477 10275 40511
rect 15761 40477 15795 40511
rect 16405 40477 16439 40511
rect 17049 40477 17083 40511
rect 17693 40477 17727 40511
rect 19257 40477 19291 40511
rect 20085 40477 20119 40511
rect 23121 40477 23155 40511
rect 23581 40477 23615 40511
rect 23857 40477 23891 40511
rect 25145 40477 25179 40511
rect 27169 40477 27203 40511
rect 27261 40477 27295 40511
rect 27353 40477 27387 40511
rect 27549 40477 27583 40511
rect 27997 40477 28031 40511
rect 29929 40477 29963 40511
rect 8401 40409 8435 40443
rect 18521 40409 18555 40443
rect 25881 40409 25915 40443
rect 26065 40409 26099 40443
rect 26249 40409 26283 40443
rect 26893 40409 26927 40443
rect 9597 40341 9631 40375
rect 15945 40341 15979 40375
rect 16589 40341 16623 40375
rect 18613 40341 18647 40375
rect 1409 40137 1443 40171
rect 8677 40137 8711 40171
rect 19993 40137 20027 40171
rect 21103 40137 21137 40171
rect 22753 40137 22787 40171
rect 23213 40137 23247 40171
rect 27261 40137 27295 40171
rect 27629 40137 27663 40171
rect 8493 40069 8527 40103
rect 11989 40069 12023 40103
rect 15945 40069 15979 40103
rect 17049 40069 17083 40103
rect 19809 40069 19843 40103
rect 20085 40069 20119 40103
rect 21005 40069 21039 40103
rect 24133 40069 24167 40103
rect 1593 40001 1627 40035
rect 8309 40001 8343 40035
rect 9853 40001 9887 40035
rect 9946 40001 9980 40035
rect 10057 40001 10091 40035
rect 10241 40001 10275 40035
rect 21189 40001 21223 40035
rect 21281 40001 21315 40035
rect 22109 40001 22143 40035
rect 23397 40001 23431 40035
rect 24317 40001 24351 40035
rect 26157 40001 26191 40035
rect 27445 40001 27479 40035
rect 27721 40001 27755 40035
rect 28457 40001 28491 40035
rect 29837 40001 29871 40035
rect 23673 39933 23707 39967
rect 24501 39933 24535 39967
rect 28181 39933 28215 39967
rect 18337 39865 18371 39899
rect 26341 39865 26375 39899
rect 9597 39797 9631 39831
rect 12081 39797 12115 39831
rect 16037 39797 16071 39831
rect 19533 39797 19567 39831
rect 23581 39797 23615 39831
rect 30021 39797 30055 39831
rect 13001 39593 13035 39627
rect 14289 39593 14323 39627
rect 16221 39593 16255 39627
rect 18705 39593 18739 39627
rect 23397 39593 23431 39627
rect 26985 39593 27019 39627
rect 10609 39457 10643 39491
rect 16589 39457 16623 39491
rect 20913 39457 20947 39491
rect 24777 39457 24811 39491
rect 24869 39457 24903 39491
rect 1593 39389 1627 39423
rect 10333 39389 10367 39423
rect 11621 39389 11655 39423
rect 17325 39389 17359 39423
rect 17592 39389 17626 39423
rect 21180 39389 21214 39423
rect 23305 39389 23339 39423
rect 24593 39389 24627 39423
rect 24685 39389 24719 39423
rect 26801 39389 26835 39423
rect 27997 39389 28031 39423
rect 28733 39389 28767 39423
rect 29837 39389 29871 39423
rect 11866 39321 11900 39355
rect 14197 39321 14231 39355
rect 15117 39321 15151 39355
rect 15301 39321 15335 39355
rect 16773 39321 16807 39355
rect 19717 39321 19751 39355
rect 23121 39321 23155 39355
rect 1409 39253 1443 39287
rect 16681 39253 16715 39287
rect 19809 39253 19843 39287
rect 22293 39253 22327 39287
rect 24409 39253 24443 39287
rect 28181 39253 28215 39287
rect 28917 39253 28951 39287
rect 30021 39253 30055 39287
rect 11529 39049 11563 39083
rect 12817 39049 12851 39083
rect 17233 39049 17267 39083
rect 18797 39049 18831 39083
rect 24869 39049 24903 39083
rect 24961 39049 24995 39083
rect 27169 39049 27203 39083
rect 8401 38981 8435 39015
rect 8585 38981 8619 39015
rect 14350 38981 14384 39015
rect 17049 38981 17083 39015
rect 19533 38981 19567 39015
rect 20821 38981 20855 39015
rect 20913 38981 20947 39015
rect 1593 38913 1627 38947
rect 11785 38913 11819 38947
rect 11894 38913 11928 38947
rect 12010 38913 12044 38947
rect 12173 38913 12207 38947
rect 13093 38913 13127 38947
rect 13182 38913 13216 38947
rect 13277 38913 13311 38947
rect 13473 38913 13507 38947
rect 17969 38913 18003 38947
rect 18613 38913 18647 38947
rect 19349 38913 19383 38947
rect 22293 38913 22327 38947
rect 24777 38913 24811 38947
rect 25145 38913 25179 38947
rect 26985 38913 27019 38947
rect 28365 38913 28399 38947
rect 29101 38913 29135 38947
rect 29837 38913 29871 38947
rect 14105 38845 14139 38879
rect 17325 38845 17359 38879
rect 20821 38845 20855 38879
rect 23029 38845 23063 38879
rect 23305 38845 23339 38879
rect 1409 38777 1443 38811
rect 16773 38777 16807 38811
rect 24593 38777 24627 38811
rect 8769 38709 8803 38743
rect 15485 38709 15519 38743
rect 18061 38709 18095 38743
rect 20361 38709 20395 38743
rect 22477 38709 22511 38743
rect 28549 38709 28583 38743
rect 29285 38709 29319 38743
rect 30021 38709 30055 38743
rect 11069 38505 11103 38539
rect 17233 38505 17267 38539
rect 18061 38505 18095 38539
rect 20453 38505 20487 38539
rect 21097 38505 21131 38539
rect 11805 38369 11839 38403
rect 23490 38369 23524 38403
rect 23765 38369 23799 38403
rect 24685 38369 24719 38403
rect 25973 38369 26007 38403
rect 1593 38301 1627 38335
rect 9689 38301 9723 38335
rect 9956 38301 9990 38335
rect 12081 38301 12115 38335
rect 14105 38301 14139 38335
rect 17969 38301 18003 38335
rect 19257 38301 19291 38335
rect 20361 38301 20395 38335
rect 21005 38301 21039 38335
rect 23581 38301 23615 38335
rect 23673 38301 23707 38335
rect 24409 38301 24443 38335
rect 25697 38301 25731 38335
rect 27353 38301 27387 38335
rect 29837 38301 29871 38335
rect 14372 38233 14406 38267
rect 17141 38233 17175 38267
rect 28181 38233 28215 38267
rect 1409 38165 1443 38199
rect 15485 38165 15519 38199
rect 19441 38165 19475 38199
rect 23305 38165 23339 38199
rect 27537 38165 27571 38199
rect 28273 38165 28307 38199
rect 30021 38165 30055 38199
rect 8125 37961 8159 37995
rect 9229 37961 9263 37995
rect 10977 37961 11011 37995
rect 13001 37961 13035 37995
rect 15301 37961 15335 37995
rect 16681 37961 16715 37995
rect 18705 37961 18739 37995
rect 23673 37961 23707 37995
rect 26065 37961 26099 37995
rect 27261 37961 27295 37995
rect 29929 37961 29963 37995
rect 9045 37893 9079 37927
rect 9873 37893 9907 37927
rect 14013 37893 14047 37927
rect 18613 37893 18647 37927
rect 24685 37893 24719 37927
rect 24887 37893 24921 37927
rect 25881 37893 25915 37927
rect 1593 37825 1627 37859
rect 8309 37825 8343 37859
rect 8861 37825 8895 37859
rect 9689 37825 9723 37859
rect 10793 37825 10827 37859
rect 11888 37825 11922 37859
rect 16957 37825 16991 37859
rect 17049 37825 17083 37859
rect 17141 37825 17175 37859
rect 17325 37825 17359 37859
rect 17785 37825 17819 37859
rect 19993 37825 20027 37859
rect 23673 37825 23707 37859
rect 24797 37825 24831 37859
rect 25053 37825 25087 37859
rect 27445 37825 27479 37859
rect 27629 37825 27663 37859
rect 27721 37825 27755 37859
rect 28273 37825 28307 37859
rect 29745 37825 29779 37859
rect 30021 37825 30055 37859
rect 11621 37757 11655 37791
rect 26157 37757 26191 37791
rect 28549 37757 28583 37791
rect 24501 37689 24535 37723
rect 1409 37621 1443 37655
rect 10057 37621 10091 37655
rect 17969 37621 18003 37655
rect 20177 37621 20211 37655
rect 25605 37621 25639 37655
rect 29561 37621 29595 37655
rect 4353 37417 4387 37451
rect 9597 37417 9631 37451
rect 12449 37417 12483 37451
rect 17233 37417 17267 37451
rect 21281 37417 21315 37451
rect 26525 37417 26559 37451
rect 28365 37417 28399 37451
rect 18245 37281 18279 37315
rect 18705 37281 18739 37315
rect 24593 37281 24627 37315
rect 24685 37281 24719 37315
rect 24869 37281 24903 37315
rect 8953 37213 8987 37247
rect 11621 37213 11655 37247
rect 11713 37213 11747 37247
rect 11805 37213 11839 37247
rect 11989 37213 12023 37247
rect 12725 37213 12759 37247
rect 12817 37213 12851 37247
rect 12909 37213 12943 37247
rect 13093 37213 13127 37247
rect 15117 37213 15151 37247
rect 17141 37213 17175 37247
rect 18429 37213 18463 37247
rect 18613 37213 18647 37247
rect 19257 37213 19291 37247
rect 19513 37213 19547 37247
rect 21281 37213 21315 37247
rect 21925 37213 21959 37247
rect 22385 37213 22419 37247
rect 24777 37213 24811 37247
rect 26709 37213 26743 37247
rect 26985 37213 27019 37247
rect 27629 37213 27663 37247
rect 27813 37213 27847 37247
rect 27905 37213 27939 37247
rect 28641 37213 28675 37247
rect 28733 37213 28767 37247
rect 28825 37213 28859 37247
rect 29009 37213 29043 37247
rect 29745 37213 29779 37247
rect 30021 37213 30055 37247
rect 4261 37145 4295 37179
rect 15362 37145 15396 37179
rect 29561 37145 29595 37179
rect 11345 37077 11379 37111
rect 16497 37077 16531 37111
rect 20637 37077 20671 37111
rect 22569 37077 22603 37111
rect 24409 37077 24443 37111
rect 26893 37077 26927 37111
rect 27445 37077 27479 37111
rect 29929 37077 29963 37111
rect 1409 36873 1443 36907
rect 9321 36873 9355 36907
rect 15025 36873 15059 36907
rect 26341 36873 26375 36907
rect 8309 36805 8343 36839
rect 9137 36805 9171 36839
rect 27813 36805 27847 36839
rect 1593 36737 1627 36771
rect 8125 36737 8159 36771
rect 8953 36737 8987 36771
rect 13461 36737 13495 36771
rect 13737 36737 13771 36771
rect 15301 36737 15335 36771
rect 15393 36737 15427 36771
rect 15485 36740 15519 36774
rect 15669 36737 15703 36771
rect 17877 36737 17911 36771
rect 18981 36737 19015 36771
rect 21833 36737 21867 36771
rect 22109 36737 22143 36771
rect 26065 36737 26099 36771
rect 27629 36737 27663 36771
rect 27905 36737 27939 36771
rect 28641 36737 28675 36771
rect 28733 36737 28767 36771
rect 28825 36737 28859 36771
rect 29009 36737 29043 36771
rect 29699 36737 29733 36771
rect 29837 36737 29871 36771
rect 29929 36737 29963 36771
rect 30113 36737 30147 36771
rect 22293 36669 22327 36703
rect 22477 36669 22511 36703
rect 25697 36669 25731 36703
rect 25973 36669 26007 36703
rect 26157 36669 26191 36703
rect 8493 36601 8527 36635
rect 18061 36601 18095 36635
rect 27445 36601 27479 36635
rect 20269 36533 20303 36567
rect 28365 36533 28399 36567
rect 29469 36533 29503 36567
rect 8217 36329 8251 36363
rect 11069 36329 11103 36363
rect 15209 36329 15243 36363
rect 18245 36329 18279 36363
rect 19441 36329 19475 36363
rect 25145 36329 25179 36363
rect 1409 36261 1443 36295
rect 20821 36261 20855 36295
rect 25697 36261 25731 36295
rect 19993 36193 20027 36227
rect 21465 36193 21499 36227
rect 26249 36193 26283 36227
rect 28089 36193 28123 36227
rect 1593 36125 1627 36159
rect 8401 36125 8435 36159
rect 9689 36125 9723 36159
rect 9945 36125 9979 36159
rect 15025 36125 15059 36159
rect 16957 36125 16991 36159
rect 19257 36125 19291 36159
rect 20177 36125 20211 36159
rect 21189 36125 21223 36159
rect 22017 36125 22051 36159
rect 22845 36125 22879 36159
rect 24961 36125 24995 36159
rect 25973 36125 26007 36159
rect 27353 36125 27387 36159
rect 27629 36125 27663 36159
rect 28365 36125 28399 36159
rect 29745 36125 29779 36159
rect 29929 36125 29963 36159
rect 30021 36125 30055 36159
rect 22201 36057 22235 36091
rect 22385 36057 22419 36091
rect 25881 36057 25915 36091
rect 27537 36057 27571 36091
rect 20361 35989 20395 36023
rect 21281 35989 21315 36023
rect 23029 35989 23063 36023
rect 26065 35989 26099 36023
rect 27169 35989 27203 36023
rect 29561 35989 29595 36023
rect 21189 35785 21223 35819
rect 23765 35785 23799 35819
rect 27721 35785 27755 35819
rect 8861 35717 8895 35751
rect 9045 35717 9079 35751
rect 25329 35717 25363 35751
rect 1593 35649 1627 35683
rect 19257 35649 19291 35683
rect 20177 35649 20211 35683
rect 21005 35649 21039 35683
rect 22385 35649 22419 35683
rect 22641 35649 22675 35683
rect 24777 35649 24811 35683
rect 25053 35649 25087 35683
rect 26985 35649 27019 35683
rect 27997 35649 28031 35683
rect 28089 35649 28123 35683
rect 28181 35649 28215 35683
rect 28365 35649 28399 35683
rect 20821 35581 20855 35615
rect 24317 35581 24351 35615
rect 28825 35581 28859 35615
rect 29101 35581 29135 35615
rect 19441 35513 19475 35547
rect 1409 35445 1443 35479
rect 9229 35445 9263 35479
rect 19993 35445 20027 35479
rect 27169 35445 27203 35479
rect 10885 35241 10919 35275
rect 11713 35241 11747 35275
rect 12357 35241 12391 35275
rect 13461 35241 13495 35275
rect 18061 35241 18095 35275
rect 20821 35241 20855 35275
rect 23765 35241 23799 35275
rect 24593 35241 24627 35275
rect 16589 35173 16623 35207
rect 26985 35173 27019 35207
rect 17049 35105 17083 35139
rect 18521 35105 18555 35139
rect 1593 35037 1627 35071
rect 10701 35037 10735 35071
rect 11529 35037 11563 35071
rect 12173 35037 12207 35071
rect 13277 35037 13311 35071
rect 14565 35037 14599 35071
rect 14749 35037 14783 35071
rect 15853 35037 15887 35071
rect 18613 35037 18647 35071
rect 19441 35037 19475 35071
rect 21833 35037 21867 35071
rect 22109 35037 22143 35071
rect 23673 35037 23707 35071
rect 23857 35037 23891 35071
rect 24409 35037 24443 35071
rect 27077 35037 27111 35071
rect 27629 35037 27663 35071
rect 28181 35037 28215 35071
rect 29837 35037 29871 35071
rect 17141 34969 17175 35003
rect 19708 34969 19742 35003
rect 28365 34969 28399 35003
rect 1409 34901 1443 34935
rect 16037 34901 16071 34935
rect 17049 34901 17083 34935
rect 18521 34901 18555 34935
rect 21925 34901 21959 34935
rect 30021 34901 30055 34935
rect 1409 34697 1443 34731
rect 9873 34697 9907 34731
rect 14289 34697 14323 34731
rect 17325 34697 17359 34731
rect 19073 34697 19107 34731
rect 20453 34697 20487 34731
rect 28181 34697 28215 34731
rect 28917 34697 28951 34731
rect 10425 34629 10459 34663
rect 15945 34629 15979 34663
rect 18153 34629 18187 34663
rect 18981 34629 19015 34663
rect 27353 34629 27387 34663
rect 1593 34561 1627 34595
rect 9689 34561 9723 34595
rect 11621 34561 11655 34595
rect 12357 34561 12391 34595
rect 13093 34561 13127 34595
rect 14105 34561 14139 34595
rect 14749 34561 14783 34595
rect 19625 34561 19659 34595
rect 20269 34561 20303 34595
rect 27169 34561 27203 34595
rect 27997 34561 28031 34595
rect 28733 34561 28767 34595
rect 29745 34561 29779 34595
rect 29837 34561 29871 34595
rect 29929 34561 29963 34595
rect 30113 34561 30147 34595
rect 13277 34493 13311 34527
rect 16129 34493 16163 34527
rect 17325 34493 17359 34527
rect 17417 34493 17451 34527
rect 18337 34493 18371 34527
rect 10609 34425 10643 34459
rect 11805 34357 11839 34391
rect 12449 34357 12483 34391
rect 14933 34357 14967 34391
rect 16865 34357 16899 34391
rect 19809 34357 19843 34391
rect 27445 34357 27479 34391
rect 29469 34357 29503 34391
rect 10517 34153 10551 34187
rect 16589 34153 16623 34187
rect 20085 34153 20119 34187
rect 28181 34153 28215 34187
rect 17601 34085 17635 34119
rect 25145 34085 25179 34119
rect 26341 34085 26375 34119
rect 11069 34017 11103 34051
rect 12725 34017 12759 34051
rect 17969 34017 18003 34051
rect 1593 33949 1627 33983
rect 10793 33949 10827 33983
rect 13369 33949 13403 33983
rect 15301 33949 15335 33983
rect 19993 33949 20027 33983
rect 24593 33949 24627 33983
rect 24777 33949 24811 33983
rect 24961 33949 24995 33983
rect 25789 33949 25823 33983
rect 26157 33949 26191 33983
rect 27997 33949 28031 33983
rect 28733 33949 28767 33983
rect 29837 33949 29871 33983
rect 12817 33881 12851 33915
rect 14197 33881 14231 33915
rect 18061 33881 18095 33915
rect 18153 33881 18187 33915
rect 19349 33881 19383 33915
rect 24869 33881 24903 33915
rect 25973 33881 26007 33915
rect 26065 33881 26099 33915
rect 1409 33813 1443 33847
rect 10977 33813 11011 33847
rect 12247 33813 12281 33847
rect 12725 33813 12759 33847
rect 13553 33813 13587 33847
rect 14289 33813 14323 33847
rect 19441 33813 19475 33847
rect 28917 33813 28951 33847
rect 30021 33813 30055 33847
rect 11805 33609 11839 33643
rect 15485 33609 15519 33643
rect 17601 33609 17635 33643
rect 26249 33609 26283 33643
rect 9781 33541 9815 33575
rect 10793 33541 10827 33575
rect 13093 33541 13127 33575
rect 14289 33541 14323 33575
rect 16773 33541 16807 33575
rect 18245 33541 18279 33575
rect 19901 33541 19935 33575
rect 24961 33541 24995 33575
rect 25881 33541 25915 33575
rect 25973 33541 26007 33575
rect 1593 33473 1627 33507
rect 9597 33473 9631 33507
rect 10885 33473 10919 33507
rect 11621 33473 11655 33507
rect 13185 33473 13219 33507
rect 14105 33473 14139 33507
rect 15301 33473 15335 33507
rect 17509 33473 17543 33507
rect 20453 33473 20487 33507
rect 24685 33473 24719 33507
rect 24869 33473 24903 33507
rect 25053 33473 25087 33507
rect 25697 33473 25731 33507
rect 26065 33473 26099 33507
rect 29101 33473 29135 33507
rect 29837 33473 29871 33507
rect 10793 33405 10827 33439
rect 13093 33405 13127 33439
rect 14381 33405 14415 33439
rect 15577 33405 15611 33439
rect 16957 33405 16991 33439
rect 10333 33337 10367 33371
rect 12633 33337 12667 33371
rect 13829 33337 13863 33371
rect 15025 33337 15059 33371
rect 1409 33269 1443 33303
rect 20637 33269 20671 33303
rect 25237 33269 25271 33303
rect 29285 33269 29319 33303
rect 30021 33269 30055 33303
rect 10701 33065 10735 33099
rect 16221 33065 16255 33099
rect 18337 33065 18371 33099
rect 19349 33065 19383 33099
rect 15577 32997 15611 33031
rect 16865 32997 16899 33031
rect 25697 32997 25731 33031
rect 11161 32929 11195 32963
rect 17417 32929 17451 32963
rect 19717 32929 19751 32963
rect 1593 32861 1627 32895
rect 9781 32861 9815 32895
rect 11253 32861 11287 32895
rect 13553 32861 13587 32895
rect 14197 32861 14231 32895
rect 17141 32861 17175 32895
rect 18153 32861 18187 32895
rect 20545 32861 20579 32895
rect 20637 32861 20671 32895
rect 21281 32861 21315 32895
rect 21465 32861 21499 32895
rect 21833 32861 21867 32895
rect 22477 32861 22511 32895
rect 22661 32861 22695 32895
rect 22753 32861 22787 32895
rect 25145 32861 25179 32895
rect 25513 32861 25547 32895
rect 28733 32861 28767 32895
rect 29837 32861 29871 32895
rect 9597 32793 9631 32827
rect 9965 32793 9999 32827
rect 11805 32793 11839 32827
rect 14464 32793 14498 32827
rect 16129 32793 16163 32827
rect 19809 32793 19843 32827
rect 19901 32793 19935 32827
rect 25329 32793 25363 32827
rect 25421 32793 25455 32827
rect 1409 32725 1443 32759
rect 11161 32725 11195 32759
rect 17325 32725 17359 32759
rect 20821 32725 20855 32759
rect 21741 32725 21775 32759
rect 22293 32725 22327 32759
rect 28917 32725 28951 32759
rect 30021 32725 30055 32759
rect 9965 32521 9999 32555
rect 13185 32521 13219 32555
rect 14105 32521 14139 32555
rect 17233 32521 17267 32555
rect 18981 32521 19015 32555
rect 21833 32521 21867 32555
rect 9781 32453 9815 32487
rect 11897 32453 11931 32487
rect 15301 32453 15335 32487
rect 17049 32453 17083 32487
rect 17325 32453 17359 32487
rect 22201 32453 22235 32487
rect 22339 32453 22373 32487
rect 28181 32453 28215 32487
rect 29101 32453 29135 32487
rect 1593 32385 1627 32419
rect 9597 32385 9631 32419
rect 14381 32385 14415 32419
rect 14470 32385 14504 32419
rect 14570 32385 14604 32419
rect 14749 32385 14783 32419
rect 15945 32385 15979 32419
rect 18797 32385 18831 32419
rect 19625 32385 19659 32419
rect 19892 32385 19926 32419
rect 22017 32385 22051 32419
rect 22109 32385 22143 32419
rect 23397 32385 23431 32419
rect 23765 32385 23799 32419
rect 25605 32385 25639 32419
rect 27997 32385 28031 32419
rect 28257 32385 28291 32419
rect 28733 32385 28767 32419
rect 29377 32385 29411 32419
rect 29469 32385 29503 32419
rect 29561 32385 29595 32419
rect 29745 32385 29779 32419
rect 19073 32317 19107 32351
rect 22477 32317 22511 32351
rect 25881 32317 25915 32351
rect 21005 32249 21039 32283
rect 1409 32181 1443 32215
rect 15393 32181 15427 32215
rect 16129 32181 16163 32215
rect 16773 32181 16807 32215
rect 18521 32181 18555 32215
rect 27813 32181 27847 32215
rect 2789 31977 2823 32011
rect 11621 31977 11655 32011
rect 13369 31977 13403 32011
rect 14289 31977 14323 32011
rect 16313 31977 16347 32011
rect 20085 31977 20119 32011
rect 21465 31977 21499 32011
rect 24409 31977 24443 32011
rect 26893 31977 26927 32011
rect 28089 31977 28123 32011
rect 30113 31977 30147 32011
rect 9505 31909 9539 31943
rect 10425 31909 10459 31943
rect 17877 31909 17911 31943
rect 10885 31841 10919 31875
rect 11989 31841 12023 31875
rect 18337 31841 18371 31875
rect 22477 31841 22511 31875
rect 27261 31841 27295 31875
rect 28549 31841 28583 31875
rect 1869 31773 1903 31807
rect 2421 31773 2455 31807
rect 2605 31773 2639 31807
rect 9689 31773 9723 31807
rect 10977 31773 11011 31807
rect 12173 31773 12207 31807
rect 13277 31773 13311 31807
rect 14105 31773 14139 31807
rect 16221 31773 16255 31807
rect 18429 31773 18463 31807
rect 20269 31773 20303 31807
rect 21649 31773 21683 31807
rect 21741 31773 21775 31807
rect 21925 31773 21959 31807
rect 22017 31773 22051 31807
rect 24593 31773 24627 31807
rect 24777 31773 24811 31807
rect 24869 31773 24903 31807
rect 26157 31773 26191 31807
rect 26341 31773 26375 31807
rect 27445 31773 27479 31807
rect 29745 31773 29779 31807
rect 18337 31705 18371 31739
rect 22744 31705 22778 31739
rect 27353 31705 27387 31739
rect 28641 31705 28675 31739
rect 29929 31705 29963 31739
rect 1685 31637 1719 31671
rect 10885 31637 10919 31671
rect 12081 31637 12115 31671
rect 23857 31637 23891 31671
rect 28549 31637 28583 31671
rect 12449 31433 12483 31467
rect 13277 31433 13311 31467
rect 14059 31433 14093 31467
rect 17233 31433 17267 31467
rect 22661 31433 22695 31467
rect 23121 31433 23155 31467
rect 24041 31433 24075 31467
rect 24961 31433 24995 31467
rect 26433 31433 26467 31467
rect 27629 31433 27663 31467
rect 2421 31365 2455 31399
rect 9873 31365 9907 31399
rect 10701 31365 10735 31399
rect 12357 31365 12391 31399
rect 19349 31365 19383 31399
rect 28733 31365 28767 31399
rect 29653 31365 29687 31399
rect 1869 31297 1903 31331
rect 2605 31297 2639 31331
rect 9689 31297 9723 31331
rect 10517 31297 10551 31331
rect 13185 31297 13219 31331
rect 15761 31297 15795 31331
rect 15853 31297 15887 31331
rect 15945 31297 15979 31331
rect 16129 31297 16163 31331
rect 17325 31297 17359 31331
rect 22293 31297 22327 31331
rect 22477 31297 22511 31331
rect 23305 31297 23339 31331
rect 23581 31297 23615 31331
rect 24225 31297 24259 31331
rect 25145 31297 25179 31331
rect 25881 31297 25915 31331
rect 26065 31297 26099 31331
rect 26157 31297 26191 31331
rect 26249 31297 26283 31331
rect 28273 31297 28307 31331
rect 28457 31297 28491 31331
rect 13829 31229 13863 31263
rect 17233 31229 17267 31263
rect 18245 31229 18279 31263
rect 24501 31229 24535 31263
rect 25421 31229 25455 31263
rect 27537 31229 27571 31263
rect 27721 31229 27755 31263
rect 29561 31229 29595 31263
rect 29745 31229 29779 31263
rect 2789 31161 2823 31195
rect 10057 31161 10091 31195
rect 15485 31161 15519 31195
rect 19533 31161 19567 31195
rect 29193 31161 29227 31195
rect 1685 31093 1719 31127
rect 10885 31093 10919 31127
rect 16773 31093 16807 31127
rect 18797 31093 18831 31127
rect 23489 31093 23523 31127
rect 24409 31093 24443 31127
rect 25329 31093 25363 31127
rect 27169 31093 27203 31127
rect 26065 30889 26099 30923
rect 28365 30889 28399 30923
rect 30113 30889 30147 30923
rect 20177 30821 20211 30855
rect 24409 30821 24443 30855
rect 24777 30753 24811 30787
rect 26433 30753 26467 30787
rect 28089 30753 28123 30787
rect 1409 30685 1443 30719
rect 2329 30685 2363 30719
rect 9689 30685 9723 30719
rect 9873 30685 9907 30719
rect 11069 30685 11103 30719
rect 15439 30685 15473 30719
rect 15577 30685 15611 30719
rect 15669 30685 15703 30719
rect 15853 30685 15887 30719
rect 18705 30685 18739 30719
rect 19349 30685 19383 30719
rect 19993 30685 20027 30719
rect 24593 30685 24627 30719
rect 24869 30685 24903 30719
rect 26249 30685 26283 30719
rect 26525 30685 26559 30719
rect 28641 30685 28675 30719
rect 28730 30685 28764 30719
rect 28846 30685 28880 30719
rect 29009 30685 29043 30719
rect 29929 30685 29963 30719
rect 10057 30617 10091 30651
rect 16313 30617 16347 30651
rect 29745 30617 29779 30651
rect 1593 30549 1627 30583
rect 2145 30549 2179 30583
rect 11253 30549 11287 30583
rect 15209 30549 15243 30583
rect 17601 30549 17635 30583
rect 18521 30549 18555 30583
rect 19533 30549 19567 30583
rect 12909 30345 12943 30379
rect 11774 30277 11808 30311
rect 19441 30277 19475 30311
rect 19657 30277 19691 30311
rect 28641 30277 28675 30311
rect 29561 30277 29595 30311
rect 29653 30277 29687 30311
rect 1409 30209 1443 30243
rect 2329 30209 2363 30243
rect 11529 30209 11563 30243
rect 13829 30209 13863 30243
rect 13921 30209 13955 30243
rect 14013 30209 14047 30243
rect 14197 30209 14231 30243
rect 17601 30209 17635 30243
rect 17868 30209 17902 30243
rect 27537 30209 27571 30243
rect 28089 30209 28123 30243
rect 25605 30141 25639 30175
rect 25881 30141 25915 30175
rect 29561 30141 29595 30175
rect 1593 30005 1627 30039
rect 2145 30005 2179 30039
rect 13553 30005 13587 30039
rect 18981 30005 19015 30039
rect 19625 30005 19659 30039
rect 19809 30005 19843 30039
rect 27721 30005 27755 30039
rect 28273 30005 28307 30039
rect 29101 30005 29135 30039
rect 17049 29801 17083 29835
rect 18705 29801 18739 29835
rect 19901 29801 19935 29835
rect 25789 29801 25823 29835
rect 30021 29801 30055 29835
rect 27077 29733 27111 29767
rect 26157 29665 26191 29699
rect 1409 29597 1443 29631
rect 2329 29597 2363 29631
rect 12725 29597 12759 29631
rect 13001 29597 13035 29631
rect 14361 29597 14395 29631
rect 14473 29597 14507 29631
rect 14565 29594 14599 29628
rect 14749 29597 14783 29631
rect 15761 29597 15795 29631
rect 18061 29597 18095 29631
rect 19257 29597 19291 29631
rect 21097 29597 21131 29631
rect 21189 29597 21223 29631
rect 21281 29597 21315 29631
rect 21465 29597 21499 29631
rect 25973 29597 26007 29631
rect 26249 29597 26283 29631
rect 26893 29597 26927 29631
rect 27832 29597 27866 29631
rect 28089 29575 28123 29609
rect 28733 29597 28767 29631
rect 29837 29597 29871 29631
rect 27997 29529 28031 29563
rect 1593 29461 1627 29495
rect 2145 29461 2179 29495
rect 14105 29461 14139 29495
rect 20821 29461 20855 29495
rect 27629 29461 27663 29495
rect 28917 29461 28951 29495
rect 15209 29257 15243 29291
rect 18061 29257 18095 29291
rect 21833 29257 21867 29291
rect 22845 29257 22879 29291
rect 28365 29257 28399 29291
rect 30021 29257 30055 29291
rect 13921 29189 13955 29223
rect 16948 29189 16982 29223
rect 19800 29189 19834 29223
rect 1409 29121 1443 29155
rect 12771 29121 12805 29155
rect 12909 29121 12943 29155
rect 13001 29121 13035 29155
rect 13185 29121 13219 29155
rect 19533 29121 19567 29155
rect 22017 29121 22051 29155
rect 22293 29121 22327 29155
rect 23029 29121 23063 29155
rect 23121 29121 23155 29155
rect 23305 29121 23339 29155
rect 23397 29121 23431 29155
rect 27675 29121 27709 29155
rect 27813 29121 27847 29155
rect 27905 29121 27939 29155
rect 28621 29121 28655 29155
rect 28733 29121 28767 29155
rect 28825 29121 28859 29155
rect 29009 29121 29043 29155
rect 29837 29121 29871 29155
rect 16681 29053 16715 29087
rect 27445 29053 27479 29087
rect 1593 28985 1627 29019
rect 12541 28985 12575 29019
rect 22109 28985 22143 29019
rect 22201 28985 22235 29019
rect 20913 28917 20947 28951
rect 15577 28713 15611 28747
rect 25145 28713 25179 28747
rect 18613 28577 18647 28611
rect 19349 28577 19383 28611
rect 19533 28577 19567 28611
rect 22661 28577 22695 28611
rect 28457 28577 28491 28611
rect 1409 28509 1443 28543
rect 14361 28509 14395 28543
rect 14454 28509 14488 28543
rect 14570 28509 14604 28543
rect 14749 28509 14783 28543
rect 15393 28509 15427 28543
rect 16129 28509 16163 28543
rect 16865 28509 16899 28543
rect 18521 28509 18555 28543
rect 18705 28509 18739 28543
rect 19257 28509 19291 28543
rect 21005 28509 21039 28543
rect 21189 28509 21223 28543
rect 21741 28509 21775 28543
rect 22017 28509 22051 28543
rect 22937 28509 22971 28543
rect 24593 28509 24627 28543
rect 24961 28509 24995 28543
rect 27445 28509 27479 28543
rect 27721 28509 27755 28543
rect 28181 28509 28215 28543
rect 29837 28509 29871 28543
rect 16313 28441 16347 28475
rect 20085 28441 20119 28475
rect 24777 28441 24811 28475
rect 24869 28441 24903 28475
rect 1593 28373 1627 28407
rect 14105 28373 14139 28407
rect 16957 28373 16991 28407
rect 19533 28373 19567 28407
rect 20177 28373 20211 28407
rect 21005 28373 21039 28407
rect 27261 28373 27295 28407
rect 27629 28373 27663 28407
rect 30021 28373 30055 28407
rect 14473 28169 14507 28203
rect 24041 28169 24075 28203
rect 25053 28169 25087 28203
rect 29377 28169 29411 28203
rect 13185 28101 13219 28135
rect 15945 28101 15979 28135
rect 24685 28101 24719 28135
rect 24777 28101 24811 28135
rect 16037 28033 16071 28067
rect 18429 28033 18463 28067
rect 18696 28033 18730 28067
rect 21925 28033 21959 28067
rect 22661 28033 22695 28067
rect 22928 28033 22962 28067
rect 24501 28033 24535 28067
rect 24869 28033 24903 28067
rect 27537 28033 27571 28067
rect 28549 28033 28583 28067
rect 28641 28033 28675 28067
rect 28733 28033 28767 28067
rect 28917 28033 28951 28067
rect 29653 28033 29687 28067
rect 29745 28033 29779 28067
rect 29837 28033 29871 28067
rect 30021 28033 30055 28067
rect 15853 27965 15887 27999
rect 28273 27965 28307 27999
rect 15485 27897 15519 27931
rect 27721 27897 27755 27931
rect 19809 27829 19843 27863
rect 22109 27829 22143 27863
rect 16405 27625 16439 27659
rect 21557 27625 21591 27659
rect 14565 27557 14599 27591
rect 17049 27557 17083 27591
rect 25329 27557 25363 27591
rect 30113 27557 30147 27591
rect 15025 27489 15059 27523
rect 21557 27489 21591 27523
rect 27721 27489 27755 27523
rect 27813 27489 27847 27523
rect 1409 27421 1443 27455
rect 12081 27421 12115 27455
rect 12348 27421 12382 27455
rect 14381 27421 14415 27455
rect 21649 27421 21683 27455
rect 24777 27421 24811 27455
rect 25145 27421 25179 27455
rect 25789 27421 25823 27455
rect 26065 27421 26099 27455
rect 27445 27421 27479 27455
rect 27629 27421 27663 27455
rect 28008 27421 28042 27455
rect 28733 27421 28767 27455
rect 29929 27421 29963 27455
rect 15292 27353 15326 27387
rect 17325 27353 17359 27387
rect 17601 27353 17635 27387
rect 21373 27353 21407 27387
rect 24961 27353 24995 27387
rect 25053 27353 25087 27387
rect 29745 27353 29779 27387
rect 1593 27285 1627 27319
rect 13461 27285 13495 27319
rect 17509 27285 17543 27319
rect 21833 27285 21867 27319
rect 28181 27285 28215 27319
rect 28917 27285 28951 27319
rect 2145 27081 2179 27115
rect 12541 27081 12575 27115
rect 15669 27081 15703 27115
rect 23213 27081 23247 27115
rect 24961 27081 24995 27115
rect 25421 27081 25455 27115
rect 26249 27081 26283 27115
rect 27537 27081 27571 27115
rect 27997 27081 28031 27115
rect 28733 27081 28767 27115
rect 29929 27081 29963 27115
rect 13553 27013 13587 27047
rect 15485 27013 15519 27047
rect 18889 27013 18923 27047
rect 24593 27013 24627 27047
rect 24685 27013 24719 27047
rect 26065 27013 26099 27047
rect 28549 27013 28583 27047
rect 1409 26945 1443 26979
rect 2329 26945 2363 26979
rect 12357 26945 12391 26979
rect 14473 26945 14507 26979
rect 15191 26945 15225 26979
rect 22293 26945 22327 26979
rect 23397 26945 23431 26979
rect 23673 26945 23707 26979
rect 24409 26945 24443 26979
rect 24777 26945 24811 26979
rect 26341 26945 26375 26979
rect 27629 26945 27663 26979
rect 28365 26945 28399 26979
rect 29101 26945 29135 26979
rect 15761 26877 15795 26911
rect 27445 26877 27479 26911
rect 29837 26877 29871 26911
rect 30021 26877 30055 26911
rect 22477 26809 22511 26843
rect 25789 26809 25823 26843
rect 27077 26809 27111 26843
rect 1593 26741 1627 26775
rect 13645 26741 13679 26775
rect 14657 26741 14691 26775
rect 20177 26741 20211 26775
rect 23581 26741 23615 26775
rect 29469 26741 29503 26775
rect 17049 26537 17083 26571
rect 30113 26537 30147 26571
rect 2145 26469 2179 26503
rect 25881 26469 25915 26503
rect 28089 26469 28123 26503
rect 28917 26469 28951 26503
rect 15669 26401 15703 26435
rect 1409 26333 1443 26367
rect 2329 26333 2363 26367
rect 13185 26333 13219 26367
rect 15925 26333 15959 26367
rect 25329 26333 25363 26367
rect 25697 26333 25731 26367
rect 28273 26333 28307 26367
rect 28733 26333 28767 26367
rect 29745 26333 29779 26367
rect 25513 26265 25547 26299
rect 25605 26265 25639 26299
rect 29929 26265 29963 26299
rect 1593 26197 1627 26231
rect 13277 26197 13311 26231
rect 13001 25993 13035 26027
rect 28181 25993 28215 26027
rect 28641 25993 28675 26027
rect 29101 25993 29135 26027
rect 29929 25993 29963 26027
rect 18613 25925 18647 25959
rect 30021 25925 30055 25959
rect 1409 25857 1443 25891
rect 2329 25857 2363 25891
rect 13093 25857 13127 25891
rect 17877 25857 17911 25891
rect 19349 25857 19383 25891
rect 22477 25857 22511 25891
rect 22569 25857 22603 25891
rect 22753 25857 22787 25891
rect 22845 25857 22879 25891
rect 27813 25857 27847 25891
rect 27997 25857 28031 25891
rect 28457 25857 28491 25891
rect 13001 25789 13035 25823
rect 18797 25789 18831 25823
rect 29929 25789 29963 25823
rect 2145 25721 2179 25755
rect 12541 25721 12575 25755
rect 29469 25721 29503 25755
rect 1593 25653 1627 25687
rect 17969 25653 18003 25687
rect 19533 25653 19567 25687
rect 22293 25653 22327 25687
rect 1685 25449 1719 25483
rect 24501 25449 24535 25483
rect 27445 25449 27479 25483
rect 28365 25449 28399 25483
rect 30021 25449 30055 25483
rect 17417 25381 17451 25415
rect 21005 25381 21039 25415
rect 28825 25381 28859 25415
rect 17969 25313 18003 25347
rect 19625 25313 19659 25347
rect 24961 25313 24995 25347
rect 1869 25245 1903 25279
rect 16405 25245 16439 25279
rect 18521 25245 18555 25279
rect 22385 25245 22419 25279
rect 22477 25245 22511 25279
rect 22661 25245 22695 25279
rect 22753 25245 22787 25279
rect 24685 25245 24719 25279
rect 24869 25245 24903 25279
rect 25513 25245 25547 25279
rect 26525 25245 26559 25279
rect 28181 25245 28215 25279
rect 29009 25245 29043 25279
rect 29837 25245 29871 25279
rect 17693 25177 17727 25211
rect 17877 25177 17911 25211
rect 19892 25177 19926 25211
rect 25697 25177 25731 25211
rect 27353 25177 27387 25211
rect 27997 25177 28031 25211
rect 16589 25109 16623 25143
rect 18613 25109 18647 25143
rect 22201 25109 22235 25143
rect 26709 25109 26743 25143
rect 13277 24905 13311 24939
rect 20637 24905 20671 24939
rect 26617 24905 26651 24939
rect 28273 24905 28307 24939
rect 29929 24905 29963 24939
rect 13093 24837 13127 24871
rect 28089 24837 28123 24871
rect 1409 24769 1443 24803
rect 2329 24769 2363 24803
rect 14177 24769 14211 24803
rect 17141 24769 17175 24803
rect 17233 24772 17267 24806
rect 17346 24769 17380 24803
rect 17509 24769 17543 24803
rect 17969 24769 18003 24803
rect 18236 24769 18270 24803
rect 20913 24769 20947 24803
rect 21005 24769 21039 24803
rect 21097 24769 21131 24803
rect 21281 24769 21315 24803
rect 23121 24769 23155 24803
rect 23305 24769 23339 24803
rect 23673 24769 23707 24803
rect 24317 24769 24351 24803
rect 24501 24769 24535 24803
rect 24777 24769 24811 24803
rect 26801 24769 26835 24803
rect 27445 24769 27479 24803
rect 30021 24769 30055 24803
rect 13369 24701 13403 24735
rect 13921 24701 13955 24735
rect 21833 24701 21867 24735
rect 23397 24701 23431 24735
rect 23489 24701 23523 24735
rect 25329 24701 25363 24735
rect 28365 24701 28399 24735
rect 29929 24701 29963 24735
rect 1593 24633 1627 24667
rect 2145 24633 2179 24667
rect 15301 24633 15335 24667
rect 27813 24633 27847 24667
rect 12817 24565 12851 24599
rect 16865 24565 16899 24599
rect 19349 24565 19383 24599
rect 22063 24565 22097 24599
rect 23857 24565 23891 24599
rect 24685 24565 24719 24599
rect 25559 24565 25593 24599
rect 29469 24565 29503 24599
rect 14289 24361 14323 24395
rect 17877 24361 17911 24395
rect 19257 24361 19291 24395
rect 23305 24361 23339 24395
rect 24409 24361 24443 24395
rect 28181 24361 28215 24395
rect 28825 24361 28859 24395
rect 2145 24293 2179 24327
rect 12909 24293 12943 24327
rect 1409 24157 1443 24191
rect 2329 24157 2363 24191
rect 13185 24157 13219 24191
rect 13461 24157 13495 24191
rect 14105 24157 14139 24191
rect 16497 24157 16531 24191
rect 18521 24157 18555 24191
rect 18613 24157 18647 24191
rect 19441 24157 19475 24191
rect 19533 24157 19567 24191
rect 19717 24157 19751 24191
rect 19809 24157 19843 24191
rect 21097 24157 21131 24191
rect 21189 24157 21223 24191
rect 21281 24157 21315 24191
rect 21465 24157 21499 24191
rect 24665 24157 24699 24191
rect 24777 24157 24811 24191
rect 24869 24157 24903 24191
rect 25053 24157 25087 24191
rect 25605 24157 25639 24191
rect 28365 24157 28399 24191
rect 29009 24157 29043 24191
rect 13369 24089 13403 24123
rect 16764 24089 16798 24123
rect 22017 24089 22051 24123
rect 29929 24089 29963 24123
rect 1593 24021 1627 24055
rect 20821 24021 20855 24055
rect 25697 24021 25731 24055
rect 30021 24021 30055 24055
rect 17417 23817 17451 23851
rect 17785 23817 17819 23851
rect 21189 23817 21223 23851
rect 22753 23817 22787 23851
rect 23397 23817 23431 23851
rect 24409 23817 24443 23851
rect 25421 23817 25455 23851
rect 27813 23749 27847 23783
rect 29929 23749 29963 23783
rect 1409 23681 1443 23715
rect 2329 23681 2363 23715
rect 13185 23681 13219 23715
rect 17601 23681 17635 23715
rect 17877 23681 17911 23715
rect 19533 23681 19567 23715
rect 21097 23681 21131 23715
rect 21281 23681 21315 23715
rect 22017 23681 22051 23715
rect 22201 23681 22235 23715
rect 22569 23681 22603 23715
rect 23581 23681 23615 23715
rect 24593 23681 24627 23715
rect 25329 23681 25363 23715
rect 28641 23681 28675 23715
rect 29193 23681 29227 23715
rect 22293 23613 22327 23647
rect 22385 23613 22419 23647
rect 23857 23613 23891 23647
rect 24869 23613 24903 23647
rect 30113 23613 30147 23647
rect 2145 23545 2179 23579
rect 27997 23545 28031 23579
rect 28457 23545 28491 23579
rect 1593 23477 1627 23511
rect 13369 23477 13403 23511
rect 19717 23477 19751 23511
rect 23765 23477 23799 23511
rect 24777 23477 24811 23511
rect 29285 23477 29319 23511
rect 23305 23273 23339 23307
rect 24409 23273 24443 23307
rect 28917 23273 28951 23307
rect 29929 23273 29963 23307
rect 2145 23205 2179 23239
rect 15485 23205 15519 23239
rect 26433 23205 26467 23239
rect 28089 23205 28123 23239
rect 14105 23137 14139 23171
rect 19809 23137 19843 23171
rect 21925 23137 21959 23171
rect 24869 23137 24903 23171
rect 1409 23069 1443 23103
rect 2329 23069 2363 23103
rect 14361 23069 14395 23103
rect 21649 23069 21683 23103
rect 22937 23069 22971 23103
rect 23121 23069 23155 23103
rect 24593 23069 24627 23103
rect 24777 23069 24811 23103
rect 26709 23069 26743 23103
rect 28273 23069 28307 23103
rect 28733 23069 28767 23103
rect 29745 23069 29779 23103
rect 20076 23001 20110 23035
rect 26985 23001 27019 23035
rect 29561 23001 29595 23035
rect 1593 22933 1627 22967
rect 21189 22933 21223 22967
rect 26893 22933 26927 22967
rect 17969 22729 18003 22763
rect 21005 22729 21039 22763
rect 21833 22729 21867 22763
rect 28255 22729 28289 22763
rect 29837 22729 29871 22763
rect 27353 22661 27387 22695
rect 27537 22661 27571 22695
rect 27629 22661 27663 22695
rect 28733 22661 28767 22695
rect 29653 22661 29687 22695
rect 1409 22593 1443 22627
rect 2329 22593 2363 22627
rect 17877 22593 17911 22627
rect 21005 22593 21039 22627
rect 21281 22593 21315 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 22293 22593 22327 22627
rect 23397 22593 23431 22627
rect 23581 22593 23615 22627
rect 25421 22593 25455 22627
rect 25697 22593 25731 22627
rect 28549 22593 28583 22627
rect 29469 22593 29503 22627
rect 23673 22525 23707 22559
rect 28825 22525 28859 22559
rect 2145 22457 2179 22491
rect 21097 22457 21131 22491
rect 23213 22457 23247 22491
rect 27077 22457 27111 22491
rect 1593 22389 1627 22423
rect 25237 22389 25271 22423
rect 25605 22389 25639 22423
rect 26433 22185 26467 22219
rect 30021 22185 30055 22219
rect 27169 22049 27203 22083
rect 27353 22049 27387 22083
rect 28733 22049 28767 22083
rect 1869 21981 1903 22015
rect 19257 21981 19291 22015
rect 22477 21981 22511 22015
rect 25053 21981 25087 22015
rect 25320 21981 25354 22015
rect 28163 21981 28197 22015
rect 29837 21981 29871 22015
rect 27261 21913 27295 21947
rect 27813 21913 27847 21947
rect 28457 21913 28491 21947
rect 29653 21913 29687 21947
rect 1685 21845 1719 21879
rect 19901 21845 19935 21879
rect 22569 21845 22603 21879
rect 26783 21845 26817 21879
rect 28641 21845 28675 21879
rect 18705 21641 18739 21675
rect 24041 21641 24075 21675
rect 25237 21641 25271 21675
rect 27629 21641 27663 21675
rect 29101 21641 29135 21675
rect 30113 21641 30147 21675
rect 27537 21573 27571 21607
rect 29745 21573 29779 21607
rect 29929 21573 29963 21607
rect 1409 21505 1443 21539
rect 2329 21505 2363 21539
rect 16681 21505 16715 21539
rect 17877 21505 17911 21539
rect 18521 21505 18555 21539
rect 18797 21505 18831 21539
rect 19257 21505 19291 21539
rect 19441 21505 19475 21539
rect 24225 21505 24259 21539
rect 24501 21505 24535 21539
rect 24685 21505 24719 21539
rect 25421 21505 25455 21539
rect 25697 21505 25731 21539
rect 25881 21505 25915 21539
rect 28181 21505 28215 21539
rect 29285 21505 29319 21539
rect 28457 21437 28491 21471
rect 1593 21369 1627 21403
rect 2145 21301 2179 21335
rect 16865 21301 16899 21335
rect 18061 21301 18095 21335
rect 18521 21301 18555 21335
rect 19257 21301 19291 21335
rect 16957 21097 16991 21131
rect 24409 21097 24443 21131
rect 27445 21097 27479 21131
rect 28089 21097 28123 21131
rect 30113 21097 30147 21131
rect 17877 20961 17911 20995
rect 19257 20961 19291 20995
rect 29009 20961 29043 20995
rect 1409 20893 1443 20927
rect 16773 20893 16807 20927
rect 17601 20893 17635 20927
rect 17693 20893 17727 20927
rect 19513 20893 19547 20927
rect 24593 20893 24627 20927
rect 24869 20893 24903 20927
rect 25053 20893 25087 20927
rect 27629 20893 27663 20927
rect 28273 20893 28307 20927
rect 29929 20893 29963 20927
rect 28825 20825 28859 20859
rect 29745 20825 29779 20859
rect 1593 20757 1627 20791
rect 20637 20757 20671 20791
rect 29451 20553 29485 20587
rect 29929 20553 29963 20587
rect 20085 20485 20119 20519
rect 28273 20485 28307 20519
rect 1409 20417 1443 20451
rect 16129 20417 16163 20451
rect 16681 20417 16715 20451
rect 16937 20417 16971 20451
rect 18613 20417 18647 20451
rect 29745 20417 29779 20451
rect 20269 20349 20303 20383
rect 30021 20349 30055 20383
rect 15945 20281 15979 20315
rect 18061 20281 18095 20315
rect 1593 20213 1627 20247
rect 18705 20213 18739 20247
rect 28365 20213 28399 20247
rect 2145 20009 2179 20043
rect 16865 20009 16899 20043
rect 23305 20009 23339 20043
rect 28641 20009 28675 20043
rect 30021 20009 30055 20043
rect 17601 19941 17635 19975
rect 1409 19805 1443 19839
rect 2329 19805 2363 19839
rect 16497 19805 16531 19839
rect 16681 19805 16715 19839
rect 17785 19805 17819 19839
rect 18245 19805 18279 19839
rect 20177 19805 20211 19839
rect 20361 19805 20395 19839
rect 21925 19805 21959 19839
rect 24593 19805 24627 19839
rect 24869 19805 24903 19839
rect 25053 19805 25087 19839
rect 28457 19805 28491 19839
rect 29837 19805 29871 19839
rect 20545 19737 20579 19771
rect 22192 19737 22226 19771
rect 28273 19737 28307 19771
rect 1593 19669 1627 19703
rect 24409 19669 24443 19703
rect 2145 19465 2179 19499
rect 17325 19465 17359 19499
rect 22937 19465 22971 19499
rect 27611 19465 27645 19499
rect 28089 19465 28123 19499
rect 28733 19465 28767 19499
rect 29929 19465 29963 19499
rect 17693 19397 17727 19431
rect 27905 19397 27939 19431
rect 28181 19397 28215 19431
rect 30021 19397 30055 19431
rect 1409 19329 1443 19363
rect 2329 19329 2363 19363
rect 17785 19329 17819 19363
rect 18521 19329 18555 19363
rect 18797 19329 18831 19363
rect 19165 19329 19199 19363
rect 19901 19329 19935 19363
rect 20085 19329 20119 19363
rect 20269 19329 20303 19363
rect 23121 19329 23155 19363
rect 25697 19329 25731 19363
rect 25881 19329 25915 19363
rect 26157 19329 26191 19363
rect 26341 19329 26375 19363
rect 28917 19329 28951 19363
rect 29745 19329 29779 19363
rect 17877 19261 17911 19295
rect 18981 19261 19015 19295
rect 23397 19261 23431 19295
rect 23305 19193 23339 19227
rect 29469 19193 29503 19227
rect 1593 19125 1627 19159
rect 2329 18921 2363 18955
rect 28365 18921 28399 18955
rect 29929 18921 29963 18955
rect 26985 18853 27019 18887
rect 25605 18785 25639 18819
rect 28917 18785 28951 18819
rect 1869 18717 1903 18751
rect 2513 18717 2547 18751
rect 24593 18717 24627 18751
rect 24869 18717 24903 18751
rect 25053 18717 25087 18751
rect 28641 18717 28675 18751
rect 29745 18717 29779 18751
rect 25850 18649 25884 18683
rect 29561 18649 29595 18683
rect 1685 18581 1719 18615
rect 24409 18581 24443 18615
rect 28825 18581 28859 18615
rect 23213 18377 23247 18411
rect 28641 18377 28675 18411
rect 29745 18377 29779 18411
rect 28457 18309 28491 18343
rect 29561 18309 29595 18343
rect 1409 18241 1443 18275
rect 2329 18241 2363 18275
rect 21833 18241 21867 18275
rect 22100 18241 22134 18275
rect 23857 18241 23891 18275
rect 24041 18241 24075 18275
rect 24777 18241 24811 18275
rect 25513 18241 25547 18275
rect 28273 18241 28307 18275
rect 29837 18241 29871 18275
rect 24133 18173 24167 18207
rect 25237 18173 25271 18207
rect 1593 18105 1627 18139
rect 29285 18105 29319 18139
rect 2145 18037 2179 18071
rect 23673 18037 23707 18071
rect 24593 18037 24627 18071
rect 23857 17833 23891 17867
rect 24961 17833 24995 17867
rect 25697 17833 25731 17867
rect 28825 17833 28859 17867
rect 28181 17765 28215 17799
rect 21097 17697 21131 17731
rect 26157 17697 26191 17731
rect 1409 17629 1443 17663
rect 19625 17629 19659 17663
rect 19901 17629 19935 17663
rect 20729 17629 20763 17663
rect 22477 17629 22511 17663
rect 22744 17629 22778 17663
rect 25881 17629 25915 17663
rect 26065 17629 26099 17663
rect 28365 17629 28399 17663
rect 29009 17629 29043 17663
rect 29929 17629 29963 17663
rect 19809 17561 19843 17595
rect 20913 17561 20947 17595
rect 24869 17561 24903 17595
rect 1593 17493 1627 17527
rect 19441 17493 19475 17527
rect 30021 17493 30055 17527
rect 22477 17289 22511 17323
rect 27537 17289 27571 17323
rect 29193 17289 29227 17323
rect 28273 17221 28307 17255
rect 29929 17221 29963 17255
rect 1409 17153 1443 17187
rect 2329 17153 2363 17187
rect 17877 17153 17911 17187
rect 18429 17153 18463 17187
rect 18613 17153 18647 17187
rect 18981 17153 19015 17187
rect 19625 17153 19659 17187
rect 19717 17153 19751 17187
rect 19901 17153 19935 17187
rect 19993 17153 20027 17187
rect 22661 17153 22695 17187
rect 23857 17153 23891 17187
rect 24041 17153 24075 17187
rect 24317 17153 24351 17187
rect 24501 17153 24535 17187
rect 27353 17153 27387 17187
rect 29377 17153 29411 17187
rect 18889 17085 18923 17119
rect 22937 17085 22971 17119
rect 27629 17085 27663 17119
rect 28457 17085 28491 17119
rect 2145 17017 2179 17051
rect 27077 17017 27111 17051
rect 1593 16949 1627 16983
rect 17693 16949 17727 16983
rect 19441 16949 19475 16983
rect 22845 16949 22879 16983
rect 30021 16949 30055 16983
rect 17233 16745 17267 16779
rect 18107 16745 18141 16779
rect 19257 16745 19291 16779
rect 20361 16745 20395 16779
rect 27629 16745 27663 16779
rect 16865 16609 16899 16643
rect 19901 16609 19935 16643
rect 20729 16609 20763 16643
rect 27077 16609 27111 16643
rect 1409 16541 1443 16575
rect 2329 16541 2363 16575
rect 16221 16541 16255 16575
rect 17049 16541 17083 16575
rect 17877 16541 17911 16575
rect 19442 16541 19476 16575
rect 19743 16541 19777 16575
rect 20545 16541 20579 16575
rect 20637 16541 20671 16575
rect 20821 16541 20855 16575
rect 28071 16541 28105 16575
rect 28365 16541 28399 16575
rect 30113 16541 30147 16575
rect 19533 16473 19567 16507
rect 19625 16473 19659 16507
rect 27261 16473 27295 16507
rect 28641 16473 28675 16507
rect 1593 16405 1627 16439
rect 2145 16405 2179 16439
rect 16405 16405 16439 16439
rect 26691 16405 26725 16439
rect 27169 16405 27203 16439
rect 28549 16405 28583 16439
rect 29929 16405 29963 16439
rect 28163 16201 28197 16235
rect 17132 16133 17166 16167
rect 25329 16133 25363 16167
rect 27721 16133 27755 16167
rect 28641 16133 28675 16167
rect 28733 16133 28767 16167
rect 1869 16065 1903 16099
rect 2513 16065 2547 16099
rect 16865 16065 16899 16099
rect 18705 16065 18739 16099
rect 20545 16065 20579 16099
rect 21833 16065 21867 16099
rect 25053 16065 25087 16099
rect 25237 16065 25271 16099
rect 25421 16065 25455 16099
rect 28457 16065 28491 16099
rect 29929 16065 29963 16099
rect 20269 15997 20303 16031
rect 30113 15997 30147 16031
rect 18245 15929 18279 15963
rect 22017 15929 22051 15963
rect 25605 15929 25639 15963
rect 1685 15861 1719 15895
rect 2329 15861 2363 15895
rect 19349 15861 19383 15895
rect 27169 15657 27203 15691
rect 28825 15657 28859 15691
rect 16865 15589 16899 15623
rect 18705 15589 18739 15623
rect 20637 15589 20671 15623
rect 25789 15589 25823 15623
rect 17325 15521 17359 15555
rect 21281 15521 21315 15555
rect 27721 15521 27755 15555
rect 1409 15453 1443 15487
rect 2329 15453 2363 15487
rect 16681 15453 16715 15487
rect 19349 15453 19383 15487
rect 19717 15453 19751 15487
rect 20177 15453 20211 15487
rect 20453 15453 20487 15487
rect 21557 15453 21591 15487
rect 25237 15453 25271 15487
rect 25605 15453 25639 15487
rect 27445 15453 27479 15487
rect 29009 15453 29043 15487
rect 17592 15385 17626 15419
rect 25421 15385 25455 15419
rect 25513 15385 25547 15419
rect 27629 15385 27663 15419
rect 29929 15385 29963 15419
rect 1593 15317 1627 15351
rect 2145 15317 2179 15351
rect 30021 15317 30055 15351
rect 23213 15113 23247 15147
rect 23765 15113 23799 15147
rect 24685 15113 24719 15147
rect 26249 15113 26283 15147
rect 28273 15113 28307 15147
rect 1409 14977 1443 15011
rect 19349 14977 19383 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 21097 14977 21131 15011
rect 21189 14977 21223 15011
rect 22100 14977 22134 15011
rect 23949 14977 23983 15011
rect 24869 14977 24903 15011
rect 26433 14977 26467 15011
rect 27169 14977 27203 15011
rect 28181 14977 28215 15011
rect 29561 14977 29595 15011
rect 19625 14909 19659 14943
rect 21833 14909 21867 14943
rect 24225 14909 24259 14943
rect 25145 14909 25179 14943
rect 28365 14909 28399 14943
rect 29285 14909 29319 14943
rect 27353 14841 27387 14875
rect 1593 14773 1627 14807
rect 20637 14773 20671 14807
rect 24133 14773 24167 14807
rect 25053 14773 25087 14807
rect 27813 14773 27847 14807
rect 19257 14569 19291 14603
rect 20361 14569 20395 14603
rect 20821 14569 20855 14603
rect 22477 14569 22511 14603
rect 26341 14569 26375 14603
rect 27077 14501 27111 14535
rect 28365 14501 28399 14535
rect 30021 14501 30055 14535
rect 20453 14433 20487 14467
rect 22937 14433 22971 14467
rect 27629 14433 27663 14467
rect 28825 14433 28859 14467
rect 1409 14365 1443 14399
rect 19487 14365 19521 14399
rect 19625 14365 19659 14399
rect 19717 14365 19751 14399
rect 19901 14365 19935 14399
rect 20637 14365 20671 14399
rect 22661 14365 22695 14399
rect 22845 14365 22879 14399
rect 25789 14365 25823 14399
rect 26157 14365 26191 14399
rect 27445 14365 27479 14399
rect 29837 14365 29871 14399
rect 20361 14297 20395 14331
rect 25973 14297 26007 14331
rect 26065 14297 26099 14331
rect 28917 14297 28951 14331
rect 1593 14229 1627 14263
rect 27537 14229 27571 14263
rect 28825 14229 28859 14263
rect 27537 14025 27571 14059
rect 21833 13957 21867 13991
rect 27445 13957 27479 13991
rect 28457 13957 28491 13991
rect 28641 13957 28675 13991
rect 1409 13889 1443 13923
rect 22017 13889 22051 13923
rect 23949 13889 23983 13923
rect 24225 13889 24259 13923
rect 24409 13889 24443 13923
rect 25605 13889 25639 13923
rect 29561 13889 29595 13923
rect 25881 13821 25915 13855
rect 28733 13821 28767 13855
rect 29285 13821 29319 13855
rect 1593 13685 1627 13719
rect 22201 13685 22235 13719
rect 23765 13685 23799 13719
rect 28181 13685 28215 13719
rect 23213 13481 23247 13515
rect 24409 13481 24443 13515
rect 28365 13413 28399 13447
rect 27537 13345 27571 13379
rect 27721 13345 27755 13379
rect 28917 13345 28951 13379
rect 30113 13345 30147 13379
rect 1409 13277 1443 13311
rect 20729 13277 20763 13311
rect 20822 13277 20856 13311
rect 21005 13277 21039 13311
rect 21235 13277 21269 13311
rect 21833 13277 21867 13311
rect 24593 13277 24627 13311
rect 24869 13277 24903 13311
rect 25053 13277 25087 13311
rect 26065 13277 26099 13311
rect 26433 13277 26467 13311
rect 27445 13277 27479 13311
rect 28641 13277 28675 13311
rect 21097 13209 21131 13243
rect 22100 13209 22134 13243
rect 26249 13209 26283 13243
rect 26341 13209 26375 13243
rect 29929 13209 29963 13243
rect 1593 13141 1627 13175
rect 21373 13141 21407 13175
rect 26617 13141 26651 13175
rect 27077 13141 27111 13175
rect 28825 13141 28859 13175
rect 20637 12937 20671 12971
rect 22753 12937 22787 12971
rect 24685 12937 24719 12971
rect 28641 12937 28675 12971
rect 27629 12869 27663 12903
rect 28457 12869 28491 12903
rect 28733 12869 28767 12903
rect 20545 12801 20579 12835
rect 20729 12801 20763 12835
rect 22937 12801 22971 12835
rect 24869 12801 24903 12835
rect 25605 12801 25639 12835
rect 27445 12801 27479 12835
rect 23121 12733 23155 12767
rect 23213 12733 23247 12767
rect 25145 12733 25179 12767
rect 29285 12733 29319 12767
rect 29561 12733 29595 12767
rect 28181 12665 28215 12699
rect 25053 12597 25087 12631
rect 25835 12597 25869 12631
rect 2053 12393 2087 12427
rect 25789 12393 25823 12427
rect 26985 12393 27019 12427
rect 30113 12325 30147 12359
rect 27537 12257 27571 12291
rect 1409 12189 1443 12223
rect 17325 12189 17359 12223
rect 17969 12189 18003 12223
rect 20729 12189 20763 12223
rect 20821 12189 20855 12223
rect 21005 12189 21039 12223
rect 21097 12189 21131 12223
rect 25237 12189 25271 12223
rect 25605 12189 25639 12223
rect 28181 12189 28215 12223
rect 25421 12121 25455 12155
rect 25513 12121 25547 12155
rect 26709 12121 26743 12155
rect 27445 12121 27479 12155
rect 29929 12121 29963 12155
rect 1593 12053 1627 12087
rect 17509 12053 17543 12087
rect 18153 12053 18187 12087
rect 20545 12053 20579 12087
rect 27353 12053 27387 12087
rect 28411 12053 28445 12087
rect 19257 11849 19291 11883
rect 24685 11849 24719 11883
rect 25697 11849 25731 11883
rect 28641 11849 28675 11883
rect 27721 11781 27755 11815
rect 28365 11781 28399 11815
rect 1409 11713 1443 11747
rect 17877 11713 17911 11747
rect 18144 11713 18178 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 24869 11713 24903 11747
rect 25881 11713 25915 11747
rect 27629 11713 27663 11747
rect 28825 11713 28859 11747
rect 25053 11645 25087 11679
rect 25145 11645 25179 11679
rect 26157 11645 26191 11679
rect 27813 11645 27847 11679
rect 29285 11645 29319 11679
rect 29561 11645 29595 11679
rect 26065 11577 26099 11611
rect 1593 11509 1627 11543
rect 19717 11509 19751 11543
rect 27261 11509 27295 11543
rect 19257 11305 19291 11339
rect 21281 11305 21315 11339
rect 26709 11305 26743 11339
rect 28181 11305 28215 11339
rect 28917 11305 28951 11339
rect 30021 11305 30055 11339
rect 20821 11169 20855 11203
rect 20913 11169 20947 11203
rect 25789 11169 25823 11203
rect 1409 11101 1443 11135
rect 2329 11101 2363 11135
rect 19487 11101 19521 11135
rect 19606 11101 19640 11135
rect 19717 11101 19751 11135
rect 19913 11101 19947 11135
rect 20545 11101 20579 11135
rect 20729 11101 20763 11135
rect 21097 11101 21131 11135
rect 24593 11101 24627 11135
rect 24869 11101 24903 11135
rect 25053 11101 25087 11135
rect 25605 11101 25639 11135
rect 26617 11101 26651 11135
rect 28089 11101 28123 11135
rect 28733 11101 28767 11135
rect 29837 11101 29871 11135
rect 1593 10965 1627 10999
rect 2145 10965 2179 10999
rect 24409 10965 24443 10999
rect 19257 10761 19291 10795
rect 23213 10761 23247 10795
rect 27077 10761 27111 10795
rect 27537 10761 27571 10795
rect 28089 10761 28123 10795
rect 29377 10761 29411 10795
rect 18144 10693 18178 10727
rect 26249 10693 26283 10727
rect 28365 10693 28399 10727
rect 1409 10625 1443 10659
rect 17877 10625 17911 10659
rect 20085 10625 20119 10659
rect 21097 10625 21131 10659
rect 21281 10625 21315 10659
rect 22100 10625 22134 10659
rect 24041 10625 24075 10659
rect 24317 10625 24351 10659
rect 24501 10625 24535 10659
rect 26433 10625 26467 10659
rect 27445 10625 27479 10659
rect 19809 10557 19843 10591
rect 21833 10557 21867 10591
rect 27629 10557 27663 10591
rect 1593 10421 1627 10455
rect 21097 10421 21131 10455
rect 23857 10421 23891 10455
rect 21925 10217 21959 10251
rect 22753 10217 22787 10251
rect 23121 10217 23155 10251
rect 26341 10217 26375 10251
rect 28089 10149 28123 10183
rect 20177 10081 20211 10115
rect 21465 10081 21499 10115
rect 21557 10081 21591 10115
rect 1409 10013 1443 10047
rect 2329 10013 2363 10047
rect 19901 10013 19935 10047
rect 21189 10013 21223 10047
rect 21373 10013 21407 10047
rect 21741 10013 21775 10047
rect 22937 10013 22971 10047
rect 23213 10013 23247 10047
rect 27905 10013 27939 10047
rect 28733 10013 28767 10047
rect 26249 9945 26283 9979
rect 29745 9945 29779 9979
rect 1593 9877 1627 9911
rect 2145 9877 2179 9911
rect 28825 9877 28859 9911
rect 29837 9877 29871 9911
rect 21281 9673 21315 9707
rect 24133 9673 24167 9707
rect 29377 9673 29411 9707
rect 19993 9605 20027 9639
rect 20177 9537 20211 9571
rect 20453 9537 20487 9571
rect 20913 9537 20947 9571
rect 21097 9537 21131 9571
rect 22845 9537 22879 9571
rect 24317 9537 24351 9571
rect 27077 9537 27111 9571
rect 27169 9537 27203 9571
rect 20361 9469 20395 9503
rect 23121 9469 23155 9503
rect 28365 9469 28399 9503
rect 22661 9333 22695 9367
rect 23029 9333 23063 9367
rect 27077 9333 27111 9367
rect 20269 9129 20303 9163
rect 22937 9129 22971 9163
rect 30021 9129 30055 9163
rect 20177 9061 20211 9095
rect 27077 9061 27111 9095
rect 25421 8993 25455 9027
rect 27721 8993 27755 9027
rect 28825 8993 28859 9027
rect 1409 8925 1443 8959
rect 2329 8925 2363 8959
rect 20085 8925 20119 8959
rect 21557 8925 21591 8959
rect 21824 8925 21858 8959
rect 25145 8925 25179 8959
rect 28641 8925 28675 8959
rect 29837 8925 29871 8959
rect 20361 8857 20395 8891
rect 24501 8857 24535 8891
rect 27537 8857 27571 8891
rect 28733 8857 28767 8891
rect 1593 8789 1627 8823
rect 2145 8789 2179 8823
rect 24593 8789 24627 8823
rect 27445 8789 27479 8823
rect 28273 8789 28307 8823
rect 26341 8585 26375 8619
rect 27537 8585 27571 8619
rect 29101 8585 29135 8619
rect 25421 8517 25455 8551
rect 27353 8517 27387 8551
rect 1409 8449 1443 8483
rect 24225 8449 24259 8483
rect 24501 8449 24535 8483
rect 24685 8449 24719 8483
rect 25237 8449 25271 8483
rect 26157 8449 26191 8483
rect 25973 8381 26007 8415
rect 28089 8381 28123 8415
rect 1593 8313 1627 8347
rect 26985 8313 27019 8347
rect 24041 8245 24075 8279
rect 27353 8245 27387 8279
rect 23029 8041 23063 8075
rect 2145 7973 2179 8007
rect 25513 7905 25547 7939
rect 26801 7905 26835 7939
rect 1409 7837 1443 7871
rect 2329 7837 2363 7871
rect 22845 7837 22879 7871
rect 23121 7837 23155 7871
rect 25789 7837 25823 7871
rect 27077 7837 27111 7871
rect 28273 7837 28307 7871
rect 29929 7837 29963 7871
rect 30113 7769 30147 7803
rect 1593 7701 1627 7735
rect 22661 7701 22695 7735
rect 28365 7701 28399 7735
rect 29101 7497 29135 7531
rect 28089 7429 28123 7463
rect 1409 7361 1443 7395
rect 24317 7361 24351 7395
rect 24501 7361 24535 7395
rect 24593 7361 24627 7395
rect 26341 7361 26375 7395
rect 26985 7361 27019 7395
rect 26065 7293 26099 7327
rect 26157 7293 26191 7327
rect 26249 7293 26283 7327
rect 1593 7157 1627 7191
rect 24133 7157 24167 7191
rect 25881 7157 25915 7191
rect 27169 7157 27203 7191
rect 22937 6953 22971 6987
rect 30021 6953 30055 6987
rect 25421 6817 25455 6851
rect 25697 6817 25731 6851
rect 25789 6817 25823 6851
rect 28733 6817 28767 6851
rect 21557 6749 21591 6783
rect 25605 6749 25639 6783
rect 25881 6749 25915 6783
rect 26985 6749 27019 6783
rect 27629 6749 27663 6783
rect 29837 6749 29871 6783
rect 21824 6681 21858 6715
rect 28457 6681 28491 6715
rect 26801 6613 26835 6647
rect 27445 6613 27479 6647
rect 28089 6613 28123 6647
rect 28549 6613 28583 6647
rect 2053 6409 2087 6443
rect 24685 6409 24719 6443
rect 28549 6409 28583 6443
rect 29837 6409 29871 6443
rect 23572 6341 23606 6375
rect 27445 6341 27479 6375
rect 28641 6341 28675 6375
rect 1409 6273 1443 6307
rect 29745 6273 29779 6307
rect 23305 6205 23339 6239
rect 28825 6205 28859 6239
rect 29929 6205 29963 6239
rect 1593 6137 1627 6171
rect 27537 6069 27571 6103
rect 28181 6069 28215 6103
rect 29377 6069 29411 6103
rect 28089 5865 28123 5899
rect 28825 5865 28859 5899
rect 29929 5865 29963 5899
rect 25605 5729 25639 5763
rect 26893 5729 26927 5763
rect 1409 5661 1443 5695
rect 25513 5661 25547 5695
rect 25697 5661 25731 5695
rect 25789 5661 25823 5695
rect 26617 5661 26651 5695
rect 27997 5661 28031 5695
rect 29009 5661 29043 5695
rect 30113 5661 30147 5695
rect 1593 5525 1627 5559
rect 25329 5525 25363 5559
rect 23305 5321 23339 5355
rect 27997 5321 28031 5355
rect 29837 5321 29871 5355
rect 24409 5253 24443 5287
rect 27169 5253 27203 5287
rect 28733 5253 28767 5287
rect 1409 5185 1443 5219
rect 23213 5185 23247 5219
rect 24225 5185 24259 5219
rect 24501 5185 24535 5219
rect 25605 5185 25639 5219
rect 26985 5185 27019 5219
rect 27629 5185 27663 5219
rect 28181 5185 28215 5219
rect 29745 5185 29779 5219
rect 25329 5117 25363 5151
rect 25513 5117 25547 5151
rect 25697 5117 25731 5151
rect 25789 5117 25823 5151
rect 29929 5117 29963 5151
rect 1593 4981 1627 5015
rect 24041 4981 24075 5015
rect 27353 4981 27387 5015
rect 28825 4981 28859 5015
rect 29377 4981 29411 5015
rect 26985 4777 27019 4811
rect 26893 4709 26927 4743
rect 28273 4709 28307 4743
rect 26525 4641 26559 4675
rect 28733 4641 28767 4675
rect 28917 4641 28951 4675
rect 1409 4573 1443 4607
rect 23581 4573 23615 4607
rect 23857 4573 23891 4607
rect 25237 4573 25271 4607
rect 25421 4573 25455 4607
rect 25513 4573 25547 4607
rect 27813 4573 27847 4607
rect 29929 4573 29963 4607
rect 28641 4505 28675 4539
rect 1593 4437 1627 4471
rect 23397 4437 23431 4471
rect 23765 4437 23799 4471
rect 25053 4437 25087 4471
rect 27629 4437 27663 4471
rect 30021 4437 30055 4471
rect 2053 4233 2087 4267
rect 29377 4233 29411 4267
rect 22284 4165 22318 4199
rect 24194 4165 24228 4199
rect 28549 4165 28583 4199
rect 1409 4097 1443 4131
rect 16681 4097 16715 4131
rect 27445 4097 27479 4131
rect 28181 4097 28215 4131
rect 29745 4097 29779 4131
rect 22017 4029 22051 4063
rect 23949 4029 23983 4063
rect 29009 4029 29043 4063
rect 29837 4029 29871 4063
rect 29929 4029 29963 4063
rect 23397 3961 23431 3995
rect 27997 3961 28031 3995
rect 1593 3893 1627 3927
rect 16865 3893 16899 3927
rect 25329 3893 25363 3927
rect 27261 3893 27295 3927
rect 28641 3893 28675 3927
rect 28089 3621 28123 3655
rect 24869 3553 24903 3587
rect 1409 3485 1443 3519
rect 25136 3485 25170 3519
rect 28273 3485 28307 3519
rect 28733 3485 28767 3519
rect 29929 3485 29963 3519
rect 1593 3349 1627 3383
rect 26249 3349 26283 3383
rect 28917 3349 28951 3383
rect 30021 3349 30055 3383
rect 29101 3145 29135 3179
rect 29837 3145 29871 3179
rect 1409 3009 1443 3043
rect 28917 3009 28951 3043
rect 29745 3009 29779 3043
rect 1593 2805 1627 2839
rect 28089 2601 28123 2635
rect 28917 2533 28951 2567
rect 1409 2397 1443 2431
rect 2145 2397 2179 2431
rect 3065 2397 3099 2431
rect 28273 2397 28307 2431
rect 28733 2397 28767 2431
rect 29653 2397 29687 2431
rect 29929 2329 29963 2363
rect 1593 2261 1627 2295
rect 2329 2261 2363 2295
rect 2881 2261 2915 2295
<< metal1 >>
rect 1104 77818 30820 77840
rect 1104 77766 5915 77818
rect 5967 77766 5979 77818
rect 6031 77766 6043 77818
rect 6095 77766 6107 77818
rect 6159 77766 6171 77818
rect 6223 77766 15846 77818
rect 15898 77766 15910 77818
rect 15962 77766 15974 77818
rect 16026 77766 16038 77818
rect 16090 77766 16102 77818
rect 16154 77766 25776 77818
rect 25828 77766 25840 77818
rect 25892 77766 25904 77818
rect 25956 77766 25968 77818
rect 26020 77766 26032 77818
rect 26084 77766 30820 77818
rect 1104 77744 30820 77766
rect 27433 77707 27491 77713
rect 27433 77673 27445 77707
rect 27479 77704 27491 77707
rect 27890 77704 27896 77716
rect 27479 77676 27896 77704
rect 27479 77673 27491 77676
rect 27433 77667 27491 77673
rect 27890 77664 27896 77676
rect 27948 77664 27954 77716
rect 28166 77704 28172 77716
rect 28127 77676 28172 77704
rect 28166 77664 28172 77676
rect 28224 77664 28230 77716
rect 1394 77568 1400 77580
rect 1355 77540 1400 77568
rect 1394 77528 1400 77540
rect 1452 77528 1458 77580
rect 3786 77568 3792 77580
rect 3747 77540 3792 77568
rect 3786 77528 3792 77540
rect 3844 77528 3850 77580
rect 1673 77503 1731 77509
rect 1673 77469 1685 77503
rect 1719 77469 1731 77503
rect 1673 77463 1731 77469
rect 4065 77503 4123 77509
rect 4065 77469 4077 77503
rect 4111 77500 4123 77503
rect 11698 77500 11704 77512
rect 4111 77472 11704 77500
rect 4111 77469 4123 77472
rect 4065 77463 4123 77469
rect 1688 77364 1716 77463
rect 11698 77460 11704 77472
rect 11756 77460 11762 77512
rect 27246 77500 27252 77512
rect 27207 77472 27252 77500
rect 27246 77460 27252 77472
rect 27304 77460 27310 77512
rect 27706 77460 27712 77512
rect 27764 77500 27770 77512
rect 27985 77503 28043 77509
rect 27985 77500 27997 77503
rect 27764 77472 27997 77500
rect 27764 77460 27770 77472
rect 27985 77469 27997 77472
rect 28031 77469 28043 77503
rect 27985 77463 28043 77469
rect 28721 77503 28779 77509
rect 28721 77469 28733 77503
rect 28767 77469 28779 77503
rect 28721 77463 28779 77469
rect 27154 77392 27160 77444
rect 27212 77432 27218 77444
rect 28736 77432 28764 77463
rect 29362 77460 29368 77512
rect 29420 77500 29426 77512
rect 29825 77503 29883 77509
rect 29825 77500 29837 77503
rect 29420 77472 29837 77500
rect 29420 77460 29426 77472
rect 29825 77469 29837 77472
rect 29871 77469 29883 77503
rect 29825 77463 29883 77469
rect 27212 77404 28764 77432
rect 27212 77392 27218 77404
rect 11790 77364 11796 77376
rect 1688 77336 11796 77364
rect 11790 77324 11796 77336
rect 11848 77324 11854 77376
rect 28902 77364 28908 77376
rect 28863 77336 28908 77364
rect 28902 77324 28908 77336
rect 28960 77324 28966 77376
rect 30009 77367 30067 77373
rect 30009 77333 30021 77367
rect 30055 77364 30067 77367
rect 30098 77364 30104 77376
rect 30055 77336 30104 77364
rect 30055 77333 30067 77336
rect 30009 77327 30067 77333
rect 30098 77324 30104 77336
rect 30156 77324 30162 77376
rect 1104 77274 30820 77296
rect 1104 77222 10880 77274
rect 10932 77222 10944 77274
rect 10996 77222 11008 77274
rect 11060 77222 11072 77274
rect 11124 77222 11136 77274
rect 11188 77222 20811 77274
rect 20863 77222 20875 77274
rect 20927 77222 20939 77274
rect 20991 77222 21003 77274
rect 21055 77222 21067 77274
rect 21119 77222 30820 77274
rect 1104 77200 30820 77222
rect 28534 77160 28540 77172
rect 28495 77132 28540 77160
rect 28534 77120 28540 77132
rect 28592 77120 28598 77172
rect 29270 77160 29276 77172
rect 29231 77132 29276 77160
rect 29270 77120 29276 77132
rect 29328 77120 29334 77172
rect 2685 77027 2743 77033
rect 2685 76993 2697 77027
rect 2731 77024 2743 77027
rect 2774 77024 2780 77036
rect 2731 76996 2780 77024
rect 2731 76993 2743 76996
rect 2685 76987 2743 76993
rect 2774 76984 2780 76996
rect 2832 76984 2838 77036
rect 28350 77024 28356 77036
rect 28311 76996 28356 77024
rect 28350 76984 28356 76996
rect 28408 76984 28414 77036
rect 29086 77024 29092 77036
rect 29047 76996 29092 77024
rect 29086 76984 29092 76996
rect 29144 76984 29150 77036
rect 29825 77027 29883 77033
rect 29825 76993 29837 77027
rect 29871 76993 29883 77027
rect 29825 76987 29883 76993
rect 1394 76956 1400 76968
rect 1355 76928 1400 76956
rect 1394 76916 1400 76928
rect 1452 76916 1458 76968
rect 1673 76959 1731 76965
rect 1673 76925 1685 76959
rect 1719 76925 1731 76959
rect 1673 76919 1731 76925
rect 2961 76959 3019 76965
rect 2961 76925 2973 76959
rect 3007 76956 3019 76959
rect 13722 76956 13728 76968
rect 3007 76928 13728 76956
rect 3007 76925 3019 76928
rect 2961 76919 3019 76925
rect 1688 76888 1716 76919
rect 13722 76916 13728 76928
rect 13780 76916 13786 76968
rect 28994 76916 29000 76968
rect 29052 76956 29058 76968
rect 29840 76956 29868 76987
rect 29052 76928 29868 76956
rect 29052 76916 29058 76928
rect 8294 76888 8300 76900
rect 1688 76860 8300 76888
rect 8294 76848 8300 76860
rect 8352 76848 8358 76900
rect 30006 76820 30012 76832
rect 29967 76792 30012 76820
rect 30006 76780 30012 76792
rect 30064 76780 30070 76832
rect 1104 76730 30820 76752
rect 1104 76678 5915 76730
rect 5967 76678 5979 76730
rect 6031 76678 6043 76730
rect 6095 76678 6107 76730
rect 6159 76678 6171 76730
rect 6223 76678 15846 76730
rect 15898 76678 15910 76730
rect 15962 76678 15974 76730
rect 16026 76678 16038 76730
rect 16090 76678 16102 76730
rect 16154 76678 25776 76730
rect 25828 76678 25840 76730
rect 25892 76678 25904 76730
rect 25956 76678 25968 76730
rect 26020 76678 26032 76730
rect 26084 76678 30820 76730
rect 1104 76656 30820 76678
rect 28810 76576 28816 76628
rect 28868 76616 28874 76628
rect 28905 76619 28963 76625
rect 28905 76616 28917 76619
rect 28868 76588 28917 76616
rect 28868 76576 28874 76588
rect 28905 76585 28917 76588
rect 28951 76585 28963 76619
rect 28905 76579 28963 76585
rect 1302 76440 1308 76492
rect 1360 76480 1366 76492
rect 1397 76483 1455 76489
rect 1397 76480 1409 76483
rect 1360 76452 1409 76480
rect 1360 76440 1366 76452
rect 1397 76449 1409 76452
rect 1443 76449 1455 76483
rect 1397 76443 1455 76449
rect 1673 76415 1731 76421
rect 1673 76381 1685 76415
rect 1719 76381 1731 76415
rect 2866 76412 2872 76424
rect 2827 76384 2872 76412
rect 1673 76375 1731 76381
rect 1688 76344 1716 76375
rect 2866 76372 2872 76384
rect 2924 76372 2930 76424
rect 26326 76372 26332 76424
rect 26384 76412 26390 76424
rect 28721 76415 28779 76421
rect 28721 76412 28733 76415
rect 26384 76384 28733 76412
rect 26384 76372 26390 76384
rect 28721 76381 28733 76384
rect 28767 76381 28779 76415
rect 28721 76375 28779 76381
rect 29730 76372 29736 76424
rect 29788 76412 29794 76424
rect 29825 76415 29883 76421
rect 29825 76412 29837 76415
rect 29788 76384 29837 76412
rect 29788 76372 29794 76384
rect 29825 76381 29837 76384
rect 29871 76381 29883 76415
rect 29825 76375 29883 76381
rect 10778 76344 10784 76356
rect 1688 76316 10784 76344
rect 10778 76304 10784 76316
rect 10836 76304 10842 76356
rect 2685 76279 2743 76285
rect 2685 76245 2697 76279
rect 2731 76276 2743 76279
rect 14642 76276 14648 76288
rect 2731 76248 14648 76276
rect 2731 76245 2743 76248
rect 2685 76239 2743 76245
rect 14642 76236 14648 76248
rect 14700 76236 14706 76288
rect 19978 76236 19984 76288
rect 20036 76276 20042 76288
rect 21174 76276 21180 76288
rect 20036 76248 21180 76276
rect 20036 76236 20042 76248
rect 21174 76236 21180 76248
rect 21232 76236 21238 76288
rect 30009 76279 30067 76285
rect 30009 76245 30021 76279
rect 30055 76276 30067 76279
rect 30190 76276 30196 76288
rect 30055 76248 30196 76276
rect 30055 76245 30067 76248
rect 30009 76239 30067 76245
rect 30190 76236 30196 76248
rect 30248 76236 30254 76288
rect 1104 76186 30820 76208
rect 1104 76134 10880 76186
rect 10932 76134 10944 76186
rect 10996 76134 11008 76186
rect 11060 76134 11072 76186
rect 11124 76134 11136 76186
rect 11188 76134 20811 76186
rect 20863 76134 20875 76186
rect 20927 76134 20939 76186
rect 20991 76134 21003 76186
rect 21055 76134 21067 76186
rect 21119 76134 30820 76186
rect 1104 76112 30820 76134
rect 1397 76075 1455 76081
rect 1397 76041 1409 76075
rect 1443 76072 1455 76075
rect 14550 76072 14556 76084
rect 1443 76044 14556 76072
rect 1443 76041 1455 76044
rect 1397 76035 1455 76041
rect 14550 76032 14556 76044
rect 14608 76032 14614 76084
rect 29270 76072 29276 76084
rect 29231 76044 29276 76072
rect 29270 76032 29276 76044
rect 29328 76032 29334 76084
rect 14642 76004 14648 76016
rect 14603 75976 14648 76004
rect 14642 75964 14648 75976
rect 14700 75964 14706 76016
rect 15286 75964 15292 76016
rect 15344 76004 15350 76016
rect 30098 76004 30104 76016
rect 15344 75976 20392 76004
rect 15344 75964 15350 75976
rect 1578 75936 1584 75948
rect 1539 75908 1584 75936
rect 1578 75896 1584 75908
rect 1636 75896 1642 75948
rect 14458 75936 14464 75948
rect 14419 75908 14464 75936
rect 14458 75896 14464 75908
rect 14516 75896 14522 75948
rect 15746 75896 15752 75948
rect 15804 75936 15810 75948
rect 15841 75939 15899 75945
rect 15841 75936 15853 75939
rect 15804 75908 15853 75936
rect 15804 75896 15810 75908
rect 15841 75905 15853 75908
rect 15887 75905 15899 75939
rect 15841 75899 15899 75905
rect 16758 75896 16764 75948
rect 16816 75936 16822 75948
rect 16853 75939 16911 75945
rect 16853 75936 16865 75939
rect 16816 75908 16865 75936
rect 16816 75896 16822 75908
rect 16853 75905 16865 75908
rect 16899 75905 16911 75939
rect 19058 75936 19064 75948
rect 19019 75908 19064 75936
rect 16853 75899 16911 75905
rect 19058 75896 19064 75908
rect 19116 75896 19122 75948
rect 19978 75936 19984 75948
rect 19939 75908 19984 75936
rect 19978 75896 19984 75908
rect 20036 75896 20042 75948
rect 20073 75939 20131 75945
rect 20073 75905 20085 75939
rect 20119 75905 20131 75939
rect 20073 75899 20131 75905
rect 20088 75868 20116 75899
rect 20162 75896 20168 75948
rect 20220 75936 20226 75948
rect 20364 75945 20392 75976
rect 29104 75976 30104 76004
rect 29104 75945 29132 75976
rect 30098 75964 30104 75976
rect 30156 75964 30162 76016
rect 20349 75939 20407 75945
rect 20220 75908 20265 75936
rect 20220 75896 20226 75908
rect 20349 75905 20361 75939
rect 20395 75905 20407 75939
rect 20349 75899 20407 75905
rect 29089 75939 29147 75945
rect 29089 75905 29101 75939
rect 29135 75905 29147 75939
rect 29822 75936 29828 75948
rect 29783 75908 29828 75936
rect 29089 75899 29147 75905
rect 29822 75896 29828 75908
rect 29880 75896 29886 75948
rect 21542 75868 21548 75880
rect 20088 75840 21548 75868
rect 21542 75828 21548 75840
rect 21600 75828 21606 75880
rect 14829 75803 14887 75809
rect 14829 75769 14841 75803
rect 14875 75800 14887 75803
rect 19886 75800 19892 75812
rect 14875 75772 19892 75800
rect 14875 75769 14887 75772
rect 14829 75763 14887 75769
rect 19886 75760 19892 75772
rect 19944 75760 19950 75812
rect 15194 75692 15200 75744
rect 15252 75732 15258 75744
rect 16025 75735 16083 75741
rect 16025 75732 16037 75735
rect 15252 75704 16037 75732
rect 15252 75692 15258 75704
rect 16025 75701 16037 75704
rect 16071 75701 16083 75735
rect 17034 75732 17040 75744
rect 16995 75704 17040 75732
rect 16025 75695 16083 75701
rect 17034 75692 17040 75704
rect 17092 75692 17098 75744
rect 19245 75735 19303 75741
rect 19245 75701 19257 75735
rect 19291 75732 19303 75735
rect 19610 75732 19616 75744
rect 19291 75704 19616 75732
rect 19291 75701 19303 75704
rect 19245 75695 19303 75701
rect 19610 75692 19616 75704
rect 19668 75692 19674 75744
rect 19702 75692 19708 75744
rect 19760 75732 19766 75744
rect 30006 75732 30012 75744
rect 19760 75704 19805 75732
rect 29967 75704 30012 75732
rect 19760 75692 19766 75704
rect 30006 75692 30012 75704
rect 30064 75692 30070 75744
rect 1104 75642 30820 75664
rect 1104 75590 5915 75642
rect 5967 75590 5979 75642
rect 6031 75590 6043 75642
rect 6095 75590 6107 75642
rect 6159 75590 6171 75642
rect 6223 75590 15846 75642
rect 15898 75590 15910 75642
rect 15962 75590 15974 75642
rect 16026 75590 16038 75642
rect 16090 75590 16102 75642
rect 16154 75590 25776 75642
rect 25828 75590 25840 75642
rect 25892 75590 25904 75642
rect 25956 75590 25968 75642
rect 26020 75590 26032 75642
rect 26084 75590 30820 75642
rect 1104 75568 30820 75590
rect 14737 75531 14795 75537
rect 14737 75497 14749 75531
rect 14783 75528 14795 75531
rect 21174 75528 21180 75540
rect 14783 75500 20751 75528
rect 21135 75500 21180 75528
rect 14783 75497 14795 75500
rect 14737 75491 14795 75497
rect 20723 75460 20751 75500
rect 21174 75488 21180 75500
rect 21232 75488 21238 75540
rect 22370 75460 22376 75472
rect 20723 75432 22376 75460
rect 22370 75420 22376 75432
rect 22428 75420 22434 75472
rect 15194 75392 15200 75404
rect 15155 75364 15200 75392
rect 15194 75352 15200 75364
rect 15252 75352 15258 75404
rect 17034 75352 17040 75404
rect 17092 75392 17098 75404
rect 17129 75395 17187 75401
rect 17129 75392 17141 75395
rect 17092 75364 17141 75392
rect 17092 75352 17098 75364
rect 17129 75361 17141 75364
rect 17175 75361 17187 75395
rect 17129 75355 17187 75361
rect 19610 75352 19616 75404
rect 19668 75392 19674 75404
rect 19797 75395 19855 75401
rect 19797 75392 19809 75395
rect 19668 75364 19809 75392
rect 19668 75352 19674 75364
rect 19797 75361 19809 75364
rect 19843 75361 19855 75395
rect 19797 75355 19855 75361
rect 1578 75324 1584 75336
rect 1539 75296 1584 75324
rect 1578 75284 1584 75296
rect 1636 75284 1642 75336
rect 14550 75324 14556 75336
rect 14511 75296 14556 75324
rect 14550 75284 14556 75296
rect 14608 75284 14614 75336
rect 19702 75284 19708 75336
rect 19760 75324 19766 75336
rect 20053 75327 20111 75333
rect 20053 75324 20065 75327
rect 19760 75296 20065 75324
rect 19760 75284 19766 75296
rect 20053 75293 20065 75296
rect 20099 75293 20111 75327
rect 20053 75287 20111 75293
rect 29825 75327 29883 75333
rect 29825 75293 29837 75327
rect 29871 75324 29883 75327
rect 29914 75324 29920 75336
rect 29871 75296 29920 75324
rect 29871 75293 29883 75296
rect 29825 75287 29883 75293
rect 29914 75284 29920 75296
rect 29972 75284 29978 75336
rect 14369 75259 14427 75265
rect 14369 75225 14381 75259
rect 14415 75256 14427 75259
rect 14458 75256 14464 75268
rect 14415 75228 14464 75256
rect 14415 75225 14427 75228
rect 14369 75219 14427 75225
rect 14458 75216 14464 75228
rect 14516 75216 14522 75268
rect 15464 75259 15522 75265
rect 15464 75225 15476 75259
rect 15510 75256 15522 75259
rect 16666 75256 16672 75268
rect 15510 75228 16672 75256
rect 15510 75225 15522 75228
rect 15464 75219 15522 75225
rect 16666 75216 16672 75228
rect 16724 75216 16730 75268
rect 16850 75216 16856 75268
rect 16908 75256 16914 75268
rect 17374 75259 17432 75265
rect 17374 75256 17386 75259
rect 16908 75228 17386 75256
rect 16908 75216 16914 75228
rect 17374 75225 17386 75228
rect 17420 75225 17432 75259
rect 17374 75219 17432 75225
rect 19886 75216 19892 75268
rect 19944 75256 19950 75268
rect 21266 75256 21272 75268
rect 19944 75228 21272 75256
rect 19944 75216 19950 75228
rect 21266 75216 21272 75228
rect 21324 75216 21330 75268
rect 1397 75191 1455 75197
rect 1397 75157 1409 75191
rect 1443 75188 1455 75191
rect 14642 75188 14648 75200
rect 1443 75160 14648 75188
rect 1443 75157 1455 75160
rect 1397 75151 1455 75157
rect 14642 75148 14648 75160
rect 14700 75148 14706 75200
rect 16577 75191 16635 75197
rect 16577 75157 16589 75191
rect 16623 75188 16635 75191
rect 16942 75188 16948 75200
rect 16623 75160 16948 75188
rect 16623 75157 16635 75160
rect 16577 75151 16635 75157
rect 16942 75148 16948 75160
rect 17000 75148 17006 75200
rect 17034 75148 17040 75200
rect 17092 75188 17098 75200
rect 18509 75191 18567 75197
rect 18509 75188 18521 75191
rect 17092 75160 18521 75188
rect 17092 75148 17098 75160
rect 18509 75157 18521 75160
rect 18555 75157 18567 75191
rect 18509 75151 18567 75157
rect 21174 75148 21180 75200
rect 21232 75188 21238 75200
rect 24946 75188 24952 75200
rect 21232 75160 24952 75188
rect 21232 75148 21238 75160
rect 24946 75148 24952 75160
rect 25004 75148 25010 75200
rect 30009 75191 30067 75197
rect 30009 75157 30021 75191
rect 30055 75188 30067 75191
rect 30190 75188 30196 75200
rect 30055 75160 30196 75188
rect 30055 75157 30067 75160
rect 30009 75151 30067 75157
rect 30190 75148 30196 75160
rect 30248 75148 30254 75200
rect 1104 75098 30820 75120
rect 1104 75046 10880 75098
rect 10932 75046 10944 75098
rect 10996 75046 11008 75098
rect 11060 75046 11072 75098
rect 11124 75046 11136 75098
rect 11188 75046 20811 75098
rect 20863 75046 20875 75098
rect 20927 75046 20939 75098
rect 20991 75046 21003 75098
rect 21055 75046 21067 75098
rect 21119 75046 30820 75098
rect 1104 75024 30820 75046
rect 14829 74987 14887 74993
rect 14829 74953 14841 74987
rect 14875 74984 14887 74987
rect 15286 74984 15292 74996
rect 14875 74956 15292 74984
rect 14875 74953 14887 74956
rect 14829 74947 14887 74953
rect 15286 74944 15292 74956
rect 15344 74944 15350 74996
rect 15657 74987 15715 74993
rect 15657 74953 15669 74987
rect 15703 74984 15715 74987
rect 21450 74984 21456 74996
rect 15703 74956 21456 74984
rect 15703 74953 15715 74956
rect 15657 74947 15715 74953
rect 21450 74944 21456 74956
rect 21508 74944 21514 74996
rect 14642 74916 14648 74928
rect 14603 74888 14648 74916
rect 14642 74876 14648 74888
rect 14700 74876 14706 74928
rect 17218 74916 17224 74928
rect 17179 74888 17224 74916
rect 17218 74876 17224 74888
rect 17276 74876 17282 74928
rect 20162 74876 20168 74928
rect 20220 74916 20226 74928
rect 20714 74916 20720 74928
rect 20220 74888 20720 74916
rect 20220 74876 20226 74888
rect 20714 74876 20720 74888
rect 20772 74916 20778 74928
rect 20772 74888 21128 74916
rect 20772 74876 20778 74888
rect 1578 74848 1584 74860
rect 1539 74820 1584 74848
rect 1578 74808 1584 74820
rect 1636 74808 1642 74860
rect 14461 74851 14519 74857
rect 14461 74817 14473 74851
rect 14507 74848 14519 74851
rect 14550 74848 14556 74860
rect 14507 74820 14556 74848
rect 14507 74817 14519 74820
rect 14461 74811 14519 74817
rect 14550 74808 14556 74820
rect 14608 74848 14614 74860
rect 15289 74851 15347 74857
rect 15289 74848 15301 74851
rect 14608 74820 15301 74848
rect 14608 74808 14614 74820
rect 15289 74817 15301 74820
rect 15335 74817 15347 74851
rect 15289 74811 15347 74817
rect 15473 74851 15531 74857
rect 15473 74817 15485 74851
rect 15519 74817 15531 74851
rect 15473 74811 15531 74817
rect 1397 74715 1455 74721
rect 1397 74681 1409 74715
rect 1443 74712 1455 74715
rect 15488 74712 15516 74811
rect 16482 74808 16488 74860
rect 16540 74848 16546 74860
rect 17037 74851 17095 74857
rect 17037 74848 17049 74851
rect 16540 74820 17049 74848
rect 16540 74808 16546 74820
rect 17037 74817 17049 74820
rect 17083 74817 17095 74851
rect 17037 74811 17095 74817
rect 17954 74808 17960 74860
rect 18012 74848 18018 74860
rect 21100 74857 21128 74888
rect 18489 74851 18547 74857
rect 18489 74848 18501 74851
rect 18012 74820 18501 74848
rect 18012 74808 18018 74820
rect 18489 74817 18501 74820
rect 18535 74817 18547 74851
rect 18489 74811 18547 74817
rect 20901 74851 20959 74857
rect 20901 74817 20913 74851
rect 20947 74817 20959 74851
rect 20901 74811 20959 74817
rect 20993 74851 21051 74857
rect 20993 74817 21005 74851
rect 21039 74817 21051 74851
rect 20993 74811 21051 74817
rect 21085 74851 21143 74857
rect 21085 74817 21097 74851
rect 21131 74817 21143 74851
rect 21266 74848 21272 74860
rect 21227 74820 21272 74848
rect 21085 74811 21143 74817
rect 16574 74740 16580 74792
rect 16632 74780 16638 74792
rect 17313 74783 17371 74789
rect 17313 74780 17325 74783
rect 16632 74752 17325 74780
rect 16632 74740 16638 74752
rect 17313 74749 17325 74752
rect 17359 74749 17371 74783
rect 18230 74780 18236 74792
rect 18191 74752 18236 74780
rect 17313 74743 17371 74749
rect 18230 74740 18236 74752
rect 18288 74740 18294 74792
rect 16758 74712 16764 74724
rect 1443 74684 15516 74712
rect 16719 74684 16764 74712
rect 1443 74681 1455 74684
rect 1397 74675 1455 74681
rect 16758 74672 16764 74684
rect 16816 74672 16822 74724
rect 20916 74712 20944 74811
rect 21008 74780 21036 74811
rect 21266 74808 21272 74820
rect 21324 74808 21330 74860
rect 21358 74808 21364 74860
rect 21416 74848 21422 74860
rect 22077 74851 22135 74857
rect 22077 74848 22089 74851
rect 21416 74820 22089 74848
rect 21416 74808 21422 74820
rect 22077 74817 22089 74820
rect 22123 74817 22135 74851
rect 22077 74811 22135 74817
rect 27430 74808 27436 74860
rect 27488 74848 27494 74860
rect 29825 74851 29883 74857
rect 29825 74848 29837 74851
rect 27488 74820 29837 74848
rect 27488 74808 27494 74820
rect 29825 74817 29837 74820
rect 29871 74817 29883 74851
rect 29825 74811 29883 74817
rect 21542 74780 21548 74792
rect 21008 74752 21548 74780
rect 21542 74740 21548 74752
rect 21600 74740 21606 74792
rect 21818 74780 21824 74792
rect 21779 74752 21824 74780
rect 21818 74740 21824 74752
rect 21876 74740 21882 74792
rect 20916 74684 21496 74712
rect 19613 74647 19671 74653
rect 19613 74613 19625 74647
rect 19659 74644 19671 74647
rect 20070 74644 20076 74656
rect 19659 74616 20076 74644
rect 19659 74613 19671 74616
rect 19613 74607 19671 74613
rect 20070 74604 20076 74616
rect 20128 74604 20134 74656
rect 20625 74647 20683 74653
rect 20625 74613 20637 74647
rect 20671 74644 20683 74647
rect 21266 74644 21272 74656
rect 20671 74616 21272 74644
rect 20671 74613 20683 74616
rect 20625 74607 20683 74613
rect 21266 74604 21272 74616
rect 21324 74604 21330 74656
rect 21468 74644 21496 74684
rect 22554 74644 22560 74656
rect 21468 74616 22560 74644
rect 22554 74604 22560 74616
rect 22612 74604 22618 74656
rect 22830 74604 22836 74656
rect 22888 74644 22894 74656
rect 23201 74647 23259 74653
rect 23201 74644 23213 74647
rect 22888 74616 23213 74644
rect 22888 74604 22894 74616
rect 23201 74613 23213 74616
rect 23247 74613 23259 74647
rect 30006 74644 30012 74656
rect 29967 74616 30012 74644
rect 23201 74607 23259 74613
rect 30006 74604 30012 74616
rect 30064 74604 30070 74656
rect 1104 74554 30820 74576
rect 1104 74502 5915 74554
rect 5967 74502 5979 74554
rect 6031 74502 6043 74554
rect 6095 74502 6107 74554
rect 6159 74502 6171 74554
rect 6223 74502 15846 74554
rect 15898 74502 15910 74554
rect 15962 74502 15974 74554
rect 16026 74502 16038 74554
rect 16090 74502 16102 74554
rect 16154 74502 25776 74554
rect 25828 74502 25840 74554
rect 25892 74502 25904 74554
rect 25956 74502 25968 74554
rect 26020 74502 26032 74554
rect 26084 74502 30820 74554
rect 1104 74480 30820 74502
rect 15746 74400 15752 74452
rect 15804 74440 15810 74452
rect 16025 74443 16083 74449
rect 16025 74440 16037 74443
rect 15804 74412 16037 74440
rect 15804 74400 15810 74412
rect 16025 74409 16037 74412
rect 16071 74409 16083 74443
rect 16025 74403 16083 74409
rect 17497 74443 17555 74449
rect 17497 74409 17509 74443
rect 17543 74440 17555 74443
rect 18230 74440 18236 74452
rect 17543 74412 18236 74440
rect 17543 74409 17555 74412
rect 17497 74403 17555 74409
rect 18230 74400 18236 74412
rect 18288 74400 18294 74452
rect 19886 74440 19892 74452
rect 19260 74412 19892 74440
rect 14921 74375 14979 74381
rect 14921 74341 14933 74375
rect 14967 74372 14979 74375
rect 18049 74375 18107 74381
rect 14967 74344 18000 74372
rect 14967 74341 14979 74344
rect 14921 74335 14979 74341
rect 16482 74304 16488 74316
rect 16443 74276 16488 74304
rect 16482 74264 16488 74276
rect 16540 74264 16546 74316
rect 17972 74304 18000 74344
rect 18049 74341 18061 74375
rect 18095 74372 18107 74375
rect 19058 74372 19064 74384
rect 18095 74344 19064 74372
rect 18095 74341 18107 74344
rect 18049 74335 18107 74341
rect 19058 74332 19064 74344
rect 19116 74332 19122 74384
rect 18414 74304 18420 74316
rect 17972 74276 18420 74304
rect 18414 74264 18420 74276
rect 18472 74264 18478 74316
rect 18601 74307 18659 74313
rect 18601 74273 18613 74307
rect 18647 74304 18659 74307
rect 19260 74304 19288 74412
rect 19886 74400 19892 74412
rect 19944 74400 19950 74452
rect 20625 74443 20683 74449
rect 20625 74409 20637 74443
rect 20671 74440 20683 74443
rect 21818 74440 21824 74452
rect 20671 74412 21824 74440
rect 20671 74409 20683 74412
rect 20625 74403 20683 74409
rect 21818 74400 21824 74412
rect 21876 74400 21882 74452
rect 19337 74375 19395 74381
rect 19337 74341 19349 74375
rect 19383 74341 19395 74375
rect 19337 74335 19395 74341
rect 18647 74276 19288 74304
rect 18647 74273 18659 74276
rect 18601 74267 18659 74273
rect 17313 74239 17371 74245
rect 17313 74205 17325 74239
rect 17359 74236 17371 74239
rect 19352 74236 19380 74335
rect 20438 74236 20444 74248
rect 17359 74208 19380 74236
rect 20399 74208 20444 74236
rect 17359 74205 17371 74208
rect 17313 74199 17371 74205
rect 20438 74196 20444 74208
rect 20496 74196 20502 74248
rect 21174 74236 21180 74248
rect 21135 74208 21180 74236
rect 21174 74196 21180 74208
rect 21232 74196 21238 74248
rect 21266 74196 21272 74248
rect 21324 74236 21330 74248
rect 21433 74239 21491 74245
rect 21433 74236 21445 74239
rect 21324 74208 21445 74236
rect 21324 74196 21330 74208
rect 21433 74205 21445 74208
rect 21479 74205 21491 74239
rect 21433 74199 21491 74205
rect 26234 74196 26240 74248
rect 26292 74236 26298 74248
rect 29825 74239 29883 74245
rect 29825 74236 29837 74239
rect 26292 74208 29837 74236
rect 26292 74196 26298 74208
rect 29825 74205 29837 74208
rect 29871 74205 29883 74239
rect 29825 74199 29883 74205
rect 14550 74168 14556 74180
rect 14511 74140 14556 74168
rect 14550 74128 14556 74140
rect 14608 74128 14614 74180
rect 14734 74168 14740 74180
rect 14695 74140 14740 74168
rect 14734 74128 14740 74140
rect 14792 74128 14798 74180
rect 16574 74168 16580 74180
rect 16535 74140 16580 74168
rect 16574 74128 16580 74140
rect 16632 74128 16638 74180
rect 18325 74171 18383 74177
rect 18325 74137 18337 74171
rect 18371 74168 18383 74171
rect 19518 74168 19524 74180
rect 18371 74140 19524 74168
rect 18371 74137 18383 74140
rect 18325 74131 18383 74137
rect 19518 74128 19524 74140
rect 19576 74168 19582 74180
rect 19613 74171 19671 74177
rect 19613 74168 19625 74171
rect 19576 74140 19625 74168
rect 19576 74128 19582 74140
rect 19613 74137 19625 74140
rect 19659 74137 19671 74171
rect 19886 74168 19892 74180
rect 19847 74140 19892 74168
rect 19613 74131 19671 74137
rect 19886 74128 19892 74140
rect 19944 74128 19950 74180
rect 16485 74103 16543 74109
rect 16485 74069 16497 74103
rect 16531 74100 16543 74103
rect 17218 74100 17224 74112
rect 16531 74072 17224 74100
rect 16531 74069 16543 74072
rect 16485 74063 16543 74069
rect 17218 74060 17224 74072
rect 17276 74060 17282 74112
rect 18509 74103 18567 74109
rect 18509 74069 18521 74103
rect 18555 74100 18567 74103
rect 19702 74100 19708 74112
rect 18555 74072 19708 74100
rect 18555 74069 18567 74072
rect 18509 74063 18567 74069
rect 19702 74060 19708 74072
rect 19760 74100 19766 74112
rect 19797 74103 19855 74109
rect 19797 74100 19809 74103
rect 19760 74072 19809 74100
rect 19760 74060 19766 74072
rect 19797 74069 19809 74072
rect 19843 74069 19855 74103
rect 19797 74063 19855 74069
rect 22557 74103 22615 74109
rect 22557 74069 22569 74103
rect 22603 74100 22615 74103
rect 22646 74100 22652 74112
rect 22603 74072 22652 74100
rect 22603 74069 22615 74072
rect 22557 74063 22615 74069
rect 22646 74060 22652 74072
rect 22704 74060 22710 74112
rect 30009 74103 30067 74109
rect 30009 74069 30021 74103
rect 30055 74100 30067 74103
rect 30190 74100 30196 74112
rect 30055 74072 30196 74100
rect 30055 74069 30067 74072
rect 30009 74063 30067 74069
rect 30190 74060 30196 74072
rect 30248 74060 30254 74112
rect 1104 74010 30820 74032
rect 1104 73958 10880 74010
rect 10932 73958 10944 74010
rect 10996 73958 11008 74010
rect 11060 73958 11072 74010
rect 11124 73958 11136 74010
rect 11188 73958 20811 74010
rect 20863 73958 20875 74010
rect 20927 73958 20939 74010
rect 20991 73958 21003 74010
rect 21055 73958 21067 74010
rect 21119 73958 30820 74010
rect 1104 73936 30820 73958
rect 13725 73899 13783 73905
rect 13725 73865 13737 73899
rect 13771 73896 13783 73899
rect 14550 73896 14556 73908
rect 13771 73868 14556 73896
rect 13771 73865 13783 73868
rect 13725 73859 13783 73865
rect 14550 73856 14556 73868
rect 14608 73856 14614 73908
rect 16666 73896 16672 73908
rect 16627 73868 16672 73896
rect 16666 73856 16672 73868
rect 16724 73856 16730 73908
rect 17954 73896 17960 73908
rect 17915 73868 17960 73896
rect 17954 73856 17960 73868
rect 18012 73856 18018 73908
rect 19702 73896 19708 73908
rect 19663 73868 19708 73896
rect 19702 73856 19708 73868
rect 19760 73856 19766 73908
rect 20625 73899 20683 73905
rect 20625 73865 20637 73899
rect 20671 73896 20683 73899
rect 21358 73896 21364 73908
rect 20671 73868 21364 73896
rect 20671 73865 20683 73868
rect 20625 73859 20683 73865
rect 21358 73856 21364 73868
rect 21416 73856 21422 73908
rect 17862 73828 17868 73840
rect 17052 73800 17868 73828
rect 1578 73760 1584 73772
rect 1539 73732 1584 73760
rect 1578 73720 1584 73732
rect 1636 73720 1642 73772
rect 13538 73720 13544 73772
rect 13596 73760 13602 73772
rect 13909 73763 13967 73769
rect 13909 73760 13921 73763
rect 13596 73732 13921 73760
rect 13596 73720 13602 73732
rect 13909 73729 13921 73732
rect 13955 73729 13967 73763
rect 16942 73760 16948 73772
rect 16903 73732 16948 73760
rect 13909 73723 13967 73729
rect 16942 73720 16948 73732
rect 17000 73720 17006 73772
rect 17052 73769 17080 73800
rect 17862 73788 17868 73800
rect 17920 73788 17926 73840
rect 19518 73828 19524 73840
rect 18340 73800 18736 73828
rect 19479 73800 19524 73828
rect 17037 73763 17095 73769
rect 17037 73729 17049 73763
rect 17083 73729 17095 73763
rect 17037 73723 17095 73729
rect 17129 73763 17187 73769
rect 17129 73729 17141 73763
rect 17175 73729 17187 73763
rect 17129 73723 17187 73729
rect 17325 73763 17383 73769
rect 17325 73729 17337 73763
rect 17371 73760 17383 73763
rect 17494 73760 17500 73772
rect 17371 73732 17500 73760
rect 17371 73729 17383 73732
rect 17325 73723 17383 73729
rect 17144 73692 17172 73723
rect 17494 73720 17500 73732
rect 17552 73720 17558 73772
rect 18230 73760 18236 73772
rect 18191 73732 18236 73760
rect 18230 73720 18236 73732
rect 18288 73720 18294 73772
rect 18340 73769 18368 73800
rect 18325 73763 18383 73769
rect 18325 73729 18337 73763
rect 18371 73729 18383 73763
rect 18325 73723 18383 73729
rect 18417 73763 18475 73769
rect 18417 73729 18429 73763
rect 18463 73729 18475 73763
rect 18417 73723 18475 73729
rect 18601 73763 18659 73769
rect 18601 73729 18613 73763
rect 18647 73729 18659 73763
rect 18708 73760 18736 73800
rect 19518 73788 19524 73800
rect 19576 73788 19582 73840
rect 20640 73800 21036 73828
rect 20640 73760 20668 73800
rect 21008 73769 21036 73800
rect 18708 73732 20668 73760
rect 20901 73763 20959 73769
rect 18601 73723 18659 73729
rect 20901 73729 20913 73763
rect 20947 73729 20959 73763
rect 20901 73723 20959 73729
rect 20993 73763 21051 73769
rect 20993 73729 21005 73763
rect 21039 73729 21051 73763
rect 20993 73723 21051 73729
rect 18432 73692 18460 73723
rect 17144 73664 18460 73692
rect 17328 73636 17356 73664
rect 1397 73627 1455 73633
rect 1397 73593 1409 73627
rect 1443 73624 1455 73627
rect 14734 73624 14740 73636
rect 1443 73596 14740 73624
rect 1443 73593 1455 73596
rect 1397 73587 1455 73593
rect 14734 73584 14740 73596
rect 14792 73584 14798 73636
rect 17310 73584 17316 73636
rect 17368 73584 17374 73636
rect 18414 73584 18420 73636
rect 18472 73624 18478 73636
rect 18616 73624 18644 73723
rect 19797 73695 19855 73701
rect 19797 73661 19809 73695
rect 19843 73692 19855 73695
rect 19886 73692 19892 73704
rect 19843 73664 19892 73692
rect 19843 73661 19855 73664
rect 19797 73655 19855 73661
rect 19886 73652 19892 73664
rect 19944 73652 19950 73704
rect 18472 73596 18644 73624
rect 19245 73627 19303 73633
rect 18472 73584 18478 73596
rect 19245 73593 19257 73627
rect 19291 73624 19303 73627
rect 20438 73624 20444 73636
rect 19291 73596 20444 73624
rect 19291 73593 19303 73596
rect 19245 73587 19303 73593
rect 20438 73584 20444 73596
rect 20496 73584 20502 73636
rect 18230 73516 18236 73568
rect 18288 73556 18294 73568
rect 20070 73556 20076 73568
rect 18288 73528 20076 73556
rect 18288 73516 18294 73528
rect 20070 73516 20076 73528
rect 20128 73516 20134 73568
rect 20916 73556 20944 73723
rect 21008 73692 21036 73723
rect 21082 73720 21088 73772
rect 21140 73760 21146 73772
rect 21269 73763 21327 73769
rect 21140 73732 21185 73760
rect 21140 73720 21146 73732
rect 21269 73729 21281 73763
rect 21315 73760 21327 73763
rect 21450 73760 21456 73772
rect 21315 73732 21456 73760
rect 21315 73729 21327 73732
rect 21269 73723 21327 73729
rect 21450 73720 21456 73732
rect 21508 73720 21514 73772
rect 27338 73720 27344 73772
rect 27396 73760 27402 73772
rect 29825 73763 29883 73769
rect 29825 73760 29837 73763
rect 27396 73732 29837 73760
rect 27396 73720 27402 73732
rect 29825 73729 29837 73732
rect 29871 73729 29883 73763
rect 29825 73723 29883 73729
rect 21358 73692 21364 73704
rect 21008 73664 21364 73692
rect 21358 73652 21364 73664
rect 21416 73692 21422 73704
rect 21542 73692 21548 73704
rect 21416 73664 21548 73692
rect 21416 73652 21422 73664
rect 21542 73652 21548 73664
rect 21600 73652 21606 73704
rect 22830 73556 22836 73568
rect 20916 73528 22836 73556
rect 22830 73516 22836 73528
rect 22888 73516 22894 73568
rect 30006 73556 30012 73568
rect 29967 73528 30012 73556
rect 30006 73516 30012 73528
rect 30064 73516 30070 73568
rect 1104 73466 30820 73488
rect 1104 73414 5915 73466
rect 5967 73414 5979 73466
rect 6031 73414 6043 73466
rect 6095 73414 6107 73466
rect 6159 73414 6171 73466
rect 6223 73414 15846 73466
rect 15898 73414 15910 73466
rect 15962 73414 15974 73466
rect 16026 73414 16038 73466
rect 16090 73414 16102 73466
rect 16154 73414 25776 73466
rect 25828 73414 25840 73466
rect 25892 73414 25904 73466
rect 25956 73414 25968 73466
rect 26020 73414 26032 73466
rect 26084 73414 30820 73466
rect 1104 73392 30820 73414
rect 15013 73355 15071 73361
rect 15013 73321 15025 73355
rect 15059 73352 15071 73355
rect 17494 73352 17500 73364
rect 15059 73324 17500 73352
rect 15059 73321 15071 73324
rect 15013 73315 15071 73321
rect 17494 73312 17500 73324
rect 17552 73312 17558 73364
rect 18601 73355 18659 73361
rect 18601 73321 18613 73355
rect 18647 73352 18659 73355
rect 19518 73352 19524 73364
rect 18647 73324 19524 73352
rect 18647 73321 18659 73324
rect 18601 73315 18659 73321
rect 19518 73312 19524 73324
rect 19576 73312 19582 73364
rect 19702 73312 19708 73364
rect 19760 73352 19766 73364
rect 19797 73355 19855 73361
rect 19797 73352 19809 73355
rect 19760 73324 19809 73352
rect 19760 73312 19766 73324
rect 19797 73321 19809 73324
rect 19843 73321 19855 73355
rect 19797 73315 19855 73321
rect 20717 73355 20775 73361
rect 20717 73321 20729 73355
rect 20763 73352 20775 73355
rect 21174 73352 21180 73364
rect 20763 73324 21180 73352
rect 20763 73321 20775 73324
rect 20717 73315 20775 73321
rect 21174 73312 21180 73324
rect 21232 73312 21238 73364
rect 16942 73244 16948 73296
rect 17000 73284 17006 73296
rect 17000 73256 18000 73284
rect 17000 73244 17006 73256
rect 17310 73216 17316 73228
rect 17236 73188 17316 73216
rect 1578 73148 1584 73160
rect 1539 73120 1584 73148
rect 1578 73108 1584 73120
rect 1636 73108 1642 73160
rect 15657 73151 15715 73157
rect 15657 73148 15669 73151
rect 12406 73120 15669 73148
rect 9582 73040 9588 73092
rect 9640 73080 9646 73092
rect 9640 73052 10364 73080
rect 9640 73040 9646 73052
rect 1397 73015 1455 73021
rect 1397 72981 1409 73015
rect 1443 73012 1455 73015
rect 10226 73012 10232 73024
rect 1443 72984 10232 73012
rect 1443 72981 1455 72984
rect 1397 72975 1455 72981
rect 10226 72972 10232 72984
rect 10284 72972 10290 73024
rect 10336 73012 10364 73052
rect 12406 73012 12434 73120
rect 15657 73117 15669 73120
rect 15703 73117 15715 73151
rect 15838 73148 15844 73160
rect 15799 73120 15844 73148
rect 15657 73111 15715 73117
rect 15838 73108 15844 73120
rect 15896 73108 15902 73160
rect 17236 73157 17264 73188
rect 17310 73176 17316 73188
rect 17368 73176 17374 73228
rect 17017 73151 17075 73157
rect 17017 73117 17029 73151
rect 17063 73148 17075 73151
rect 17126 73148 17184 73154
rect 17063 73117 17080 73148
rect 17017 73111 17080 73117
rect 14642 73080 14648 73092
rect 14603 73052 14648 73080
rect 14642 73040 14648 73052
rect 14700 73040 14706 73092
rect 14734 73040 14740 73092
rect 14792 73080 14798 73092
rect 14829 73083 14887 73089
rect 14829 73080 14841 73083
rect 14792 73052 14841 73080
rect 14792 73040 14798 73052
rect 14829 73049 14841 73052
rect 14875 73049 14887 73083
rect 14829 73043 14887 73049
rect 14918 73040 14924 73092
rect 14976 73080 14982 73092
rect 15473 73083 15531 73089
rect 15473 73080 15485 73083
rect 14976 73052 15485 73080
rect 14976 73040 14982 73052
rect 15473 73049 15485 73052
rect 15519 73049 15531 73083
rect 15473 73043 15531 73049
rect 16761 73083 16819 73089
rect 16761 73049 16773 73083
rect 16807 73080 16819 73083
rect 16850 73080 16856 73092
rect 16807 73052 16856 73080
rect 16807 73049 16819 73052
rect 16761 73043 16819 73049
rect 16850 73040 16856 73052
rect 16908 73040 16914 73092
rect 17052 73024 17080 73111
rect 17126 73114 17138 73148
rect 17172 73114 17184 73148
rect 17126 73108 17184 73114
rect 17221 73151 17279 73157
rect 17221 73117 17233 73151
rect 17267 73117 17279 73151
rect 17221 73111 17279 73117
rect 17402 73108 17408 73160
rect 17460 73148 17466 73160
rect 17972 73148 18000 73256
rect 20530 73148 20536 73160
rect 17460 73120 17505 73148
rect 17972 73120 19840 73148
rect 20491 73120 20536 73148
rect 17460 73108 17466 73120
rect 17141 73080 17169 73108
rect 18509 73083 18567 73089
rect 17141 73052 17172 73080
rect 10336 72984 12434 73012
rect 17034 72972 17040 73024
rect 17092 72972 17098 73024
rect 17144 73012 17172 73052
rect 18509 73049 18521 73083
rect 18555 73049 18567 73083
rect 19702 73080 19708 73092
rect 19663 73052 19708 73080
rect 18509 73043 18567 73049
rect 17862 73012 17868 73024
rect 17144 72984 17868 73012
rect 17862 72972 17868 72984
rect 17920 72972 17926 73024
rect 18524 73012 18552 73043
rect 19702 73040 19708 73052
rect 19760 73040 19766 73092
rect 19812 73080 19840 73120
rect 20530 73108 20536 73120
rect 20588 73108 20594 73160
rect 26786 73108 26792 73160
rect 26844 73148 26850 73160
rect 29825 73151 29883 73157
rect 29825 73148 29837 73151
rect 26844 73120 29837 73148
rect 26844 73108 26850 73120
rect 29825 73117 29837 73120
rect 29871 73117 29883 73151
rect 29825 73111 29883 73117
rect 26142 73080 26148 73092
rect 19812 73052 26148 73080
rect 26142 73040 26148 73052
rect 26200 73040 26206 73092
rect 20714 73012 20720 73024
rect 18524 72984 20720 73012
rect 20714 72972 20720 72984
rect 20772 72972 20778 73024
rect 30006 73012 30012 73024
rect 29967 72984 30012 73012
rect 30006 72972 30012 72984
rect 30064 72972 30070 73024
rect 1104 72922 30820 72944
rect 1104 72870 10880 72922
rect 10932 72870 10944 72922
rect 10996 72870 11008 72922
rect 11060 72870 11072 72922
rect 11124 72870 11136 72922
rect 11188 72870 20811 72922
rect 20863 72870 20875 72922
rect 20927 72870 20939 72922
rect 20991 72870 21003 72922
rect 21055 72870 21067 72922
rect 21119 72870 30820 72922
rect 1104 72848 30820 72870
rect 10226 72700 10232 72752
rect 10284 72740 10290 72752
rect 14829 72743 14887 72749
rect 14829 72740 14841 72743
rect 10284 72712 14841 72740
rect 10284 72700 10290 72712
rect 14829 72709 14841 72712
rect 14875 72709 14887 72743
rect 14829 72703 14887 72709
rect 16117 72743 16175 72749
rect 16117 72709 16129 72743
rect 16163 72740 16175 72743
rect 16482 72740 16488 72752
rect 16163 72712 16488 72740
rect 16163 72709 16175 72712
rect 16117 72703 16175 72709
rect 16482 72700 16488 72712
rect 16540 72700 16546 72752
rect 1578 72672 1584 72684
rect 1539 72644 1584 72672
rect 1578 72632 1584 72644
rect 1636 72632 1642 72684
rect 14642 72672 14648 72684
rect 14555 72644 14648 72672
rect 14642 72632 14648 72644
rect 14700 72672 14706 72684
rect 14918 72672 14924 72684
rect 14700 72644 14924 72672
rect 14700 72632 14706 72644
rect 14918 72632 14924 72644
rect 14976 72632 14982 72684
rect 15933 72675 15991 72681
rect 15933 72641 15945 72675
rect 15979 72641 15991 72675
rect 17126 72672 17132 72684
rect 17087 72644 17132 72672
rect 15933 72635 15991 72641
rect 15948 72604 15976 72635
rect 17126 72632 17132 72644
rect 17184 72632 17190 72684
rect 29638 72632 29644 72684
rect 29696 72672 29702 72684
rect 29825 72675 29883 72681
rect 29825 72672 29837 72675
rect 29696 72644 29837 72672
rect 29696 72632 29702 72644
rect 29825 72641 29837 72644
rect 29871 72641 29883 72675
rect 29825 72635 29883 72641
rect 18230 72604 18236 72616
rect 15948 72576 18236 72604
rect 18230 72564 18236 72576
rect 18288 72564 18294 72616
rect 15013 72539 15071 72545
rect 15013 72505 15025 72539
rect 15059 72536 15071 72539
rect 17954 72536 17960 72548
rect 15059 72508 17960 72536
rect 15059 72505 15071 72508
rect 15013 72499 15071 72505
rect 17954 72496 17960 72508
rect 18012 72496 18018 72548
rect 1397 72471 1455 72477
rect 1397 72437 1409 72471
rect 1443 72468 1455 72471
rect 14826 72468 14832 72480
rect 1443 72440 14832 72468
rect 1443 72437 1455 72440
rect 1397 72431 1455 72437
rect 14826 72428 14832 72440
rect 14884 72428 14890 72480
rect 17218 72468 17224 72480
rect 17179 72440 17224 72468
rect 17218 72428 17224 72440
rect 17276 72428 17282 72480
rect 30006 72468 30012 72480
rect 29967 72440 30012 72468
rect 30006 72428 30012 72440
rect 30064 72428 30070 72480
rect 1104 72378 30820 72400
rect 1104 72326 5915 72378
rect 5967 72326 5979 72378
rect 6031 72326 6043 72378
rect 6095 72326 6107 72378
rect 6159 72326 6171 72378
rect 6223 72326 15846 72378
rect 15898 72326 15910 72378
rect 15962 72326 15974 72378
rect 16026 72326 16038 72378
rect 16090 72326 16102 72378
rect 16154 72326 25776 72378
rect 25828 72326 25840 72378
rect 25892 72326 25904 72378
rect 25956 72326 25968 72378
rect 26020 72326 26032 72378
rect 26084 72326 30820 72378
rect 1104 72304 30820 72326
rect 13357 72267 13415 72273
rect 13357 72233 13369 72267
rect 13403 72264 13415 72267
rect 14642 72264 14648 72276
rect 13403 72236 14648 72264
rect 13403 72233 13415 72236
rect 13357 72227 13415 72233
rect 14642 72224 14648 72236
rect 14700 72224 14706 72276
rect 18138 72264 18144 72276
rect 17144 72236 18144 72264
rect 1397 72199 1455 72205
rect 1397 72165 1409 72199
rect 1443 72196 1455 72199
rect 14734 72196 14740 72208
rect 1443 72168 14740 72196
rect 1443 72165 1455 72168
rect 1397 72159 1455 72165
rect 14734 72156 14740 72168
rect 14792 72156 14798 72208
rect 1578 72060 1584 72072
rect 1539 72032 1584 72060
rect 1578 72020 1584 72032
rect 1636 72020 1642 72072
rect 13538 72060 13544 72072
rect 13499 72032 13544 72060
rect 13538 72020 13544 72032
rect 13596 72020 13602 72072
rect 14642 72060 14648 72072
rect 14603 72032 14648 72060
rect 14642 72020 14648 72032
rect 14700 72020 14706 72072
rect 14826 72060 14832 72072
rect 14787 72032 14832 72060
rect 14826 72020 14832 72032
rect 14884 72020 14890 72072
rect 17144 72069 17172 72236
rect 18138 72224 18144 72236
rect 18196 72224 18202 72276
rect 17862 72128 17868 72140
rect 17236 72100 17868 72128
rect 17236 72069 17264 72100
rect 17862 72088 17868 72100
rect 17920 72088 17926 72140
rect 17129 72063 17187 72069
rect 17129 72029 17141 72063
rect 17175 72029 17187 72063
rect 17129 72023 17187 72029
rect 17221 72063 17279 72069
rect 17221 72029 17233 72063
rect 17267 72029 17279 72063
rect 17221 72023 17279 72029
rect 17310 72020 17316 72072
rect 17368 72060 17374 72072
rect 17497 72063 17555 72069
rect 17368 72032 17413 72060
rect 17368 72020 17374 72032
rect 17497 72029 17509 72063
rect 17543 72029 17555 72063
rect 17497 72023 17555 72029
rect 29825 72063 29883 72069
rect 29825 72029 29837 72063
rect 29871 72060 29883 72063
rect 30190 72060 30196 72072
rect 29871 72032 30196 72060
rect 29871 72029 29883 72032
rect 29825 72023 29883 72029
rect 15013 71995 15071 72001
rect 15013 71961 15025 71995
rect 15059 71992 15071 71995
rect 17512 71992 17540 72023
rect 30190 72020 30196 72032
rect 30248 72020 30254 72072
rect 15059 71964 17540 71992
rect 15059 71961 15071 71964
rect 15013 71955 15071 71961
rect 16853 71927 16911 71933
rect 16853 71893 16865 71927
rect 16899 71924 16911 71927
rect 16942 71924 16948 71936
rect 16899 71896 16948 71924
rect 16899 71893 16911 71896
rect 16853 71887 16911 71893
rect 16942 71884 16948 71896
rect 17000 71884 17006 71936
rect 30006 71924 30012 71936
rect 29967 71896 30012 71924
rect 30006 71884 30012 71896
rect 30064 71884 30070 71936
rect 1104 71834 30820 71856
rect 1104 71782 10880 71834
rect 10932 71782 10944 71834
rect 10996 71782 11008 71834
rect 11060 71782 11072 71834
rect 11124 71782 11136 71834
rect 11188 71782 20811 71834
rect 20863 71782 20875 71834
rect 20927 71782 20939 71834
rect 20991 71782 21003 71834
rect 21055 71782 21067 71834
rect 21119 71782 30820 71834
rect 1104 71760 30820 71782
rect 17310 71680 17316 71732
rect 17368 71720 17374 71732
rect 17368 71692 17908 71720
rect 17368 71680 17374 71692
rect 8294 71612 8300 71664
rect 8352 71652 8358 71664
rect 12989 71655 13047 71661
rect 12989 71652 13001 71655
rect 8352 71624 13001 71652
rect 8352 71612 8358 71624
rect 12989 71621 13001 71624
rect 13035 71621 13047 71655
rect 12989 71615 13047 71621
rect 12802 71584 12808 71596
rect 12763 71556 12808 71584
rect 12802 71544 12808 71556
rect 12860 71544 12866 71596
rect 17494 71544 17500 71596
rect 17552 71593 17558 71596
rect 17552 71587 17601 71593
rect 17552 71553 17555 71587
rect 17589 71553 17601 71587
rect 17552 71547 17601 71553
rect 17681 71587 17739 71593
rect 17681 71553 17693 71587
rect 17727 71553 17739 71587
rect 17681 71547 17739 71553
rect 17778 71587 17836 71593
rect 17778 71553 17790 71587
rect 17824 71584 17836 71587
rect 17880 71584 17908 71692
rect 20165 71655 20223 71661
rect 20165 71621 20177 71655
rect 20211 71652 20223 71655
rect 21266 71652 21272 71664
rect 20211 71624 21272 71652
rect 20211 71621 20223 71624
rect 20165 71615 20223 71621
rect 21266 71612 21272 71624
rect 21324 71612 21330 71664
rect 17824 71556 17908 71584
rect 17824 71553 17836 71556
rect 17778 71547 17836 71553
rect 17552 71544 17558 71547
rect 17696 71516 17724 71547
rect 17954 71544 17960 71596
rect 18012 71584 18018 71596
rect 20993 71587 21051 71593
rect 18012 71556 18057 71584
rect 18012 71544 18018 71556
rect 20993 71553 21005 71587
rect 21039 71584 21051 71587
rect 21450 71584 21456 71596
rect 21039 71556 21456 71584
rect 21039 71553 21051 71556
rect 20993 71547 21051 71553
rect 21450 71544 21456 71556
rect 21508 71544 21514 71596
rect 29825 71587 29883 71593
rect 29825 71553 29837 71587
rect 29871 71584 29883 71587
rect 30834 71584 30840 71596
rect 29871 71556 30840 71584
rect 29871 71553 29883 71556
rect 29825 71547 29883 71553
rect 30834 71544 30840 71556
rect 30892 71544 30898 71596
rect 17862 71516 17868 71528
rect 17696 71488 17868 71516
rect 17862 71476 17868 71488
rect 17920 71476 17926 71528
rect 18414 71476 18420 71528
rect 18472 71516 18478 71528
rect 19334 71516 19340 71528
rect 18472 71488 19340 71516
rect 18472 71476 18478 71488
rect 19334 71476 19340 71488
rect 19392 71476 19398 71528
rect 13173 71451 13231 71457
rect 13173 71417 13185 71451
rect 13219 71448 13231 71451
rect 22462 71448 22468 71460
rect 13219 71420 22468 71448
rect 13219 71417 13231 71420
rect 13173 71411 13231 71417
rect 22462 71408 22468 71420
rect 22520 71408 22526 71460
rect 17313 71383 17371 71389
rect 17313 71349 17325 71383
rect 17359 71380 17371 71383
rect 17954 71380 17960 71392
rect 17359 71352 17960 71380
rect 17359 71349 17371 71352
rect 17313 71343 17371 71349
rect 17954 71340 17960 71352
rect 18012 71340 18018 71392
rect 19794 71340 19800 71392
rect 19852 71380 19858 71392
rect 20257 71383 20315 71389
rect 20257 71380 20269 71383
rect 19852 71352 20269 71380
rect 19852 71340 19858 71352
rect 20257 71349 20269 71352
rect 20303 71349 20315 71383
rect 20257 71343 20315 71349
rect 21085 71383 21143 71389
rect 21085 71349 21097 71383
rect 21131 71380 21143 71383
rect 21358 71380 21364 71392
rect 21131 71352 21364 71380
rect 21131 71349 21143 71352
rect 21085 71343 21143 71349
rect 21358 71340 21364 71352
rect 21416 71340 21422 71392
rect 30006 71380 30012 71392
rect 29967 71352 30012 71380
rect 30006 71340 30012 71352
rect 30064 71340 30070 71392
rect 1104 71290 30820 71312
rect 1104 71238 5915 71290
rect 5967 71238 5979 71290
rect 6031 71238 6043 71290
rect 6095 71238 6107 71290
rect 6159 71238 6171 71290
rect 6223 71238 15846 71290
rect 15898 71238 15910 71290
rect 15962 71238 15974 71290
rect 16026 71238 16038 71290
rect 16090 71238 16102 71290
rect 16154 71238 25776 71290
rect 25828 71238 25840 71290
rect 25892 71238 25904 71290
rect 25956 71238 25968 71290
rect 26020 71238 26032 71290
rect 26084 71238 30820 71290
rect 1104 71216 30820 71238
rect 15013 71179 15071 71185
rect 15013 71145 15025 71179
rect 15059 71176 15071 71179
rect 16390 71176 16396 71188
rect 15059 71148 16396 71176
rect 15059 71145 15071 71148
rect 15013 71139 15071 71145
rect 16390 71136 16396 71148
rect 16448 71136 16454 71188
rect 18230 71176 18236 71188
rect 18191 71148 18236 71176
rect 18230 71136 18236 71148
rect 18288 71136 18294 71188
rect 20714 71136 20720 71188
rect 20772 71176 20778 71188
rect 20901 71179 20959 71185
rect 20901 71176 20913 71179
rect 20772 71148 20913 71176
rect 20772 71136 20778 71148
rect 20901 71145 20913 71148
rect 20947 71145 20959 71179
rect 20901 71139 20959 71145
rect 13173 71111 13231 71117
rect 13173 71077 13185 71111
rect 13219 71108 13231 71111
rect 19518 71108 19524 71120
rect 13219 71080 19524 71108
rect 13219 71077 13231 71080
rect 13173 71071 13231 71077
rect 19518 71068 19524 71080
rect 19576 71068 19582 71120
rect 1486 71000 1492 71052
rect 1544 71040 1550 71052
rect 16301 71043 16359 71049
rect 1544 71012 10916 71040
rect 1544 71000 1550 71012
rect 1394 70972 1400 70984
rect 1355 70944 1400 70972
rect 1394 70932 1400 70944
rect 1452 70932 1458 70984
rect 1673 70975 1731 70981
rect 1673 70941 1685 70975
rect 1719 70972 1731 70975
rect 9582 70972 9588 70984
rect 1719 70944 9588 70972
rect 1719 70941 1731 70944
rect 1673 70935 1731 70941
rect 9582 70932 9588 70944
rect 9640 70932 9646 70984
rect 10888 70836 10916 71012
rect 16301 71009 16313 71043
rect 16347 71040 16359 71043
rect 16482 71040 16488 71052
rect 16347 71012 16488 71040
rect 16347 71009 16359 71012
rect 16301 71003 16359 71009
rect 16482 71000 16488 71012
rect 16540 71000 16546 71052
rect 11790 70932 11796 70984
rect 11848 70972 11854 70984
rect 12989 70975 13047 70981
rect 12989 70972 13001 70975
rect 11848 70944 13001 70972
rect 11848 70932 11854 70944
rect 12989 70941 13001 70944
rect 13035 70941 13047 70975
rect 14829 70975 14887 70981
rect 14829 70972 14841 70975
rect 12989 70935 13047 70941
rect 13096 70944 14841 70972
rect 12802 70904 12808 70916
rect 12763 70876 12808 70904
rect 12802 70864 12808 70876
rect 12860 70864 12866 70916
rect 13096 70836 13124 70944
rect 14829 70941 14841 70944
rect 14875 70941 14887 70975
rect 14829 70935 14887 70941
rect 16574 70932 16580 70984
rect 16632 70972 16638 70984
rect 17402 70972 17408 70984
rect 16632 70944 17408 70972
rect 16632 70932 16638 70944
rect 17402 70932 17408 70944
rect 17460 70932 17466 70984
rect 29825 70975 29883 70981
rect 29825 70941 29837 70975
rect 29871 70972 29883 70975
rect 30282 70972 30288 70984
rect 29871 70944 30288 70972
rect 29871 70941 29883 70944
rect 29825 70935 29883 70941
rect 30282 70932 30288 70944
rect 30340 70932 30346 70984
rect 14642 70904 14648 70916
rect 14603 70876 14648 70904
rect 14642 70864 14648 70876
rect 14700 70864 14706 70916
rect 16393 70907 16451 70913
rect 16393 70873 16405 70907
rect 16439 70904 16451 70907
rect 16592 70904 16620 70932
rect 16439 70876 16620 70904
rect 16945 70907 17003 70913
rect 16439 70873 16451 70876
rect 16393 70867 16451 70873
rect 16945 70873 16957 70907
rect 16991 70904 17003 70907
rect 18414 70904 18420 70916
rect 16991 70876 18420 70904
rect 16991 70873 17003 70876
rect 16945 70867 17003 70873
rect 18414 70864 18420 70876
rect 18472 70864 18478 70916
rect 19610 70904 19616 70916
rect 19571 70876 19616 70904
rect 19610 70864 19616 70876
rect 19668 70864 19674 70916
rect 10888 70808 13124 70836
rect 15562 70796 15568 70848
rect 15620 70836 15626 70848
rect 15823 70839 15881 70845
rect 15823 70836 15835 70839
rect 15620 70808 15835 70836
rect 15620 70796 15626 70808
rect 15823 70805 15835 70808
rect 15869 70805 15881 70839
rect 15823 70799 15881 70805
rect 16301 70839 16359 70845
rect 16301 70805 16313 70839
rect 16347 70836 16359 70839
rect 17218 70836 17224 70848
rect 16347 70808 17224 70836
rect 16347 70805 16359 70808
rect 16301 70799 16359 70805
rect 17218 70796 17224 70808
rect 17276 70796 17282 70848
rect 30006 70836 30012 70848
rect 29967 70808 30012 70836
rect 30006 70796 30012 70808
rect 30064 70796 30070 70848
rect 1104 70746 30820 70768
rect 1104 70694 10880 70746
rect 10932 70694 10944 70746
rect 10996 70694 11008 70746
rect 11060 70694 11072 70746
rect 11124 70694 11136 70746
rect 11188 70694 20811 70746
rect 20863 70694 20875 70746
rect 20927 70694 20939 70746
rect 20991 70694 21003 70746
rect 21055 70694 21067 70746
rect 21119 70694 30820 70746
rect 1104 70672 30820 70694
rect 1397 70635 1455 70641
rect 1397 70601 1409 70635
rect 1443 70632 1455 70635
rect 1486 70632 1492 70644
rect 1443 70604 1492 70632
rect 1443 70601 1455 70604
rect 1397 70595 1455 70601
rect 1486 70592 1492 70604
rect 1544 70592 1550 70644
rect 12161 70635 12219 70641
rect 12161 70601 12173 70635
rect 12207 70632 12219 70635
rect 12802 70632 12808 70644
rect 12207 70604 12808 70632
rect 12207 70601 12219 70604
rect 12161 70595 12219 70601
rect 12802 70592 12808 70604
rect 12860 70592 12866 70644
rect 15105 70635 15163 70641
rect 15105 70601 15117 70635
rect 15151 70632 15163 70635
rect 15151 70604 16896 70632
rect 15151 70601 15163 70604
rect 15105 70595 15163 70601
rect 11698 70524 11704 70576
rect 11756 70564 11762 70576
rect 12989 70567 13047 70573
rect 12989 70564 13001 70567
rect 11756 70536 13001 70564
rect 11756 70524 11762 70536
rect 12989 70533 13001 70536
rect 13035 70533 13047 70567
rect 12989 70527 13047 70533
rect 13173 70567 13231 70573
rect 13173 70533 13185 70567
rect 13219 70564 13231 70567
rect 15470 70564 15476 70576
rect 13219 70536 15476 70564
rect 13219 70533 13231 70536
rect 13173 70527 13231 70533
rect 15470 70524 15476 70536
rect 15528 70524 15534 70576
rect 1578 70496 1584 70508
rect 1539 70468 1584 70496
rect 1578 70456 1584 70468
rect 1636 70456 1642 70508
rect 12345 70499 12403 70505
rect 12345 70465 12357 70499
rect 12391 70465 12403 70499
rect 12802 70496 12808 70508
rect 12715 70468 12808 70496
rect 12345 70459 12403 70465
rect 12360 70428 12388 70459
rect 12802 70456 12808 70468
rect 12860 70496 12866 70508
rect 13633 70499 13691 70505
rect 13633 70496 13645 70499
rect 12860 70468 13645 70496
rect 12860 70456 12866 70468
rect 13633 70465 13645 70468
rect 13679 70465 13691 70499
rect 13633 70459 13691 70465
rect 13722 70456 13728 70508
rect 13780 70496 13786 70508
rect 13817 70499 13875 70505
rect 13817 70496 13829 70499
rect 13780 70468 13829 70496
rect 13780 70456 13786 70468
rect 13817 70465 13829 70468
rect 13863 70465 13875 70499
rect 13817 70459 13875 70465
rect 14921 70499 14979 70505
rect 14921 70465 14933 70499
rect 14967 70465 14979 70499
rect 15562 70496 15568 70508
rect 15523 70468 15568 70496
rect 14921 70459 14979 70465
rect 13538 70428 13544 70440
rect 12360 70400 13544 70428
rect 13538 70388 13544 70400
rect 13596 70388 13602 70440
rect 14001 70431 14059 70437
rect 14001 70397 14013 70431
rect 14047 70428 14059 70431
rect 14826 70428 14832 70440
rect 14047 70400 14832 70428
rect 14047 70397 14059 70400
rect 14001 70391 14059 70397
rect 14826 70388 14832 70400
rect 14884 70388 14890 70440
rect 14936 70428 14964 70459
rect 15562 70456 15568 70468
rect 15620 70456 15626 70508
rect 16868 70505 16896 70604
rect 18138 70592 18144 70644
rect 18196 70632 18202 70644
rect 18233 70635 18291 70641
rect 18233 70632 18245 70635
rect 18196 70604 18245 70632
rect 18196 70592 18202 70604
rect 18233 70601 18245 70604
rect 18279 70632 18291 70635
rect 18322 70632 18328 70644
rect 18279 70604 18328 70632
rect 18279 70601 18291 70604
rect 18233 70595 18291 70601
rect 18322 70592 18328 70604
rect 18380 70592 18386 70644
rect 19702 70592 19708 70644
rect 19760 70632 19766 70644
rect 19978 70632 19984 70644
rect 19760 70604 19984 70632
rect 19760 70592 19766 70604
rect 19978 70592 19984 70604
rect 20036 70592 20042 70644
rect 22370 70524 22376 70576
rect 22428 70564 22434 70576
rect 22428 70536 22508 70564
rect 22428 70524 22434 70536
rect 16853 70499 16911 70505
rect 16853 70465 16865 70499
rect 16899 70465 16911 70499
rect 16853 70459 16911 70465
rect 16942 70456 16948 70508
rect 17000 70496 17006 70508
rect 17109 70499 17167 70505
rect 17109 70496 17121 70499
rect 17000 70468 17121 70496
rect 17000 70456 17006 70468
rect 17109 70465 17121 70468
rect 17155 70465 17167 70499
rect 17109 70459 17167 70465
rect 18693 70499 18751 70505
rect 18693 70465 18705 70499
rect 18739 70496 18751 70499
rect 19426 70496 19432 70508
rect 18739 70468 19432 70496
rect 18739 70465 18751 70468
rect 18693 70459 18751 70465
rect 19426 70456 19432 70468
rect 19484 70456 19490 70508
rect 19518 70456 19524 70508
rect 19576 70496 19582 70508
rect 19702 70496 19708 70508
rect 19576 70468 19708 70496
rect 19576 70456 19582 70468
rect 19702 70456 19708 70468
rect 19760 70456 19766 70508
rect 20806 70456 20812 70508
rect 20864 70496 20870 70508
rect 20901 70499 20959 70505
rect 20901 70496 20913 70499
rect 20864 70468 20913 70496
rect 20864 70456 20870 70468
rect 20901 70465 20913 70468
rect 20947 70465 20959 70499
rect 20901 70459 20959 70465
rect 22002 70456 22008 70508
rect 22060 70505 22066 70508
rect 22060 70499 22109 70505
rect 22186 70502 22244 70508
rect 22186 70499 22198 70502
rect 22060 70465 22063 70499
rect 22097 70465 22109 70499
rect 22060 70459 22109 70465
rect 22185 70468 22198 70499
rect 22232 70468 22244 70502
rect 22185 70462 22244 70468
rect 22060 70456 22066 70459
rect 16758 70428 16764 70440
rect 14936 70400 16764 70428
rect 16758 70388 16764 70400
rect 16816 70388 16822 70440
rect 21358 70388 21364 70440
rect 21416 70428 21422 70440
rect 22185 70428 22213 70462
rect 22278 70456 22284 70508
rect 22336 70505 22342 70508
rect 22480 70505 22508 70536
rect 22336 70496 22344 70505
rect 22465 70499 22523 70505
rect 22336 70468 22381 70496
rect 22336 70459 22344 70468
rect 22465 70465 22477 70499
rect 22511 70465 22523 70499
rect 22465 70459 22523 70465
rect 22336 70456 22342 70459
rect 29178 70456 29184 70508
rect 29236 70496 29242 70508
rect 29825 70499 29883 70505
rect 29825 70496 29837 70499
rect 29236 70468 29837 70496
rect 29236 70456 29242 70468
rect 29825 70465 29837 70468
rect 29871 70465 29883 70499
rect 29825 70459 29883 70465
rect 21416 70400 22213 70428
rect 21416 70388 21422 70400
rect 15746 70292 15752 70304
rect 15707 70264 15752 70292
rect 15746 70252 15752 70264
rect 15804 70252 15810 70304
rect 21082 70292 21088 70304
rect 21043 70264 21088 70292
rect 21082 70252 21088 70264
rect 21140 70252 21146 70304
rect 21818 70292 21824 70304
rect 21779 70264 21824 70292
rect 21818 70252 21824 70264
rect 21876 70252 21882 70304
rect 30006 70292 30012 70304
rect 29967 70264 30012 70292
rect 30006 70252 30012 70264
rect 30064 70252 30070 70304
rect 1104 70202 30820 70224
rect 1104 70150 5915 70202
rect 5967 70150 5979 70202
rect 6031 70150 6043 70202
rect 6095 70150 6107 70202
rect 6159 70150 6171 70202
rect 6223 70150 15846 70202
rect 15898 70150 15910 70202
rect 15962 70150 15974 70202
rect 16026 70150 16038 70202
rect 16090 70150 16102 70202
rect 16154 70150 25776 70202
rect 25828 70150 25840 70202
rect 25892 70150 25904 70202
rect 25956 70150 25968 70202
rect 26020 70150 26032 70202
rect 26084 70150 30820 70202
rect 1104 70128 30820 70150
rect 13173 70091 13231 70097
rect 13173 70057 13185 70091
rect 13219 70088 13231 70091
rect 18506 70088 18512 70100
rect 13219 70060 18512 70088
rect 13219 70057 13231 70060
rect 13173 70051 13231 70057
rect 18506 70048 18512 70060
rect 18564 70048 18570 70100
rect 19337 70091 19395 70097
rect 19337 70057 19349 70091
rect 19383 70088 19395 70091
rect 20806 70088 20812 70100
rect 19383 70060 20812 70088
rect 19383 70057 19395 70060
rect 19337 70051 19395 70057
rect 20806 70048 20812 70060
rect 20864 70048 20870 70100
rect 21821 70091 21879 70097
rect 21821 70057 21833 70091
rect 21867 70088 21879 70091
rect 22002 70088 22008 70100
rect 21867 70060 22008 70088
rect 21867 70057 21879 70060
rect 21821 70051 21879 70057
rect 22002 70048 22008 70060
rect 22060 70088 22066 70100
rect 24210 70088 24216 70100
rect 22060 70060 24216 70088
rect 22060 70048 22066 70060
rect 24210 70048 24216 70060
rect 24268 70048 24274 70100
rect 29086 69980 29092 70032
rect 29144 69980 29150 70032
rect 1578 69884 1584 69896
rect 1539 69856 1584 69884
rect 1578 69844 1584 69856
rect 1636 69844 1642 69896
rect 10778 69844 10784 69896
rect 10836 69884 10842 69896
rect 12802 69884 12808 69896
rect 10836 69856 12434 69884
rect 12763 69856 12808 69884
rect 10836 69844 10842 69856
rect 12406 69816 12434 69856
rect 12802 69844 12808 69856
rect 12860 69844 12866 69896
rect 14737 69887 14795 69893
rect 14737 69853 14749 69887
rect 14783 69884 14795 69887
rect 15746 69884 15752 69896
rect 14783 69856 15752 69884
rect 14783 69853 14795 69856
rect 14737 69847 14795 69853
rect 15746 69844 15752 69856
rect 15804 69844 15810 69896
rect 20441 69887 20499 69893
rect 20441 69853 20453 69887
rect 20487 69884 20499 69887
rect 21082 69884 21088 69896
rect 20487 69856 21088 69884
rect 20487 69853 20499 69856
rect 20441 69847 20499 69853
rect 21082 69844 21088 69856
rect 21140 69844 21146 69896
rect 22278 69884 22284 69896
rect 22239 69856 22284 69884
rect 22278 69844 22284 69856
rect 22336 69844 22342 69896
rect 12989 69819 13047 69825
rect 12989 69816 13001 69819
rect 12406 69788 13001 69816
rect 12989 69785 13001 69788
rect 13035 69785 13047 69819
rect 12989 69779 13047 69785
rect 14642 69776 14648 69828
rect 14700 69816 14706 69828
rect 14982 69819 15040 69825
rect 14982 69816 14994 69819
rect 14700 69788 14994 69816
rect 14700 69776 14706 69788
rect 14982 69785 14994 69788
rect 15028 69785 15040 69819
rect 14982 69779 15040 69785
rect 16669 69819 16727 69825
rect 16669 69785 16681 69819
rect 16715 69816 16727 69819
rect 18046 69816 18052 69828
rect 16715 69788 18052 69816
rect 16715 69785 16727 69788
rect 16669 69779 16727 69785
rect 18046 69776 18052 69788
rect 18104 69776 18110 69828
rect 19518 69776 19524 69828
rect 19576 69816 19582 69828
rect 19613 69819 19671 69825
rect 19613 69816 19625 69819
rect 19576 69788 19625 69816
rect 19576 69776 19582 69788
rect 19613 69785 19625 69788
rect 19659 69785 19671 69819
rect 19794 69816 19800 69828
rect 19755 69788 19800 69816
rect 19613 69779 19671 69785
rect 19794 69776 19800 69788
rect 19852 69776 19858 69828
rect 19886 69776 19892 69828
rect 19944 69816 19950 69828
rect 20708 69819 20766 69825
rect 19944 69788 19989 69816
rect 19944 69776 19950 69788
rect 20708 69785 20720 69819
rect 20754 69816 20766 69819
rect 21818 69816 21824 69828
rect 20754 69788 21824 69816
rect 20754 69785 20766 69788
rect 20708 69779 20766 69785
rect 21818 69776 21824 69788
rect 21876 69776 21882 69828
rect 21910 69776 21916 69828
rect 21968 69816 21974 69828
rect 22526 69819 22584 69825
rect 22526 69816 22538 69819
rect 21968 69788 22538 69816
rect 21968 69776 21974 69788
rect 22526 69785 22538 69788
rect 22572 69785 22584 69819
rect 22526 69779 22584 69785
rect 1397 69751 1455 69757
rect 1397 69717 1409 69751
rect 1443 69748 1455 69751
rect 9950 69748 9956 69760
rect 1443 69720 9956 69748
rect 1443 69717 1455 69720
rect 1397 69711 1455 69717
rect 9950 69708 9956 69720
rect 10008 69708 10014 69760
rect 16117 69751 16175 69757
rect 16117 69717 16129 69751
rect 16163 69748 16175 69751
rect 16206 69748 16212 69760
rect 16163 69720 16212 69748
rect 16163 69717 16175 69720
rect 16117 69711 16175 69717
rect 16206 69708 16212 69720
rect 16264 69708 16270 69760
rect 17126 69708 17132 69760
rect 17184 69748 17190 69760
rect 17402 69748 17408 69760
rect 17184 69720 17408 69748
rect 17184 69708 17190 69720
rect 17402 69708 17408 69720
rect 17460 69748 17466 69760
rect 17957 69751 18015 69757
rect 17957 69748 17969 69751
rect 17460 69720 17969 69748
rect 17460 69708 17466 69720
rect 17957 69717 17969 69720
rect 18003 69717 18015 69751
rect 17957 69711 18015 69717
rect 22094 69708 22100 69760
rect 22152 69748 22158 69760
rect 23661 69751 23719 69757
rect 23661 69748 23673 69751
rect 22152 69720 23673 69748
rect 22152 69708 22158 69720
rect 23661 69717 23673 69720
rect 23707 69748 23719 69751
rect 25498 69748 25504 69760
rect 23707 69720 25504 69748
rect 23707 69717 23719 69720
rect 23661 69711 23719 69717
rect 25498 69708 25504 69720
rect 25556 69708 25562 69760
rect 28994 69708 29000 69760
rect 29052 69748 29058 69760
rect 29104 69748 29132 69980
rect 29825 69887 29883 69893
rect 29825 69853 29837 69887
rect 29871 69884 29883 69887
rect 30650 69884 30656 69896
rect 29871 69856 30656 69884
rect 29871 69853 29883 69856
rect 29825 69847 29883 69853
rect 30650 69844 30656 69856
rect 30708 69844 30714 69896
rect 30006 69748 30012 69760
rect 29052 69720 29132 69748
rect 29967 69720 30012 69748
rect 29052 69708 29058 69720
rect 30006 69708 30012 69720
rect 30064 69708 30070 69760
rect 1104 69658 30820 69680
rect 1104 69606 10880 69658
rect 10932 69606 10944 69658
rect 10996 69606 11008 69658
rect 11060 69606 11072 69658
rect 11124 69606 11136 69658
rect 11188 69606 20811 69658
rect 20863 69606 20875 69658
rect 20927 69606 20939 69658
rect 20991 69606 21003 69658
rect 21055 69606 21067 69658
rect 21119 69606 30820 69658
rect 1104 69584 30820 69606
rect 21821 69547 21879 69553
rect 21821 69513 21833 69547
rect 21867 69544 21879 69547
rect 21910 69544 21916 69556
rect 21867 69516 21916 69544
rect 21867 69513 21879 69516
rect 21821 69507 21879 69513
rect 21910 69504 21916 69516
rect 21968 69504 21974 69556
rect 29178 69504 29184 69556
rect 29236 69544 29242 69556
rect 29822 69544 29828 69556
rect 29236 69516 29828 69544
rect 29236 69504 29242 69516
rect 29822 69504 29828 69516
rect 29880 69504 29886 69556
rect 9950 69436 9956 69488
rect 10008 69476 10014 69488
rect 12989 69479 13047 69485
rect 12989 69476 13001 69479
rect 10008 69448 13001 69476
rect 10008 69436 10014 69448
rect 12989 69445 13001 69448
rect 13035 69445 13047 69479
rect 12989 69439 13047 69445
rect 17954 69436 17960 69488
rect 18012 69476 18018 69488
rect 18386 69479 18444 69485
rect 18386 69476 18398 69479
rect 18012 69448 18398 69476
rect 18012 69436 18018 69448
rect 18386 69445 18398 69448
rect 18432 69445 18444 69479
rect 18386 69439 18444 69445
rect 20257 69479 20315 69485
rect 20257 69445 20269 69479
rect 20303 69476 20315 69479
rect 20622 69476 20628 69488
rect 20303 69448 20628 69476
rect 20303 69445 20315 69448
rect 20257 69439 20315 69445
rect 20622 69436 20628 69448
rect 20680 69476 20686 69488
rect 22370 69476 22376 69488
rect 20680 69448 22376 69476
rect 20680 69436 20686 69448
rect 1578 69408 1584 69420
rect 1539 69380 1584 69408
rect 1578 69368 1584 69380
rect 1636 69368 1642 69420
rect 12618 69368 12624 69420
rect 12676 69408 12682 69420
rect 12805 69411 12863 69417
rect 12805 69408 12817 69411
rect 12676 69380 12817 69408
rect 12676 69368 12682 69380
rect 12805 69377 12817 69380
rect 12851 69377 12863 69411
rect 12805 69371 12863 69377
rect 13998 69368 14004 69420
rect 14056 69408 14062 69420
rect 14165 69411 14223 69417
rect 14165 69408 14177 69411
rect 14056 69380 14177 69408
rect 14056 69368 14062 69380
rect 14165 69377 14177 69380
rect 14211 69377 14223 69411
rect 14165 69371 14223 69377
rect 17129 69411 17187 69417
rect 17129 69377 17141 69411
rect 17175 69408 17187 69411
rect 17310 69408 17316 69420
rect 17175 69380 17316 69408
rect 17175 69377 17187 69380
rect 17129 69371 17187 69377
rect 17310 69368 17316 69380
rect 17368 69368 17374 69420
rect 20073 69411 20131 69417
rect 20073 69408 20085 69411
rect 17972 69380 20085 69408
rect 13906 69340 13912 69352
rect 13867 69312 13912 69340
rect 13906 69300 13912 69312
rect 13964 69300 13970 69352
rect 16666 69300 16672 69352
rect 16724 69340 16730 69352
rect 16853 69343 16911 69349
rect 16853 69340 16865 69343
rect 16724 69312 16865 69340
rect 16724 69300 16730 69312
rect 16853 69309 16865 69312
rect 16899 69340 16911 69343
rect 17972 69340 18000 69380
rect 20073 69377 20085 69380
rect 20119 69408 20131 69411
rect 20438 69408 20444 69420
rect 20119 69380 20444 69408
rect 20119 69377 20131 69380
rect 20073 69371 20131 69377
rect 20438 69368 20444 69380
rect 20496 69368 20502 69420
rect 21085 69411 21143 69417
rect 21085 69377 21097 69411
rect 21131 69408 21143 69411
rect 21450 69408 21456 69420
rect 21131 69380 21456 69408
rect 21131 69377 21143 69380
rect 21085 69371 21143 69377
rect 21450 69368 21456 69380
rect 21508 69368 21514 69420
rect 22094 69408 22100 69420
rect 22055 69380 22100 69408
rect 22094 69368 22100 69380
rect 22152 69368 22158 69420
rect 22296 69417 22324 69448
rect 22370 69436 22376 69448
rect 22428 69436 22434 69488
rect 29546 69436 29552 69488
rect 29604 69476 29610 69488
rect 29730 69476 29736 69488
rect 29604 69448 29736 69476
rect 29604 69436 29610 69448
rect 29730 69436 29736 69448
rect 29788 69436 29794 69488
rect 22189 69411 22247 69417
rect 22189 69377 22201 69411
rect 22235 69377 22247 69411
rect 22189 69371 22247 69377
rect 22281 69411 22339 69417
rect 22281 69377 22293 69411
rect 22327 69377 22339 69411
rect 22462 69408 22468 69420
rect 22423 69380 22468 69408
rect 22281 69371 22339 69377
rect 18138 69340 18144 69352
rect 16899 69312 18000 69340
rect 18099 69312 18144 69340
rect 16899 69309 16911 69312
rect 16853 69303 16911 69309
rect 18138 69300 18144 69312
rect 18196 69300 18202 69352
rect 19702 69300 19708 69352
rect 19760 69340 19766 69352
rect 20254 69340 20260 69352
rect 19760 69312 20260 69340
rect 19760 69300 19766 69312
rect 20254 69300 20260 69312
rect 20312 69300 20318 69352
rect 22204 69284 22232 69371
rect 22462 69368 22468 69380
rect 22520 69368 22526 69420
rect 28442 69368 28448 69420
rect 28500 69408 28506 69420
rect 29089 69411 29147 69417
rect 29089 69408 29101 69411
rect 28500 69380 29101 69408
rect 28500 69368 28506 69380
rect 29089 69377 29101 69380
rect 29135 69377 29147 69411
rect 29825 69411 29883 69417
rect 29825 69408 29837 69411
rect 29089 69371 29147 69377
rect 29380 69380 29837 69408
rect 29380 69352 29408 69380
rect 29825 69377 29837 69380
rect 29871 69377 29883 69411
rect 29825 69371 29883 69377
rect 29362 69300 29368 69352
rect 29420 69300 29426 69352
rect 21269 69275 21327 69281
rect 21269 69241 21281 69275
rect 21315 69272 21327 69275
rect 22186 69272 22192 69284
rect 21315 69244 22192 69272
rect 21315 69241 21327 69244
rect 21269 69235 21327 69241
rect 22186 69232 22192 69244
rect 22244 69232 22250 69284
rect 29270 69272 29276 69284
rect 29231 69244 29276 69272
rect 29270 69232 29276 69244
rect 29328 69232 29334 69284
rect 1397 69207 1455 69213
rect 1397 69173 1409 69207
rect 1443 69204 1455 69207
rect 11330 69204 11336 69216
rect 1443 69176 11336 69204
rect 1443 69173 1455 69176
rect 1397 69167 1455 69173
rect 11330 69164 11336 69176
rect 11388 69164 11394 69216
rect 13173 69207 13231 69213
rect 13173 69173 13185 69207
rect 13219 69204 13231 69207
rect 14826 69204 14832 69216
rect 13219 69176 14832 69204
rect 13219 69173 13231 69176
rect 13173 69167 13231 69173
rect 14826 69164 14832 69176
rect 14884 69164 14890 69216
rect 15289 69207 15347 69213
rect 15289 69173 15301 69207
rect 15335 69204 15347 69207
rect 16298 69204 16304 69216
rect 15335 69176 16304 69204
rect 15335 69173 15347 69176
rect 15289 69167 15347 69173
rect 16298 69164 16304 69176
rect 16356 69164 16362 69216
rect 19334 69164 19340 69216
rect 19392 69204 19398 69216
rect 19521 69207 19579 69213
rect 19521 69204 19533 69207
rect 19392 69176 19533 69204
rect 19392 69164 19398 69176
rect 19521 69173 19533 69176
rect 19567 69204 19579 69207
rect 19702 69204 19708 69216
rect 19567 69176 19708 69204
rect 19567 69173 19579 69176
rect 19521 69167 19579 69173
rect 19702 69164 19708 69176
rect 19760 69164 19766 69216
rect 29914 69164 29920 69216
rect 29972 69204 29978 69216
rect 30009 69207 30067 69213
rect 30009 69204 30021 69207
rect 29972 69176 30021 69204
rect 29972 69164 29978 69176
rect 30009 69173 30021 69176
rect 30055 69173 30067 69207
rect 30009 69167 30067 69173
rect 1104 69114 30820 69136
rect 1104 69062 5915 69114
rect 5967 69062 5979 69114
rect 6031 69062 6043 69114
rect 6095 69062 6107 69114
rect 6159 69062 6171 69114
rect 6223 69062 15846 69114
rect 15898 69062 15910 69114
rect 15962 69062 15974 69114
rect 16026 69062 16038 69114
rect 16090 69062 16102 69114
rect 16154 69062 25776 69114
rect 25828 69062 25840 69114
rect 25892 69062 25904 69114
rect 25956 69062 25968 69114
rect 26020 69062 26032 69114
rect 26084 69062 30820 69114
rect 1104 69040 30820 69062
rect 14642 69000 14648 69012
rect 14603 68972 14648 69000
rect 14642 68960 14648 68972
rect 14700 68960 14706 69012
rect 16758 68960 16764 69012
rect 16816 69000 16822 69012
rect 17037 69003 17095 69009
rect 17037 69000 17049 69003
rect 16816 68972 17049 69000
rect 16816 68960 16822 68972
rect 17037 68969 17049 68972
rect 17083 68969 17095 69003
rect 17037 68963 17095 68969
rect 19981 69003 20039 69009
rect 19981 68969 19993 69003
rect 20027 69000 20039 69003
rect 20530 69000 20536 69012
rect 20027 68972 20536 69000
rect 20027 68969 20039 68972
rect 19981 68963 20039 68969
rect 20530 68960 20536 68972
rect 20588 68960 20594 69012
rect 22005 69003 22063 69009
rect 22005 68969 22017 69003
rect 22051 69000 22063 69003
rect 22278 69000 22284 69012
rect 22051 68972 22284 69000
rect 22051 68969 22063 68972
rect 22005 68963 22063 68969
rect 22278 68960 22284 68972
rect 22336 68960 22342 69012
rect 16206 68932 16212 68944
rect 14752 68904 16212 68932
rect 1578 68796 1584 68808
rect 1539 68768 1584 68796
rect 1578 68756 1584 68768
rect 1636 68756 1642 68808
rect 12618 68796 12624 68808
rect 12579 68768 12624 68796
rect 12618 68756 12624 68768
rect 12676 68756 12682 68808
rect 14752 68796 14780 68904
rect 16206 68892 16212 68904
rect 16264 68932 16270 68944
rect 24762 68932 24768 68944
rect 16264 68904 24768 68932
rect 16264 68892 16270 68904
rect 24762 68892 24768 68904
rect 24820 68892 24826 68944
rect 14826 68824 14832 68876
rect 14884 68864 14890 68876
rect 14884 68836 15332 68864
rect 14884 68824 14890 68836
rect 14921 68799 14979 68805
rect 14921 68796 14933 68799
rect 14752 68768 14933 68796
rect 14921 68765 14933 68768
rect 14967 68765 14979 68799
rect 14921 68759 14979 68765
rect 15013 68799 15071 68805
rect 15013 68765 15025 68799
rect 15059 68765 15071 68799
rect 15013 68759 15071 68765
rect 15105 68799 15163 68805
rect 15105 68765 15117 68799
rect 15151 68796 15163 68799
rect 15194 68796 15200 68808
rect 15151 68768 15200 68796
rect 15151 68765 15163 68768
rect 15105 68759 15163 68765
rect 12802 68728 12808 68740
rect 12763 68700 12808 68728
rect 12802 68688 12808 68700
rect 12860 68688 12866 68740
rect 14182 68688 14188 68740
rect 14240 68728 14246 68740
rect 15028 68728 15056 68759
rect 15194 68756 15200 68768
rect 15252 68756 15258 68808
rect 15304 68805 15332 68836
rect 17494 68824 17500 68876
rect 17552 68864 17558 68876
rect 17589 68867 17647 68873
rect 17589 68864 17601 68867
rect 17552 68836 17601 68864
rect 17552 68824 17558 68836
rect 17589 68833 17601 68836
rect 17635 68833 17647 68867
rect 17589 68827 17647 68833
rect 20346 68824 20352 68876
rect 20404 68864 20410 68876
rect 20441 68867 20499 68873
rect 20441 68864 20453 68867
rect 20404 68836 20453 68864
rect 20404 68824 20410 68836
rect 20441 68833 20453 68836
rect 20487 68864 20499 68867
rect 21361 68867 21419 68873
rect 21361 68864 21373 68867
rect 20487 68836 21373 68864
rect 20487 68833 20499 68836
rect 20441 68827 20499 68833
rect 21361 68833 21373 68836
rect 21407 68833 21419 68867
rect 21361 68827 21419 68833
rect 15289 68799 15347 68805
rect 15289 68765 15301 68799
rect 15335 68765 15347 68799
rect 15289 68759 15347 68765
rect 18417 68799 18475 68805
rect 18417 68765 18429 68799
rect 18463 68796 18475 68799
rect 19978 68796 19984 68808
rect 18463 68768 19984 68796
rect 18463 68765 18475 68768
rect 18417 68759 18475 68765
rect 19978 68756 19984 68768
rect 20036 68756 20042 68808
rect 20070 68756 20076 68808
rect 20128 68796 20134 68808
rect 21821 68799 21879 68805
rect 21821 68796 21833 68799
rect 20128 68768 21833 68796
rect 20128 68756 20134 68768
rect 21821 68765 21833 68768
rect 21867 68765 21879 68799
rect 21821 68759 21879 68765
rect 27246 68756 27252 68808
rect 27304 68796 27310 68808
rect 28721 68799 28779 68805
rect 28721 68796 28733 68799
rect 27304 68768 28733 68796
rect 27304 68756 27310 68768
rect 28721 68765 28733 68768
rect 28767 68765 28779 68799
rect 28721 68759 28779 68765
rect 29270 68756 29276 68808
rect 29328 68796 29334 68808
rect 29825 68799 29883 68805
rect 29825 68796 29837 68799
rect 29328 68768 29837 68796
rect 29328 68756 29334 68768
rect 29825 68765 29837 68768
rect 29871 68765 29883 68799
rect 29825 68759 29883 68765
rect 17310 68728 17316 68740
rect 14240 68700 15056 68728
rect 17271 68700 17316 68728
rect 14240 68688 14246 68700
rect 17310 68688 17316 68700
rect 17368 68688 17374 68740
rect 18598 68728 18604 68740
rect 18559 68700 18604 68728
rect 18598 68688 18604 68700
rect 18656 68688 18662 68740
rect 19794 68688 19800 68740
rect 19852 68728 19858 68740
rect 20438 68728 20444 68740
rect 19852 68700 20444 68728
rect 19852 68688 19858 68700
rect 20438 68688 20444 68700
rect 20496 68688 20502 68740
rect 20530 68688 20536 68740
rect 20588 68728 20594 68740
rect 21177 68731 21235 68737
rect 20588 68700 20633 68728
rect 20588 68688 20594 68700
rect 21177 68697 21189 68731
rect 21223 68697 21235 68731
rect 21177 68691 21235 68697
rect 1394 68660 1400 68672
rect 1355 68632 1400 68660
rect 1394 68620 1400 68632
rect 1452 68620 1458 68672
rect 12989 68663 13047 68669
rect 12989 68629 13001 68663
rect 13035 68660 13047 68663
rect 14458 68660 14464 68672
rect 13035 68632 14464 68660
rect 13035 68629 13047 68632
rect 12989 68623 13047 68629
rect 14458 68620 14464 68632
rect 14516 68620 14522 68672
rect 17497 68663 17555 68669
rect 17497 68629 17509 68663
rect 17543 68660 17555 68663
rect 18616 68660 18644 68688
rect 17543 68632 18644 68660
rect 17543 68629 17555 68632
rect 17497 68623 17555 68629
rect 20622 68620 20628 68672
rect 20680 68660 20686 68672
rect 21192 68660 21220 68691
rect 28902 68660 28908 68672
rect 20680 68632 21220 68660
rect 28863 68632 28908 68660
rect 20680 68620 20686 68632
rect 28902 68620 28908 68632
rect 28960 68620 28966 68672
rect 30006 68660 30012 68672
rect 29967 68632 30012 68660
rect 30006 68620 30012 68632
rect 30064 68620 30070 68672
rect 1104 68570 30820 68592
rect 1104 68518 10880 68570
rect 10932 68518 10944 68570
rect 10996 68518 11008 68570
rect 11060 68518 11072 68570
rect 11124 68518 11136 68570
rect 11188 68518 20811 68570
rect 20863 68518 20875 68570
rect 20927 68518 20939 68570
rect 20991 68518 21003 68570
rect 21055 68518 21067 68570
rect 21119 68518 30820 68570
rect 1104 68496 30820 68518
rect 1394 68416 1400 68468
rect 1452 68456 1458 68468
rect 12802 68456 12808 68468
rect 1452 68428 12808 68456
rect 1452 68416 1458 68428
rect 12802 68416 12808 68428
rect 12860 68416 12866 68468
rect 13357 68459 13415 68465
rect 13357 68425 13369 68459
rect 13403 68456 13415 68459
rect 13906 68456 13912 68468
rect 13403 68428 13912 68456
rect 13403 68425 13415 68428
rect 13357 68419 13415 68425
rect 13906 68416 13912 68428
rect 13964 68416 13970 68468
rect 16298 68456 16304 68468
rect 14108 68428 16304 68456
rect 13173 68323 13231 68329
rect 13173 68289 13185 68323
rect 13219 68320 13231 68323
rect 13814 68320 13820 68332
rect 13219 68292 13820 68320
rect 13219 68289 13231 68292
rect 13173 68283 13231 68289
rect 13814 68280 13820 68292
rect 13872 68280 13878 68332
rect 14108 68329 14136 68428
rect 16298 68416 16304 68428
rect 16356 68416 16362 68468
rect 20438 68416 20444 68468
rect 20496 68456 20502 68468
rect 20533 68459 20591 68465
rect 20533 68456 20545 68459
rect 20496 68428 20545 68456
rect 20496 68416 20502 68428
rect 20533 68425 20545 68428
rect 20579 68425 20591 68459
rect 20533 68419 20591 68425
rect 26973 68459 27031 68465
rect 26973 68425 26985 68459
rect 27019 68456 27031 68459
rect 29454 68456 29460 68468
rect 27019 68428 29460 68456
rect 27019 68425 27031 68428
rect 26973 68419 27031 68425
rect 29454 68416 29460 68428
rect 29512 68416 29518 68468
rect 15194 68388 15200 68400
rect 14292 68360 15200 68388
rect 14292 68329 14320 68360
rect 15194 68348 15200 68360
rect 15252 68348 15258 68400
rect 17313 68391 17371 68397
rect 17313 68357 17325 68391
rect 17359 68388 17371 68391
rect 18230 68388 18236 68400
rect 17359 68360 18236 68388
rect 17359 68357 17371 68360
rect 17313 68351 17371 68357
rect 18230 68348 18236 68360
rect 18288 68348 18294 68400
rect 19518 68388 19524 68400
rect 19479 68360 19524 68388
rect 19518 68348 19524 68360
rect 19576 68348 19582 68400
rect 20346 68388 20352 68400
rect 20307 68360 20352 68388
rect 20346 68348 20352 68360
rect 20404 68348 20410 68400
rect 27080 68360 27381 68388
rect 14073 68323 14136 68329
rect 14073 68289 14085 68323
rect 14119 68292 14136 68323
rect 14182 68323 14240 68329
rect 14119 68289 14131 68292
rect 14073 68283 14131 68289
rect 14182 68289 14194 68323
rect 14228 68289 14240 68323
rect 14292 68323 14356 68329
rect 14292 68292 14310 68323
rect 14182 68283 14240 68289
rect 14298 68289 14310 68292
rect 14344 68289 14356 68323
rect 14458 68320 14464 68332
rect 14419 68292 14464 68320
rect 14298 68283 14356 68289
rect 14200 68196 14228 68283
rect 14458 68280 14464 68292
rect 14516 68280 14522 68332
rect 19337 68323 19395 68329
rect 19337 68289 19349 68323
rect 19383 68320 19395 68323
rect 20714 68320 20720 68332
rect 19383 68292 20720 68320
rect 19383 68289 19395 68292
rect 19337 68283 19395 68289
rect 20714 68280 20720 68292
rect 20772 68280 20778 68332
rect 26418 68280 26424 68332
rect 26476 68320 26482 68332
rect 27080 68320 27108 68360
rect 27353 68329 27381 68360
rect 26476 68292 27108 68320
rect 27203 68323 27261 68329
rect 26476 68280 26482 68292
rect 27203 68289 27215 68323
rect 27249 68289 27261 68323
rect 27203 68283 27261 68289
rect 27341 68323 27399 68329
rect 27341 68289 27353 68323
rect 27387 68289 27399 68323
rect 27341 68283 27399 68289
rect 27433 68326 27491 68329
rect 27522 68326 27528 68332
rect 27433 68323 27528 68326
rect 27433 68289 27445 68323
rect 27479 68298 27528 68323
rect 27479 68289 27491 68298
rect 27433 68283 27491 68289
rect 14918 68212 14924 68264
rect 14976 68252 14982 68264
rect 14976 68224 20208 68252
rect 14976 68212 14982 68224
rect 13817 68187 13875 68193
rect 13817 68153 13829 68187
rect 13863 68184 13875 68187
rect 13998 68184 14004 68196
rect 13863 68156 14004 68184
rect 13863 68153 13875 68156
rect 13817 68147 13875 68153
rect 13998 68144 14004 68156
rect 14056 68144 14062 68196
rect 14182 68144 14188 68196
rect 14240 68144 14246 68196
rect 20070 68184 20076 68196
rect 20031 68156 20076 68184
rect 20070 68144 20076 68156
rect 20128 68144 20134 68196
rect 20180 68184 20208 68224
rect 20530 68212 20536 68264
rect 20588 68252 20594 68264
rect 20625 68255 20683 68261
rect 20625 68252 20637 68255
rect 20588 68224 20637 68252
rect 20588 68212 20594 68224
rect 20625 68221 20637 68224
rect 20671 68252 20683 68255
rect 21174 68252 21180 68264
rect 20671 68224 21180 68252
rect 20671 68221 20683 68224
rect 20625 68215 20683 68221
rect 21174 68212 21180 68224
rect 21232 68212 21238 68264
rect 27062 68212 27068 68264
rect 27120 68252 27126 68264
rect 27218 68252 27246 68283
rect 27522 68280 27528 68298
rect 27580 68280 27586 68332
rect 27617 68323 27675 68329
rect 27617 68289 27629 68323
rect 27663 68289 27675 68323
rect 27617 68283 27675 68289
rect 29825 68323 29883 68329
rect 29825 68289 29837 68323
rect 29871 68320 29883 68323
rect 30466 68320 30472 68332
rect 29871 68292 30472 68320
rect 29871 68289 29883 68292
rect 29825 68283 29883 68289
rect 27120 68224 27246 68252
rect 27120 68212 27126 68224
rect 22462 68184 22468 68196
rect 20180 68156 22468 68184
rect 22462 68144 22468 68156
rect 22520 68144 22526 68196
rect 26510 68144 26516 68196
rect 26568 68184 26574 68196
rect 26568 68156 27246 68184
rect 26568 68144 26574 68156
rect 17310 68076 17316 68128
rect 17368 68116 17374 68128
rect 17405 68119 17463 68125
rect 17405 68116 17417 68119
rect 17368 68088 17417 68116
rect 17368 68076 17374 68088
rect 17405 68085 17417 68088
rect 17451 68085 17463 68119
rect 27218 68116 27246 68156
rect 27632 68116 27660 68283
rect 30466 68280 30472 68292
rect 30524 68280 30530 68332
rect 27218 68088 27660 68116
rect 17405 68079 17463 68085
rect 29914 68076 29920 68128
rect 29972 68116 29978 68128
rect 30009 68119 30067 68125
rect 30009 68116 30021 68119
rect 29972 68088 30021 68116
rect 29972 68076 29978 68088
rect 30009 68085 30021 68088
rect 30055 68085 30067 68119
rect 30009 68079 30067 68085
rect 1104 68026 30820 68048
rect 1104 67974 5915 68026
rect 5967 67974 5979 68026
rect 6031 67974 6043 68026
rect 6095 67974 6107 68026
rect 6159 67974 6171 68026
rect 6223 67974 15846 68026
rect 15898 67974 15910 68026
rect 15962 67974 15974 68026
rect 16026 67974 16038 68026
rect 16090 67974 16102 68026
rect 16154 67974 25776 68026
rect 25828 67974 25840 68026
rect 25892 67974 25904 68026
rect 25956 67974 25968 68026
rect 26020 67974 26032 68026
rect 26084 67974 30820 68026
rect 1104 67952 30820 67974
rect 18138 67872 18144 67924
rect 18196 67912 18202 67924
rect 18509 67915 18567 67921
rect 18509 67912 18521 67915
rect 18196 67884 18521 67912
rect 18196 67872 18202 67884
rect 18509 67881 18521 67884
rect 18555 67881 18567 67915
rect 26234 67912 26240 67924
rect 26195 67884 26240 67912
rect 18509 67875 18567 67881
rect 26234 67872 26240 67884
rect 26292 67872 26298 67924
rect 27341 67915 27399 67921
rect 27341 67881 27353 67915
rect 27387 67912 27399 67915
rect 27430 67912 27436 67924
rect 27387 67884 27436 67912
rect 27387 67881 27399 67884
rect 27341 67875 27399 67881
rect 27430 67872 27436 67884
rect 27488 67872 27494 67924
rect 1397 67847 1455 67853
rect 1397 67813 1409 67847
rect 1443 67844 1455 67847
rect 11238 67844 11244 67856
rect 1443 67816 11244 67844
rect 1443 67813 1455 67816
rect 1397 67807 1455 67813
rect 11238 67804 11244 67816
rect 11296 67804 11302 67856
rect 21266 67844 21272 67856
rect 21227 67816 21272 67844
rect 21266 67804 21272 67816
rect 21324 67804 21330 67856
rect 24857 67847 24915 67853
rect 24857 67813 24869 67847
rect 24903 67844 24915 67847
rect 26050 67844 26056 67856
rect 24903 67816 26056 67844
rect 24903 67813 24915 67816
rect 24857 67807 24915 67813
rect 26050 67804 26056 67816
rect 26108 67804 26114 67856
rect 26602 67804 26608 67856
rect 26660 67804 26666 67856
rect 27062 67804 27068 67856
rect 27120 67844 27126 67856
rect 27614 67844 27620 67856
rect 27120 67816 27620 67844
rect 27120 67804 27126 67816
rect 27614 67804 27620 67816
rect 27672 67804 27678 67856
rect 28902 67844 28908 67856
rect 28863 67816 28908 67844
rect 28902 67804 28908 67816
rect 28960 67804 28966 67856
rect 30006 67844 30012 67856
rect 29967 67816 30012 67844
rect 30006 67804 30012 67816
rect 30064 67804 30070 67856
rect 1578 67708 1584 67720
rect 1539 67680 1584 67708
rect 1578 67668 1584 67680
rect 1636 67668 1642 67720
rect 11330 67668 11336 67720
rect 11388 67708 11394 67720
rect 12897 67711 12955 67717
rect 12897 67708 12909 67711
rect 11388 67680 12909 67708
rect 11388 67668 11394 67680
rect 12897 67677 12909 67680
rect 12943 67677 12955 67711
rect 16666 67708 16672 67720
rect 16627 67680 16672 67708
rect 12897 67671 12955 67677
rect 16666 67668 16672 67680
rect 16724 67668 16730 67720
rect 17402 67708 17408 67720
rect 17363 67680 17408 67708
rect 17402 67668 17408 67680
rect 17460 67668 17466 67720
rect 18325 67711 18383 67717
rect 18325 67677 18337 67711
rect 18371 67708 18383 67711
rect 18690 67708 18696 67720
rect 18371 67680 18696 67708
rect 18371 67677 18383 67680
rect 18325 67671 18383 67677
rect 18690 67668 18696 67680
rect 18748 67668 18754 67720
rect 25041 67711 25099 67717
rect 25041 67677 25053 67711
rect 25087 67708 25099 67711
rect 25130 67708 25136 67720
rect 25087 67680 25136 67708
rect 25087 67677 25099 67680
rect 25041 67671 25099 67677
rect 25130 67668 25136 67680
rect 25188 67668 25194 67720
rect 25317 67711 25375 67717
rect 25317 67677 25329 67711
rect 25363 67708 25375 67711
rect 25406 67708 25412 67720
rect 25363 67680 25412 67708
rect 25363 67677 25375 67680
rect 25317 67671 25375 67677
rect 25406 67668 25412 67680
rect 25464 67668 25470 67720
rect 26620 67717 26648 67804
rect 27264 67748 28028 67776
rect 26493 67711 26551 67717
rect 26493 67677 26505 67711
rect 26539 67708 26551 67711
rect 26602 67711 26660 67717
rect 26539 67677 26556 67708
rect 26493 67671 26556 67677
rect 26602 67677 26614 67711
rect 26648 67677 26660 67711
rect 26602 67671 26660 67677
rect 12618 67600 12624 67652
rect 12676 67640 12682 67652
rect 12713 67643 12771 67649
rect 12713 67640 12725 67643
rect 12676 67612 12725 67640
rect 12676 67600 12682 67612
rect 12713 67609 12725 67612
rect 12759 67609 12771 67643
rect 17586 67640 17592 67652
rect 17547 67612 17592 67640
rect 12713 67603 12771 67609
rect 17586 67600 17592 67612
rect 17644 67600 17650 67652
rect 19978 67640 19984 67652
rect 19939 67612 19984 67640
rect 19978 67600 19984 67612
rect 20036 67600 20042 67652
rect 24946 67600 24952 67652
rect 25004 67640 25010 67652
rect 25222 67640 25228 67652
rect 25004 67612 25228 67640
rect 25004 67600 25010 67612
rect 25222 67600 25228 67612
rect 25280 67600 25286 67652
rect 26528 67640 26556 67671
rect 26694 67668 26700 67720
rect 26752 67708 26758 67720
rect 26752 67680 26797 67708
rect 26752 67668 26758 67680
rect 26878 67668 26884 67720
rect 26936 67708 26942 67720
rect 26936 67680 26981 67708
rect 26936 67668 26942 67680
rect 27062 67668 27068 67720
rect 27120 67708 27126 67720
rect 27264 67708 27292 67748
rect 27614 67708 27620 67720
rect 27120 67680 27292 67708
rect 27575 67680 27620 67708
rect 27120 67668 27126 67680
rect 27614 67668 27620 67680
rect 27672 67668 27678 67720
rect 27709 67711 27767 67717
rect 27709 67677 27721 67711
rect 27755 67677 27767 67711
rect 27709 67671 27767 67677
rect 26528 67612 26648 67640
rect 13078 67572 13084 67584
rect 13039 67544 13084 67572
rect 13078 67532 13084 67544
rect 13136 67532 13142 67584
rect 15194 67532 15200 67584
rect 15252 67572 15258 67584
rect 16761 67575 16819 67581
rect 16761 67572 16773 67575
rect 15252 67544 16773 67572
rect 15252 67532 15258 67544
rect 16761 67541 16773 67544
rect 16807 67572 16819 67575
rect 17678 67572 17684 67584
rect 16807 67544 17684 67572
rect 16807 67541 16819 67544
rect 16761 67535 16819 67541
rect 17678 67532 17684 67544
rect 17736 67532 17742 67584
rect 25590 67532 25596 67584
rect 25648 67572 25654 67584
rect 26142 67572 26148 67584
rect 25648 67544 26148 67572
rect 25648 67532 25654 67544
rect 26142 67532 26148 67544
rect 26200 67532 26206 67584
rect 26620 67572 26648 67612
rect 27614 67572 27620 67584
rect 26620 67544 27620 67572
rect 27614 67532 27620 67544
rect 27672 67532 27678 67584
rect 27724 67572 27752 67671
rect 27798 67668 27804 67720
rect 27856 67708 27862 67720
rect 28000 67717 28028 67748
rect 27985 67711 28043 67717
rect 27856 67680 27901 67708
rect 27856 67668 27862 67680
rect 27985 67677 27997 67711
rect 28031 67677 28043 67711
rect 27985 67671 28043 67677
rect 28721 67711 28779 67717
rect 28721 67677 28733 67711
rect 28767 67708 28779 67711
rect 28994 67708 29000 67720
rect 28767 67680 29000 67708
rect 28767 67677 28779 67680
rect 28721 67671 28779 67677
rect 28994 67668 29000 67680
rect 29052 67668 29058 67720
rect 29454 67668 29460 67720
rect 29512 67708 29518 67720
rect 29825 67711 29883 67717
rect 29825 67708 29837 67711
rect 29512 67680 29837 67708
rect 29512 67668 29518 67680
rect 29825 67677 29837 67680
rect 29871 67677 29883 67711
rect 29825 67671 29883 67677
rect 27798 67572 27804 67584
rect 27724 67544 27804 67572
rect 27798 67532 27804 67544
rect 27856 67532 27862 67584
rect 1104 67482 30820 67504
rect 1104 67430 10880 67482
rect 10932 67430 10944 67482
rect 10996 67430 11008 67482
rect 11060 67430 11072 67482
rect 11124 67430 11136 67482
rect 11188 67430 20811 67482
rect 20863 67430 20875 67482
rect 20927 67430 20939 67482
rect 20991 67430 21003 67482
rect 21055 67430 21067 67482
rect 21119 67430 30820 67482
rect 1104 67408 30820 67430
rect 18598 67328 18604 67380
rect 18656 67368 18662 67380
rect 19153 67371 19211 67377
rect 19153 67368 19165 67371
rect 18656 67340 19165 67368
rect 18656 67328 18662 67340
rect 19153 67337 19165 67340
rect 19199 67337 19211 67371
rect 19153 67331 19211 67337
rect 24857 67371 24915 67377
rect 24857 67337 24869 67371
rect 24903 67368 24915 67371
rect 26878 67368 26884 67380
rect 24903 67340 26884 67368
rect 24903 67337 24915 67340
rect 24857 67331 24915 67337
rect 26878 67328 26884 67340
rect 26936 67328 26942 67380
rect 27614 67368 27620 67380
rect 27264 67340 27620 67368
rect 11238 67260 11244 67312
rect 11296 67300 11302 67312
rect 12805 67303 12863 67309
rect 12805 67300 12817 67303
rect 11296 67272 12817 67300
rect 11296 67260 11302 67272
rect 12805 67269 12817 67272
rect 12851 67269 12863 67303
rect 12805 67263 12863 67269
rect 13078 67260 13084 67312
rect 13136 67300 13142 67312
rect 18969 67303 19027 67309
rect 13136 67272 15516 67300
rect 13136 67260 13142 67272
rect 1578 67232 1584 67244
rect 1539 67204 1584 67232
rect 1578 67192 1584 67204
rect 1636 67192 1642 67244
rect 12618 67232 12624 67244
rect 12579 67204 12624 67232
rect 12618 67192 12624 67204
rect 12676 67192 12682 67244
rect 14918 67192 14924 67244
rect 14976 67232 14982 67244
rect 15488 67241 15516 67272
rect 18969 67269 18981 67303
rect 19015 67300 19027 67303
rect 19518 67300 19524 67312
rect 19015 67272 19524 67300
rect 19015 67269 19027 67272
rect 18969 67263 19027 67269
rect 19518 67260 19524 67272
rect 19576 67260 19582 67312
rect 25148 67272 26004 67300
rect 25148 67244 25176 67272
rect 15059 67235 15117 67241
rect 15059 67232 15071 67235
rect 14976 67204 15071 67232
rect 14976 67192 14982 67204
rect 15059 67201 15071 67204
rect 15105 67201 15117 67235
rect 15059 67195 15117 67201
rect 15194 67235 15252 67241
rect 15194 67201 15206 67235
rect 15240 67201 15252 67235
rect 15194 67195 15252 67201
rect 15294 67235 15352 67241
rect 15294 67201 15306 67235
rect 15340 67201 15352 67235
rect 15294 67195 15352 67201
rect 15473 67235 15531 67241
rect 15473 67201 15485 67235
rect 15519 67201 15531 67235
rect 15473 67195 15531 67201
rect 14182 67124 14188 67176
rect 14240 67164 14246 67176
rect 15212 67164 15240 67195
rect 14240 67136 15240 67164
rect 14240 67124 14246 67136
rect 14550 67056 14556 67108
rect 14608 67096 14614 67108
rect 15194 67096 15200 67108
rect 14608 67068 15200 67096
rect 14608 67056 14614 67068
rect 15194 67056 15200 67068
rect 15252 67096 15258 67108
rect 15304 67096 15332 67195
rect 19702 67192 19708 67244
rect 19760 67232 19766 67244
rect 23293 67235 23351 67241
rect 23293 67232 23305 67235
rect 19760 67204 23305 67232
rect 19760 67192 19766 67204
rect 23293 67201 23305 67204
rect 23339 67201 23351 67235
rect 23293 67195 23351 67201
rect 23477 67235 23535 67241
rect 23477 67201 23489 67235
rect 23523 67232 23535 67235
rect 23566 67232 23572 67244
rect 23523 67204 23572 67232
rect 23523 67201 23535 67204
rect 23477 67195 23535 67201
rect 23566 67192 23572 67204
rect 23624 67192 23630 67244
rect 25041 67235 25099 67241
rect 25041 67201 25053 67235
rect 25087 67232 25099 67235
rect 25130 67232 25136 67244
rect 25087 67204 25136 67232
rect 25087 67201 25099 67204
rect 25041 67195 25099 67201
rect 25130 67192 25136 67204
rect 25188 67192 25194 67244
rect 25225 67235 25283 67241
rect 25225 67201 25237 67235
rect 25271 67201 25283 67235
rect 25225 67195 25283 67201
rect 25317 67235 25375 67241
rect 25317 67201 25329 67235
rect 25363 67232 25375 67235
rect 25406 67232 25412 67244
rect 25363 67204 25412 67232
rect 25363 67201 25375 67204
rect 25317 67195 25375 67201
rect 17034 67124 17040 67176
rect 17092 67164 17098 67176
rect 19245 67167 19303 67173
rect 17092 67136 18828 67164
rect 17092 67124 17098 67136
rect 18690 67096 18696 67108
rect 15252 67068 15332 67096
rect 18651 67068 18696 67096
rect 15252 67056 15258 67068
rect 18690 67056 18696 67068
rect 18748 67056 18754 67108
rect 18800 67096 18828 67136
rect 19245 67133 19257 67167
rect 19291 67164 19303 67167
rect 19886 67164 19892 67176
rect 19291 67136 19892 67164
rect 19291 67133 19303 67136
rect 19245 67127 19303 67133
rect 19886 67124 19892 67136
rect 19944 67164 19950 67176
rect 20070 67164 20076 67176
rect 19944 67136 20076 67164
rect 19944 67124 19950 67136
rect 20070 67124 20076 67136
rect 20128 67124 20134 67176
rect 25240 67164 25268 67195
rect 25406 67192 25412 67204
rect 25464 67192 25470 67244
rect 25976 67241 26004 67272
rect 25961 67235 26019 67241
rect 25961 67201 25973 67235
rect 26007 67201 26019 67235
rect 25961 67195 26019 67201
rect 26050 67192 26056 67244
rect 26108 67232 26114 67244
rect 26145 67235 26203 67241
rect 26145 67232 26157 67235
rect 26108 67204 26157 67232
rect 26108 67192 26114 67204
rect 26145 67201 26157 67204
rect 26191 67201 26203 67235
rect 26145 67195 26203 67201
rect 26234 67192 26240 67244
rect 26292 67232 26298 67244
rect 27264 67241 27292 67340
rect 27614 67328 27620 67340
rect 27672 67368 27678 67380
rect 27798 67368 27804 67380
rect 27672 67340 27804 67368
rect 27672 67328 27678 67340
rect 27798 67328 27804 67340
rect 27856 67328 27862 67380
rect 27890 67300 27896 67312
rect 27377 67272 27896 67300
rect 27377 67241 27405 67272
rect 27890 67260 27896 67272
rect 27948 67260 27954 67312
rect 27249 67235 27307 67241
rect 26292 67204 26337 67232
rect 26292 67192 26298 67204
rect 27249 67201 27261 67235
rect 27295 67201 27307 67235
rect 27249 67195 27307 67201
rect 27338 67235 27405 67241
rect 27338 67201 27350 67235
rect 27384 67204 27405 67235
rect 27438 67235 27496 67241
rect 27384 67201 27396 67204
rect 27338 67195 27396 67201
rect 27438 67201 27450 67235
rect 27484 67201 27496 67235
rect 27614 67232 27620 67244
rect 27575 67204 27620 67232
rect 27438 67195 27496 67201
rect 25498 67164 25504 67176
rect 25056 67136 25268 67164
rect 25424 67136 25504 67164
rect 25056 67108 25084 67136
rect 25038 67096 25044 67108
rect 18800 67068 25044 67096
rect 25038 67056 25044 67068
rect 25096 67056 25102 67108
rect 1397 67031 1455 67037
rect 1397 66997 1409 67031
rect 1443 67028 1455 67031
rect 11238 67028 11244 67040
rect 1443 67000 11244 67028
rect 1443 66997 1455 67000
rect 1397 66991 1455 66997
rect 11238 66988 11244 67000
rect 11296 66988 11302 67040
rect 12989 67031 13047 67037
rect 12989 66997 13001 67031
rect 13035 67028 13047 67031
rect 14734 67028 14740 67040
rect 13035 67000 14740 67028
rect 13035 66997 13047 67000
rect 12989 66991 13047 66997
rect 14734 66988 14740 67000
rect 14792 66988 14798 67040
rect 14829 67031 14887 67037
rect 14829 66997 14841 67031
rect 14875 67028 14887 67031
rect 15378 67028 15384 67040
rect 14875 67000 15384 67028
rect 14875 66997 14887 67000
rect 14829 66991 14887 66997
rect 15378 66988 15384 67000
rect 15436 66988 15442 67040
rect 23661 67031 23719 67037
rect 23661 66997 23673 67031
rect 23707 67028 23719 67031
rect 23934 67028 23940 67040
rect 23707 67000 23940 67028
rect 23707 66997 23719 67000
rect 23661 66991 23719 66997
rect 23934 66988 23940 67000
rect 23992 66988 23998 67040
rect 24854 66988 24860 67040
rect 24912 67028 24918 67040
rect 25424 67028 25452 67136
rect 25498 67124 25504 67136
rect 25556 67124 25562 67176
rect 25777 67167 25835 67173
rect 25777 67133 25789 67167
rect 25823 67164 25835 67167
rect 27062 67164 27068 67176
rect 25823 67136 27068 67164
rect 25823 67133 25835 67136
rect 25777 67127 25835 67133
rect 27062 67124 27068 67136
rect 27120 67124 27126 67176
rect 27445 67164 27473 67195
rect 27614 67192 27620 67204
rect 27672 67192 27678 67244
rect 28258 67192 28264 67244
rect 28316 67232 28322 67244
rect 29089 67235 29147 67241
rect 29089 67232 29101 67235
rect 28316 67204 29101 67232
rect 28316 67192 28322 67204
rect 29089 67201 29101 67204
rect 29135 67201 29147 67235
rect 29089 67195 29147 67201
rect 29825 67235 29883 67241
rect 29825 67201 29837 67235
rect 29871 67201 29883 67235
rect 29825 67195 29883 67201
rect 29840 67164 29868 67195
rect 27172 67136 27473 67164
rect 27540 67136 29868 67164
rect 26878 67056 26884 67108
rect 26936 67096 26942 67108
rect 27172 67096 27200 67136
rect 26936 67068 27200 67096
rect 26936 67056 26942 67068
rect 27430 67056 27436 67108
rect 27488 67096 27494 67108
rect 27540 67096 27568 67136
rect 29086 67096 29092 67108
rect 27488 67068 27568 67096
rect 28276 67068 29092 67096
rect 27488 67056 27494 67068
rect 24912 67000 25452 67028
rect 26973 67031 27031 67037
rect 24912 66988 24918 67000
rect 26973 66997 26985 67031
rect 27019 67028 27031 67031
rect 28276 67028 28304 67068
rect 29086 67056 29092 67068
rect 29144 67056 29150 67108
rect 27019 67000 28304 67028
rect 27019 66997 27031 67000
rect 26973 66991 27031 66997
rect 28902 66988 28908 67040
rect 28960 67028 28966 67040
rect 29273 67031 29331 67037
rect 29273 67028 29285 67031
rect 28960 67000 29285 67028
rect 28960 66988 28966 67000
rect 29273 66997 29285 67000
rect 29319 66997 29331 67031
rect 29273 66991 29331 66997
rect 29822 66988 29828 67040
rect 29880 67028 29886 67040
rect 30009 67031 30067 67037
rect 30009 67028 30021 67031
rect 29880 67000 30021 67028
rect 29880 66988 29886 67000
rect 30009 66997 30021 67000
rect 30055 66997 30067 67031
rect 30009 66991 30067 66997
rect 1104 66938 30820 66960
rect 1104 66886 5915 66938
rect 5967 66886 5979 66938
rect 6031 66886 6043 66938
rect 6095 66886 6107 66938
rect 6159 66886 6171 66938
rect 6223 66886 15846 66938
rect 15898 66886 15910 66938
rect 15962 66886 15974 66938
rect 16026 66886 16038 66938
rect 16090 66886 16102 66938
rect 16154 66886 25776 66938
rect 25828 66886 25840 66938
rect 25892 66886 25904 66938
rect 25956 66886 25968 66938
rect 26020 66886 26032 66938
rect 26084 66886 30820 66938
rect 1104 66864 30820 66886
rect 14918 66784 14924 66836
rect 14976 66824 14982 66836
rect 18414 66824 18420 66836
rect 14976 66796 16712 66824
rect 18375 66796 18420 66824
rect 14976 66784 14982 66796
rect 16684 66765 16712 66796
rect 18414 66784 18420 66796
rect 18472 66784 18478 66836
rect 19429 66827 19487 66833
rect 19429 66793 19441 66827
rect 19475 66824 19487 66827
rect 19610 66824 19616 66836
rect 19475 66796 19616 66824
rect 19475 66793 19487 66796
rect 19429 66787 19487 66793
rect 19610 66784 19616 66796
rect 19668 66784 19674 66836
rect 22554 66784 22560 66836
rect 22612 66824 22618 66836
rect 23566 66824 23572 66836
rect 22612 66796 23572 66824
rect 22612 66784 22618 66796
rect 23566 66784 23572 66796
rect 23624 66784 23630 66836
rect 26421 66827 26479 66833
rect 26421 66793 26433 66827
rect 26467 66824 26479 66827
rect 26970 66824 26976 66836
rect 26467 66796 26976 66824
rect 26467 66793 26479 66796
rect 26421 66787 26479 66793
rect 26970 66784 26976 66796
rect 27028 66784 27034 66836
rect 28810 66784 28816 66836
rect 28868 66824 28874 66836
rect 29086 66824 29092 66836
rect 28868 66796 29092 66824
rect 28868 66784 28874 66796
rect 29086 66784 29092 66796
rect 29144 66784 29150 66836
rect 16669 66759 16727 66765
rect 16669 66725 16681 66759
rect 16715 66756 16727 66759
rect 23290 66756 23296 66768
rect 16715 66728 23296 66756
rect 16715 66725 16727 66728
rect 16669 66719 16727 66725
rect 23290 66716 23296 66728
rect 23348 66716 23354 66768
rect 25317 66759 25375 66765
rect 25317 66725 25329 66759
rect 25363 66756 25375 66759
rect 26510 66756 26516 66768
rect 25363 66728 26516 66756
rect 25363 66725 25375 66728
rect 25317 66719 25375 66725
rect 26510 66716 26516 66728
rect 26568 66716 26574 66768
rect 26620 66728 27844 66756
rect 14182 66648 14188 66700
rect 14240 66688 14246 66700
rect 14240 66660 14504 66688
rect 14240 66648 14246 66660
rect 1578 66620 1584 66632
rect 1539 66592 1584 66620
rect 1578 66580 1584 66592
rect 1636 66580 1642 66632
rect 14476 66629 14504 66660
rect 16390 66648 16396 66700
rect 16448 66688 16454 66700
rect 16448 66660 17816 66688
rect 16448 66648 16454 66660
rect 14369 66623 14427 66629
rect 14369 66589 14381 66623
rect 14415 66589 14427 66623
rect 14369 66583 14427 66589
rect 14461 66623 14519 66629
rect 14461 66589 14473 66623
rect 14507 66589 14519 66623
rect 14461 66583 14519 66589
rect 14384 66552 14412 66583
rect 14550 66580 14556 66632
rect 14608 66620 14614 66632
rect 14734 66620 14740 66632
rect 14608 66592 14653 66620
rect 14695 66592 14740 66620
rect 14608 66580 14614 66592
rect 14734 66580 14740 66592
rect 14792 66580 14798 66632
rect 15286 66620 15292 66632
rect 15247 66592 15292 66620
rect 15286 66580 15292 66592
rect 15344 66580 15350 66632
rect 15378 66580 15384 66632
rect 15436 66620 15442 66632
rect 15545 66623 15603 66629
rect 15545 66620 15557 66623
rect 15436 66592 15557 66620
rect 15436 66580 15442 66592
rect 15545 66589 15557 66592
rect 15591 66589 15603 66623
rect 15545 66583 15603 66589
rect 17385 66623 17443 66629
rect 17385 66589 17397 66623
rect 17431 66620 17443 66623
rect 17497 66623 17555 66629
rect 17431 66589 17448 66620
rect 17385 66583 17448 66589
rect 17497 66589 17509 66623
rect 17543 66589 17555 66623
rect 17497 66583 17555 66589
rect 17589 66623 17647 66629
rect 17589 66589 17601 66623
rect 17635 66620 17647 66623
rect 17678 66620 17684 66632
rect 17635 66592 17684 66620
rect 17635 66589 17647 66592
rect 17589 66583 17647 66589
rect 14826 66552 14832 66564
rect 14384 66524 14832 66552
rect 14826 66512 14832 66524
rect 14884 66512 14890 66564
rect 1397 66487 1455 66493
rect 1397 66453 1409 66487
rect 1443 66484 1455 66487
rect 11330 66484 11336 66496
rect 1443 66456 11336 66484
rect 1443 66453 1455 66456
rect 1397 66447 1455 66453
rect 11330 66444 11336 66456
rect 11388 66444 11394 66496
rect 14090 66484 14096 66496
rect 14051 66456 14096 66484
rect 14090 66444 14096 66456
rect 14148 66444 14154 66496
rect 17126 66484 17132 66496
rect 17087 66456 17132 66484
rect 17126 66444 17132 66456
rect 17184 66444 17190 66496
rect 17420 66484 17448 66583
rect 17512 66552 17540 66583
rect 17678 66580 17684 66592
rect 17736 66580 17742 66632
rect 17788 66629 17816 66660
rect 18322 66648 18328 66700
rect 18380 66688 18386 66700
rect 18380 66660 20116 66688
rect 18380 66648 18386 66660
rect 17773 66623 17831 66629
rect 17773 66589 17785 66623
rect 17819 66589 17831 66623
rect 17773 66583 17831 66589
rect 18233 66623 18291 66629
rect 18233 66589 18245 66623
rect 18279 66620 18291 66623
rect 18598 66620 18604 66632
rect 18279 66592 18604 66620
rect 18279 66589 18291 66592
rect 18233 66583 18291 66589
rect 18598 66580 18604 66592
rect 18656 66620 18662 66632
rect 19245 66623 19303 66629
rect 19245 66620 19257 66623
rect 18656 66592 19257 66620
rect 18656 66580 18662 66592
rect 19245 66589 19257 66592
rect 19291 66589 19303 66623
rect 19245 66583 19303 66589
rect 17862 66552 17868 66564
rect 17512 66524 17868 66552
rect 17862 66512 17868 66524
rect 17920 66512 17926 66564
rect 20088 66552 20116 66660
rect 20162 66648 20168 66700
rect 20220 66688 20226 66700
rect 22373 66691 22431 66697
rect 22373 66688 22385 66691
rect 20220 66660 22385 66688
rect 20220 66648 20226 66660
rect 22373 66657 22385 66660
rect 22419 66657 22431 66691
rect 22373 66651 22431 66657
rect 22830 66648 22836 66700
rect 22888 66688 22894 66700
rect 24397 66691 24455 66697
rect 24397 66688 24409 66691
rect 22888 66660 24409 66688
rect 22888 66648 22894 66660
rect 24397 66657 24409 66660
rect 24443 66657 24455 66691
rect 24397 66651 24455 66657
rect 20530 66620 20536 66632
rect 20491 66592 20536 66620
rect 20530 66580 20536 66592
rect 20588 66580 20594 66632
rect 22554 66620 22560 66632
rect 22515 66592 22560 66620
rect 22554 66580 22560 66592
rect 22612 66580 22618 66632
rect 23385 66623 23443 66629
rect 23385 66589 23397 66623
rect 23431 66589 23443 66623
rect 23385 66583 23443 66589
rect 23477 66623 23535 66629
rect 23477 66589 23489 66623
rect 23523 66620 23535 66623
rect 23566 66620 23572 66632
rect 23523 66592 23572 66620
rect 23523 66589 23535 66592
rect 23477 66583 23535 66589
rect 23400 66552 23428 66583
rect 23566 66580 23572 66592
rect 23624 66620 23630 66632
rect 24581 66623 24639 66629
rect 24581 66620 24593 66623
rect 23624 66592 24593 66620
rect 23624 66580 23630 66592
rect 24581 66589 24593 66592
rect 24627 66589 24639 66623
rect 24581 66583 24639 66589
rect 25222 66580 25228 66632
rect 25280 66620 25286 66632
rect 25501 66623 25559 66629
rect 25501 66620 25513 66623
rect 25280 66592 25513 66620
rect 25280 66580 25286 66592
rect 25501 66589 25513 66592
rect 25547 66589 25559 66623
rect 25501 66583 25559 66589
rect 25777 66623 25835 66629
rect 25777 66589 25789 66623
rect 25823 66620 25835 66623
rect 26142 66620 26148 66632
rect 25823 66592 26148 66620
rect 25823 66589 25835 66592
rect 25777 66583 25835 66589
rect 20088 66524 23428 66552
rect 24210 66512 24216 66564
rect 24268 66552 24274 66564
rect 24268 66524 24900 66552
rect 24268 66512 24274 66524
rect 18414 66484 18420 66496
rect 17420 66456 18420 66484
rect 18414 66444 18420 66456
rect 18472 66444 18478 66496
rect 20714 66484 20720 66496
rect 20675 66456 20720 66484
rect 20714 66444 20720 66456
rect 20772 66444 20778 66496
rect 22741 66487 22799 66493
rect 22741 66453 22753 66487
rect 22787 66484 22799 66487
rect 23382 66484 23388 66496
rect 22787 66456 23388 66484
rect 22787 66453 22799 66456
rect 22741 66447 22799 66453
rect 23382 66444 23388 66456
rect 23440 66444 23446 66496
rect 23658 66484 23664 66496
rect 23619 66456 23664 66484
rect 23658 66444 23664 66456
rect 23716 66444 23722 66496
rect 24670 66444 24676 66496
rect 24728 66484 24734 66496
rect 24765 66487 24823 66493
rect 24765 66484 24777 66487
rect 24728 66456 24777 66484
rect 24728 66444 24734 66456
rect 24765 66453 24777 66456
rect 24811 66453 24823 66487
rect 24872 66484 24900 66524
rect 25130 66512 25136 66564
rect 25188 66552 25194 66564
rect 25406 66552 25412 66564
rect 25188 66524 25412 66552
rect 25188 66512 25194 66524
rect 25406 66512 25412 66524
rect 25464 66552 25470 66564
rect 25792 66552 25820 66583
rect 26142 66580 26148 66592
rect 26200 66580 26206 66632
rect 26620 66622 26648 66728
rect 27816 66700 27844 66728
rect 27246 66688 27252 66700
rect 26896 66660 27252 66688
rect 26896 66629 26924 66660
rect 27246 66648 27252 66660
rect 27304 66648 27310 66700
rect 27614 66688 27620 66700
rect 27448 66660 27620 66688
rect 26697 66623 26755 66629
rect 26697 66622 26709 66623
rect 26620 66594 26709 66622
rect 26697 66589 26709 66594
rect 26743 66589 26755 66623
rect 26697 66583 26755 66589
rect 26789 66623 26847 66629
rect 26789 66589 26801 66623
rect 26835 66589 26847 66623
rect 26789 66583 26847 66589
rect 26881 66623 26939 66629
rect 26881 66589 26893 66623
rect 26927 66589 26939 66623
rect 26881 66583 26939 66589
rect 25464 66524 25820 66552
rect 26804 66552 26832 66583
rect 26970 66580 26976 66632
rect 27028 66580 27034 66632
rect 27077 66623 27135 66629
rect 27077 66589 27089 66623
rect 27123 66620 27135 66623
rect 27448 66620 27476 66660
rect 27614 66648 27620 66660
rect 27672 66648 27678 66700
rect 27798 66688 27804 66700
rect 27759 66660 27804 66688
rect 27798 66648 27804 66660
rect 27856 66648 27862 66700
rect 27123 66592 27476 66620
rect 27525 66623 27583 66629
rect 27123 66589 27135 66592
rect 27077 66583 27135 66589
rect 27525 66589 27537 66623
rect 27571 66589 27583 66623
rect 27525 66583 27583 66589
rect 26988 66552 27016 66580
rect 26804 66524 27016 66552
rect 27540 66552 27568 66583
rect 28810 66580 28816 66632
rect 28868 66620 28874 66632
rect 29825 66623 29883 66629
rect 29825 66620 29837 66623
rect 28868 66592 29837 66620
rect 28868 66580 28874 66592
rect 29825 66589 29837 66592
rect 29871 66589 29883 66623
rect 29825 66583 29883 66589
rect 27798 66552 27804 66564
rect 27540 66524 27804 66552
rect 25464 66512 25470 66524
rect 27798 66512 27804 66524
rect 27856 66512 27862 66564
rect 25685 66487 25743 66493
rect 25685 66484 25697 66487
rect 24872 66456 25697 66484
rect 24765 66447 24823 66453
rect 25685 66453 25697 66456
rect 25731 66453 25743 66487
rect 25685 66447 25743 66453
rect 26970 66444 26976 66496
rect 27028 66484 27034 66496
rect 30009 66487 30067 66493
rect 30009 66484 30021 66487
rect 27028 66456 30021 66484
rect 27028 66444 27034 66456
rect 30009 66453 30021 66456
rect 30055 66453 30067 66487
rect 30009 66447 30067 66453
rect 1104 66394 30820 66416
rect 1104 66342 10880 66394
rect 10932 66342 10944 66394
rect 10996 66342 11008 66394
rect 11060 66342 11072 66394
rect 11124 66342 11136 66394
rect 11188 66342 20811 66394
rect 20863 66342 20875 66394
rect 20927 66342 20939 66394
rect 20991 66342 21003 66394
rect 21055 66342 21067 66394
rect 21119 66342 30820 66394
rect 1104 66320 30820 66342
rect 25041 66283 25099 66289
rect 25041 66249 25053 66283
rect 25087 66280 25099 66283
rect 27614 66280 27620 66292
rect 25087 66252 27620 66280
rect 25087 66249 25099 66252
rect 25041 66243 25099 66249
rect 27614 66240 27620 66252
rect 27672 66240 27678 66292
rect 29454 66240 29460 66292
rect 29512 66280 29518 66292
rect 29512 66252 30236 66280
rect 29512 66240 29518 66252
rect 11238 66172 11244 66224
rect 11296 66212 11302 66224
rect 12805 66215 12863 66221
rect 12805 66212 12817 66215
rect 11296 66184 12817 66212
rect 11296 66172 11302 66184
rect 12805 66181 12817 66184
rect 12851 66181 12863 66215
rect 12805 66175 12863 66181
rect 13992 66215 14050 66221
rect 13992 66181 14004 66215
rect 14038 66212 14050 66215
rect 14090 66212 14096 66224
rect 14038 66184 14096 66212
rect 14038 66181 14050 66184
rect 13992 66175 14050 66181
rect 14090 66172 14096 66184
rect 14148 66172 14154 66224
rect 17126 66172 17132 66224
rect 17184 66212 17190 66224
rect 17282 66215 17340 66221
rect 17282 66212 17294 66215
rect 17184 66184 17294 66212
rect 17184 66172 17190 66184
rect 17282 66181 17294 66184
rect 17328 66181 17340 66215
rect 22370 66212 22376 66224
rect 17282 66175 17340 66181
rect 22185 66184 22376 66212
rect 22185 66156 22213 66184
rect 22370 66172 22376 66184
rect 22428 66172 22434 66224
rect 23014 66172 23020 66224
rect 23072 66212 23078 66224
rect 23661 66215 23719 66221
rect 23661 66212 23673 66215
rect 23072 66184 23673 66212
rect 23072 66172 23078 66184
rect 23661 66181 23673 66184
rect 23707 66181 23719 66215
rect 30098 66212 30104 66224
rect 30059 66184 30104 66212
rect 23661 66175 23719 66181
rect 30098 66172 30104 66184
rect 30156 66172 30162 66224
rect 1578 66144 1584 66156
rect 1539 66116 1584 66144
rect 1578 66104 1584 66116
rect 1636 66104 1642 66156
rect 12618 66144 12624 66156
rect 12579 66116 12624 66144
rect 12618 66104 12624 66116
rect 12676 66104 12682 66156
rect 15933 66147 15991 66153
rect 15933 66113 15945 66147
rect 15979 66144 15991 66147
rect 16850 66144 16856 66156
rect 15979 66116 16856 66144
rect 15979 66113 15991 66116
rect 15933 66107 15991 66113
rect 16850 66104 16856 66116
rect 16908 66104 16914 66156
rect 18690 66104 18696 66156
rect 18748 66144 18754 66156
rect 19521 66147 19579 66153
rect 19521 66144 19533 66147
rect 18748 66116 19533 66144
rect 18748 66104 18754 66116
rect 19521 66113 19533 66116
rect 19567 66113 19579 66147
rect 19521 66107 19579 66113
rect 21910 66104 21916 66156
rect 21968 66144 21974 66156
rect 22051 66147 22109 66153
rect 22051 66144 22063 66147
rect 21968 66116 22063 66144
rect 21968 66104 21974 66116
rect 22051 66113 22063 66116
rect 22097 66113 22109 66147
rect 22051 66107 22109 66113
rect 22170 66150 22228 66156
rect 22170 66116 22182 66150
rect 22216 66116 22228 66150
rect 22170 66110 22228 66116
rect 22281 66147 22339 66153
rect 22281 66113 22293 66147
rect 22327 66144 22339 66147
rect 22465 66147 22523 66153
rect 22327 66116 22416 66144
rect 22327 66113 22339 66116
rect 22281 66107 22339 66113
rect 22388 66088 22416 66116
rect 22465 66113 22477 66147
rect 22511 66144 22523 66147
rect 22554 66144 22560 66156
rect 22511 66116 22560 66144
rect 22511 66113 22523 66116
rect 22465 66107 22523 66113
rect 22554 66104 22560 66116
rect 22612 66104 22618 66156
rect 23290 66144 23296 66156
rect 23251 66116 23296 66144
rect 23290 66104 23296 66116
rect 23348 66104 23354 66156
rect 23477 66147 23535 66153
rect 23477 66113 23489 66147
rect 23523 66144 23535 66147
rect 23566 66144 23572 66156
rect 23523 66116 23572 66144
rect 23523 66113 23535 66116
rect 23477 66107 23535 66113
rect 23566 66104 23572 66116
rect 23624 66104 23630 66156
rect 25222 66144 25228 66156
rect 25183 66116 25228 66144
rect 25222 66104 25228 66116
rect 25280 66104 25286 66156
rect 25406 66144 25412 66156
rect 25367 66116 25412 66144
rect 25406 66104 25412 66116
rect 25464 66104 25470 66156
rect 25501 66147 25559 66153
rect 25501 66113 25513 66147
rect 25547 66144 25559 66147
rect 26142 66144 26148 66156
rect 25547 66116 26148 66144
rect 25547 66113 25559 66116
rect 25501 66107 25559 66113
rect 26142 66104 26148 66116
rect 26200 66104 26206 66156
rect 27893 66147 27951 66153
rect 27893 66113 27905 66147
rect 27939 66144 27951 66147
rect 27982 66144 27988 66156
rect 27939 66116 27988 66144
rect 27939 66113 27951 66116
rect 27893 66107 27951 66113
rect 27982 66104 27988 66116
rect 28040 66104 28046 66156
rect 28626 66144 28632 66156
rect 28587 66116 28632 66144
rect 28626 66104 28632 66116
rect 28684 66104 28690 66156
rect 28718 66104 28724 66156
rect 28776 66144 28782 66156
rect 29365 66147 29423 66153
rect 29365 66144 29377 66147
rect 28776 66116 29377 66144
rect 28776 66104 28782 66116
rect 29365 66113 29377 66116
rect 29411 66113 29423 66147
rect 29549 66147 29607 66153
rect 29549 66144 29561 66147
rect 29365 66107 29423 66113
rect 29472 66116 29561 66144
rect 13722 66076 13728 66088
rect 13683 66048 13728 66076
rect 13722 66036 13728 66048
rect 13780 66036 13786 66088
rect 17037 66079 17095 66085
rect 17037 66076 17049 66079
rect 16132 66048 17049 66076
rect 16132 66017 16160 66048
rect 17037 66045 17049 66048
rect 17083 66045 17095 66079
rect 17037 66039 17095 66045
rect 22370 66036 22376 66088
rect 22428 66036 22434 66088
rect 28902 66036 28908 66088
rect 28960 66076 28966 66088
rect 29472 66076 29500 66116
rect 29549 66113 29561 66116
rect 29595 66113 29607 66147
rect 29549 66107 29607 66113
rect 29641 66147 29699 66153
rect 29641 66113 29653 66147
rect 29687 66144 29699 66147
rect 29917 66147 29975 66153
rect 29687 66116 29868 66144
rect 29687 66113 29699 66116
rect 29641 66107 29699 66113
rect 28960 66048 29500 66076
rect 29733 66079 29791 66085
rect 28960 66036 28966 66048
rect 29733 66045 29745 66079
rect 29779 66045 29791 66079
rect 29733 66039 29791 66045
rect 16117 66011 16175 66017
rect 16117 65977 16129 66011
rect 16163 65977 16175 66011
rect 16117 65971 16175 65977
rect 20622 65968 20628 66020
rect 20680 66008 20686 66020
rect 20809 66011 20867 66017
rect 20809 66008 20821 66011
rect 20680 65980 20821 66008
rect 20680 65968 20686 65980
rect 20809 65977 20821 65980
rect 20855 65977 20867 66011
rect 20809 65971 20867 65977
rect 20916 65980 22094 66008
rect 1397 65943 1455 65949
rect 1397 65909 1409 65943
rect 1443 65940 1455 65943
rect 11422 65940 11428 65952
rect 1443 65912 11428 65940
rect 1443 65909 1455 65912
rect 1397 65903 1455 65909
rect 11422 65900 11428 65912
rect 11480 65900 11486 65952
rect 12986 65940 12992 65952
rect 12947 65912 12992 65940
rect 12986 65900 12992 65912
rect 13044 65900 13050 65952
rect 14826 65900 14832 65952
rect 14884 65940 14890 65952
rect 15105 65943 15163 65949
rect 15105 65940 15117 65943
rect 14884 65912 15117 65940
rect 14884 65900 14890 65912
rect 15105 65909 15117 65912
rect 15151 65909 15163 65943
rect 18414 65940 18420 65952
rect 18327 65912 18420 65940
rect 15105 65903 15163 65909
rect 18414 65900 18420 65912
rect 18472 65940 18478 65952
rect 20916 65940 20944 65980
rect 21818 65940 21824 65952
rect 18472 65912 20944 65940
rect 21779 65912 21824 65940
rect 18472 65900 18478 65912
rect 21818 65900 21824 65912
rect 21876 65900 21882 65952
rect 22066 65940 22094 65980
rect 25516 65980 28948 66008
rect 23474 65940 23480 65952
rect 22066 65912 23480 65940
rect 23474 65900 23480 65912
rect 23532 65900 23538 65952
rect 24670 65900 24676 65952
rect 24728 65940 24734 65952
rect 25516 65940 25544 65980
rect 28074 65940 28080 65952
rect 24728 65912 25544 65940
rect 28035 65912 28080 65940
rect 24728 65900 24734 65912
rect 28074 65900 28080 65912
rect 28132 65900 28138 65952
rect 28166 65900 28172 65952
rect 28224 65940 28230 65952
rect 28813 65943 28871 65949
rect 28813 65940 28825 65943
rect 28224 65912 28825 65940
rect 28224 65900 28230 65912
rect 28813 65909 28825 65912
rect 28859 65909 28871 65943
rect 28920 65940 28948 65980
rect 29546 65968 29552 66020
rect 29604 66008 29610 66020
rect 29748 66008 29776 66039
rect 29604 65980 29776 66008
rect 29604 65968 29610 65980
rect 29840 65940 29868 66116
rect 29917 66113 29929 66147
rect 29963 66113 29975 66147
rect 29917 66107 29975 66113
rect 29932 66008 29960 66107
rect 30098 66036 30104 66088
rect 30156 66076 30162 66088
rect 30208 66076 30236 66252
rect 30156 66048 30236 66076
rect 30156 66036 30162 66048
rect 30374 66008 30380 66020
rect 29932 65980 30380 66008
rect 30374 65968 30380 65980
rect 30432 65968 30438 66020
rect 29914 65940 29920 65952
rect 28920 65912 29920 65940
rect 28813 65903 28871 65909
rect 29914 65900 29920 65912
rect 29972 65900 29978 65952
rect 1104 65850 30820 65872
rect 1104 65798 5915 65850
rect 5967 65798 5979 65850
rect 6031 65798 6043 65850
rect 6095 65798 6107 65850
rect 6159 65798 6171 65850
rect 6223 65798 15846 65850
rect 15898 65798 15910 65850
rect 15962 65798 15974 65850
rect 16026 65798 16038 65850
rect 16090 65798 16102 65850
rect 16154 65798 25776 65850
rect 25828 65798 25840 65850
rect 25892 65798 25904 65850
rect 25956 65798 25968 65850
rect 26020 65798 26032 65850
rect 26084 65798 30820 65850
rect 1104 65776 30820 65798
rect 12618 65696 12624 65748
rect 12676 65736 12682 65748
rect 12713 65739 12771 65745
rect 12713 65736 12725 65739
rect 12676 65708 12725 65736
rect 12676 65696 12682 65708
rect 12713 65705 12725 65708
rect 12759 65705 12771 65739
rect 12713 65699 12771 65705
rect 15286 65696 15292 65748
rect 15344 65736 15350 65748
rect 15473 65739 15531 65745
rect 15473 65736 15485 65739
rect 15344 65708 15485 65736
rect 15344 65696 15350 65708
rect 15473 65705 15485 65708
rect 15519 65705 15531 65739
rect 16850 65736 16856 65748
rect 16811 65708 16856 65736
rect 15473 65699 15531 65705
rect 16850 65696 16856 65708
rect 16908 65696 16914 65748
rect 18046 65696 18052 65748
rect 18104 65736 18110 65748
rect 18141 65739 18199 65745
rect 18141 65736 18153 65739
rect 18104 65708 18153 65736
rect 18104 65696 18110 65708
rect 18141 65705 18153 65708
rect 18187 65705 18199 65739
rect 19426 65736 19432 65748
rect 19387 65708 19432 65736
rect 18141 65699 18199 65705
rect 19426 65696 19432 65708
rect 19484 65696 19490 65748
rect 19981 65739 20039 65745
rect 19981 65705 19993 65739
rect 20027 65736 20039 65739
rect 20530 65736 20536 65748
rect 20027 65708 20536 65736
rect 20027 65705 20039 65708
rect 19981 65699 20039 65705
rect 20530 65696 20536 65708
rect 20588 65696 20594 65748
rect 27338 65696 27344 65748
rect 27396 65736 27402 65748
rect 27433 65739 27491 65745
rect 27433 65736 27445 65739
rect 27396 65708 27445 65736
rect 27396 65696 27402 65708
rect 27433 65705 27445 65708
rect 27479 65705 27491 65739
rect 27433 65699 27491 65705
rect 27798 65696 27804 65748
rect 27856 65736 27862 65748
rect 28721 65739 28779 65745
rect 28721 65736 28733 65739
rect 27856 65708 28733 65736
rect 27856 65696 27862 65708
rect 28721 65705 28733 65708
rect 28767 65705 28779 65739
rect 28721 65699 28779 65705
rect 20806 65668 20812 65680
rect 20548 65640 20812 65668
rect 17310 65600 17316 65612
rect 17271 65572 17316 65600
rect 17310 65560 17316 65572
rect 17368 65560 17374 65612
rect 17405 65603 17463 65609
rect 17405 65569 17417 65603
rect 17451 65600 17463 65603
rect 17494 65600 17500 65612
rect 17451 65572 17500 65600
rect 17451 65569 17463 65572
rect 17405 65563 17463 65569
rect 17494 65560 17500 65572
rect 17552 65560 17558 65612
rect 20548 65609 20576 65640
rect 20806 65628 20812 65640
rect 20864 65668 20870 65680
rect 21174 65668 21180 65680
rect 20864 65640 21180 65668
rect 20864 65628 20870 65640
rect 21174 65628 21180 65640
rect 21232 65628 21238 65680
rect 24302 65628 24308 65680
rect 24360 65668 24366 65680
rect 24360 65640 28120 65668
rect 24360 65628 24366 65640
rect 20533 65603 20591 65609
rect 20533 65569 20545 65603
rect 20579 65569 20591 65603
rect 20533 65563 20591 65569
rect 20714 65560 20720 65612
rect 20772 65600 20778 65612
rect 21361 65603 21419 65609
rect 21361 65600 21373 65603
rect 20772 65572 21373 65600
rect 20772 65560 20778 65572
rect 21361 65569 21373 65572
rect 21407 65569 21419 65603
rect 25222 65600 25228 65612
rect 25183 65572 25228 65600
rect 21361 65563 21419 65569
rect 25222 65560 25228 65572
rect 25280 65560 25286 65612
rect 1578 65532 1584 65544
rect 1539 65504 1584 65532
rect 1578 65492 1584 65504
rect 1636 65492 1642 65544
rect 12894 65532 12900 65544
rect 12855 65504 12900 65532
rect 12894 65492 12900 65504
rect 12952 65492 12958 65544
rect 15286 65532 15292 65544
rect 15247 65504 15292 65532
rect 15286 65492 15292 65504
rect 15344 65492 15350 65544
rect 17957 65535 18015 65541
rect 17957 65501 17969 65535
rect 18003 65532 18015 65535
rect 19245 65535 19303 65541
rect 19245 65532 19257 65535
rect 18003 65504 19257 65532
rect 18003 65501 18015 65504
rect 17957 65495 18015 65501
rect 19245 65501 19257 65504
rect 19291 65532 19303 65535
rect 19334 65532 19340 65544
rect 19291 65504 19340 65532
rect 19291 65501 19303 65504
rect 19245 65495 19303 65501
rect 19334 65492 19340 65504
rect 19392 65492 19398 65544
rect 24578 65492 24584 65544
rect 24636 65532 24642 65544
rect 24949 65535 25007 65541
rect 24949 65532 24961 65535
rect 24636 65504 24961 65532
rect 24636 65492 24642 65504
rect 24949 65501 24961 65504
rect 24995 65501 25007 65535
rect 24949 65495 25007 65501
rect 27614 65492 27620 65544
rect 27672 65532 27678 65544
rect 27709 65535 27767 65541
rect 27709 65532 27721 65535
rect 27672 65504 27721 65532
rect 27672 65492 27678 65504
rect 27709 65501 27721 65504
rect 27755 65501 27767 65535
rect 27709 65495 27767 65501
rect 27801 65535 27859 65541
rect 27801 65501 27813 65535
rect 27847 65501 27859 65535
rect 27801 65495 27859 65501
rect 20254 65464 20260 65476
rect 20215 65436 20260 65464
rect 20254 65424 20260 65436
rect 20312 65424 20318 65476
rect 21174 65424 21180 65476
rect 21232 65464 21238 65476
rect 21606 65467 21664 65473
rect 21606 65464 21618 65467
rect 21232 65436 21618 65464
rect 21232 65424 21238 65436
rect 21606 65433 21618 65436
rect 21652 65433 21664 65467
rect 27816 65464 27844 65495
rect 27890 65492 27896 65544
rect 27948 65532 27954 65544
rect 28092 65541 28120 65640
rect 29914 65628 29920 65680
rect 29972 65668 29978 65680
rect 31846 65668 31852 65680
rect 29972 65640 31852 65668
rect 29972 65628 29978 65640
rect 31846 65628 31852 65640
rect 31904 65628 31910 65680
rect 28077 65535 28135 65541
rect 27948 65504 27993 65532
rect 27948 65492 27954 65504
rect 28077 65501 28089 65535
rect 28123 65501 28135 65535
rect 28077 65495 28135 65501
rect 29825 65535 29883 65541
rect 29825 65501 29837 65535
rect 29871 65532 29883 65535
rect 29914 65532 29920 65544
rect 29871 65504 29920 65532
rect 29871 65501 29883 65504
rect 29825 65495 29883 65501
rect 29914 65492 29920 65504
rect 29972 65492 29978 65544
rect 28442 65464 28448 65476
rect 27816 65436 28448 65464
rect 21606 65427 21664 65433
rect 28442 65424 28448 65436
rect 28500 65424 28506 65476
rect 28629 65467 28687 65473
rect 28629 65433 28641 65467
rect 28675 65433 28687 65467
rect 28629 65427 28687 65433
rect 1397 65399 1455 65405
rect 1397 65365 1409 65399
rect 1443 65396 1455 65399
rect 11238 65396 11244 65408
rect 1443 65368 11244 65396
rect 1443 65365 1455 65368
rect 1397 65359 1455 65365
rect 11238 65356 11244 65368
rect 11296 65356 11302 65408
rect 17313 65399 17371 65405
rect 17313 65365 17325 65399
rect 17359 65396 17371 65399
rect 17586 65396 17592 65408
rect 17359 65368 17592 65396
rect 17359 65365 17371 65368
rect 17313 65359 17371 65365
rect 17586 65356 17592 65368
rect 17644 65356 17650 65408
rect 20438 65396 20444 65408
rect 20399 65368 20444 65396
rect 20438 65356 20444 65368
rect 20496 65356 20502 65408
rect 22738 65396 22744 65408
rect 22699 65368 22744 65396
rect 22738 65356 22744 65368
rect 22796 65356 22802 65408
rect 28350 65356 28356 65408
rect 28408 65396 28414 65408
rect 28644 65396 28672 65427
rect 28408 65368 28672 65396
rect 30009 65399 30067 65405
rect 28408 65356 28414 65368
rect 30009 65365 30021 65399
rect 30055 65396 30067 65399
rect 30558 65396 30564 65408
rect 30055 65368 30564 65396
rect 30055 65365 30067 65368
rect 30009 65359 30067 65365
rect 30558 65356 30564 65368
rect 30616 65356 30622 65408
rect 1104 65306 30820 65328
rect 1104 65254 10880 65306
rect 10932 65254 10944 65306
rect 10996 65254 11008 65306
rect 11060 65254 11072 65306
rect 11124 65254 11136 65306
rect 11188 65254 20811 65306
rect 20863 65254 20875 65306
rect 20927 65254 20939 65306
rect 20991 65254 21003 65306
rect 21055 65254 21067 65306
rect 21119 65254 30820 65306
rect 1104 65232 30820 65254
rect 13722 65152 13728 65204
rect 13780 65192 13786 65204
rect 13909 65195 13967 65201
rect 13909 65192 13921 65195
rect 13780 65164 13921 65192
rect 13780 65152 13786 65164
rect 13909 65161 13921 65164
rect 13955 65161 13967 65195
rect 13909 65155 13967 65161
rect 15286 65152 15292 65204
rect 15344 65192 15350 65204
rect 15455 65195 15513 65201
rect 15455 65192 15467 65195
rect 15344 65164 15467 65192
rect 15344 65152 15350 65164
rect 15455 65161 15467 65164
rect 15501 65161 15513 65195
rect 15455 65155 15513 65161
rect 15933 65195 15991 65201
rect 15933 65161 15945 65195
rect 15979 65192 15991 65195
rect 17586 65192 17592 65204
rect 15979 65164 17592 65192
rect 15979 65161 15991 65164
rect 15933 65155 15991 65161
rect 17586 65152 17592 65164
rect 17644 65152 17650 65204
rect 18690 65192 18696 65204
rect 18651 65164 18696 65192
rect 18690 65152 18696 65164
rect 18748 65152 18754 65204
rect 21266 65192 21272 65204
rect 19260 65164 21272 65192
rect 17494 65124 17500 65136
rect 17455 65096 17500 65124
rect 17494 65084 17500 65096
rect 17552 65084 17558 65136
rect 19260 65133 19288 65164
rect 21266 65152 21272 65164
rect 21324 65152 21330 65204
rect 21910 65152 21916 65204
rect 21968 65192 21974 65204
rect 23198 65192 23204 65204
rect 21968 65164 23204 65192
rect 21968 65152 21974 65164
rect 23198 65152 23204 65164
rect 23256 65152 23262 65204
rect 25961 65195 26019 65201
rect 25961 65161 25973 65195
rect 26007 65192 26019 65195
rect 27890 65192 27896 65204
rect 26007 65164 27896 65192
rect 26007 65161 26019 65164
rect 25961 65155 26019 65161
rect 27890 65152 27896 65164
rect 27948 65152 27954 65204
rect 19245 65127 19303 65133
rect 19245 65093 19257 65127
rect 19291 65093 19303 65127
rect 19245 65087 19303 65093
rect 19429 65127 19487 65133
rect 19429 65093 19441 65127
rect 19475 65124 19487 65127
rect 20438 65124 20444 65136
rect 19475 65096 20444 65124
rect 19475 65093 19487 65096
rect 19429 65087 19487 65093
rect 20438 65084 20444 65096
rect 20496 65084 20502 65136
rect 20533 65127 20591 65133
rect 20533 65093 20545 65127
rect 20579 65124 20591 65127
rect 20714 65124 20720 65136
rect 20579 65096 20720 65124
rect 20579 65093 20591 65096
rect 20533 65087 20591 65093
rect 20714 65084 20720 65096
rect 20772 65084 20778 65136
rect 21818 65084 21824 65136
rect 21876 65124 21882 65136
rect 22066 65127 22124 65133
rect 22066 65124 22078 65127
rect 21876 65096 22078 65124
rect 21876 65084 21882 65096
rect 22066 65093 22078 65096
rect 22112 65093 22124 65127
rect 22066 65087 22124 65093
rect 26160 65096 28028 65124
rect 12894 65056 12900 65068
rect 12855 65028 12900 65056
rect 12894 65016 12900 65028
rect 12952 65016 12958 65068
rect 13725 65059 13783 65065
rect 13725 65025 13737 65059
rect 13771 65056 13783 65059
rect 13998 65056 14004 65068
rect 13771 65028 14004 65056
rect 13771 65025 13783 65028
rect 13725 65019 13783 65025
rect 13998 65016 14004 65028
rect 14056 65016 14062 65068
rect 15562 65016 15568 65068
rect 15620 65056 15626 65068
rect 15749 65059 15807 65065
rect 15749 65056 15761 65059
rect 15620 65028 15761 65056
rect 15620 65016 15626 65028
rect 15749 65025 15761 65028
rect 15795 65025 15807 65059
rect 15749 65019 15807 65025
rect 17126 65016 17132 65068
rect 17184 65056 17190 65068
rect 17313 65059 17371 65065
rect 17313 65056 17325 65059
rect 17184 65028 17325 65056
rect 17184 65016 17190 65028
rect 17313 65025 17325 65028
rect 17359 65025 17371 65059
rect 17313 65019 17371 65025
rect 18509 65059 18567 65065
rect 18509 65025 18521 65059
rect 18555 65056 18567 65059
rect 18598 65056 18604 65068
rect 18555 65028 18604 65056
rect 18555 65025 18567 65028
rect 18509 65019 18567 65025
rect 18598 65016 18604 65028
rect 18656 65016 18662 65068
rect 20254 65056 20260 65068
rect 20215 65028 20260 65056
rect 20254 65016 20260 65028
rect 20312 65016 20318 65068
rect 21085 65059 21143 65065
rect 21085 65025 21097 65059
rect 21131 65025 21143 65059
rect 21085 65019 21143 65025
rect 14550 64948 14556 65000
rect 14608 64988 14614 65000
rect 16025 64991 16083 64997
rect 16025 64988 16037 64991
rect 14608 64960 16037 64988
rect 14608 64948 14614 64960
rect 16025 64957 16037 64960
rect 16071 64957 16083 64991
rect 16025 64951 16083 64957
rect 19981 64923 20039 64929
rect 19981 64889 19993 64923
rect 20027 64920 20039 64923
rect 21100 64920 21128 65019
rect 25498 65016 25504 65068
rect 25556 65056 25562 65068
rect 26160 65065 26188 65096
rect 26145 65059 26203 65065
rect 26145 65056 26157 65059
rect 25556 65028 26157 65056
rect 25556 65016 25562 65028
rect 26145 65025 26157 65028
rect 26191 65025 26203 65059
rect 26329 65059 26387 65065
rect 26329 65056 26341 65059
rect 26145 65019 26203 65025
rect 26252 65028 26341 65056
rect 21821 64991 21879 64997
rect 21821 64957 21833 64991
rect 21867 64957 21879 64991
rect 21821 64951 21879 64957
rect 20027 64892 21128 64920
rect 21269 64923 21327 64929
rect 20027 64889 20039 64892
rect 19981 64883 20039 64889
rect 21269 64889 21281 64923
rect 21315 64920 21327 64923
rect 21836 64920 21864 64951
rect 23474 64948 23480 65000
rect 23532 64988 23538 65000
rect 23750 64988 23756 65000
rect 23532 64960 23756 64988
rect 23532 64948 23538 64960
rect 23750 64948 23756 64960
rect 23808 64988 23814 65000
rect 26252 64988 26280 65028
rect 26329 65025 26341 65028
rect 26375 65025 26387 65059
rect 26329 65019 26387 65025
rect 26421 65059 26479 65065
rect 26421 65025 26433 65059
rect 26467 65025 26479 65059
rect 26421 65019 26479 65025
rect 26436 64988 26464 65019
rect 28000 64997 28028 65096
rect 28350 65016 28356 65068
rect 28408 65056 28414 65068
rect 29549 65059 29607 65065
rect 28408 65028 29316 65056
rect 28408 65016 28414 65028
rect 23808 64960 26280 64988
rect 26344 64960 26464 64988
rect 27985 64991 28043 64997
rect 23808 64948 23814 64960
rect 21315 64892 21864 64920
rect 21315 64889 21327 64892
rect 21269 64883 21327 64889
rect 26142 64880 26148 64932
rect 26200 64920 26206 64932
rect 26344 64920 26372 64960
rect 27985 64957 27997 64991
rect 28031 64988 28043 64991
rect 28074 64988 28080 65000
rect 28031 64960 28080 64988
rect 28031 64957 28043 64960
rect 27985 64951 28043 64957
rect 28074 64948 28080 64960
rect 28132 64948 28138 65000
rect 28261 64991 28319 64997
rect 28261 64957 28273 64991
rect 28307 64988 28319 64991
rect 28902 64988 28908 65000
rect 28307 64960 28908 64988
rect 28307 64957 28319 64960
rect 28261 64951 28319 64957
rect 28368 64932 28396 64960
rect 28902 64948 28908 64960
rect 28960 64948 28966 65000
rect 29288 64997 29316 65028
rect 29549 65025 29561 65059
rect 29595 65056 29607 65059
rect 30006 65056 30012 65068
rect 29595 65028 30012 65056
rect 29595 65025 29607 65028
rect 29549 65019 29607 65025
rect 30006 65016 30012 65028
rect 30064 65056 30070 65068
rect 30374 65056 30380 65068
rect 30064 65028 30380 65056
rect 30064 65016 30070 65028
rect 30374 65016 30380 65028
rect 30432 65016 30438 65068
rect 29273 64991 29331 64997
rect 29273 64957 29285 64991
rect 29319 64988 29331 64991
rect 29822 64988 29828 65000
rect 29319 64960 29828 64988
rect 29319 64957 29331 64960
rect 29273 64951 29331 64957
rect 29822 64948 29828 64960
rect 29880 64948 29886 65000
rect 26200 64892 26372 64920
rect 26200 64880 26206 64892
rect 28350 64880 28356 64932
rect 28408 64880 28414 64932
rect 12710 64852 12716 64864
rect 12671 64824 12716 64852
rect 12710 64812 12716 64824
rect 12768 64812 12774 64864
rect 15470 64812 15476 64864
rect 15528 64852 15534 64864
rect 21542 64852 21548 64864
rect 15528 64824 21548 64852
rect 15528 64812 15534 64824
rect 21542 64812 21548 64824
rect 21600 64812 21606 64864
rect 23382 64812 23388 64864
rect 23440 64852 23446 64864
rect 30742 64852 30748 64864
rect 23440 64824 30748 64852
rect 23440 64812 23446 64824
rect 30742 64812 30748 64824
rect 30800 64812 30806 64864
rect 1104 64762 30820 64784
rect 1104 64710 5915 64762
rect 5967 64710 5979 64762
rect 6031 64710 6043 64762
rect 6095 64710 6107 64762
rect 6159 64710 6171 64762
rect 6223 64710 15846 64762
rect 15898 64710 15910 64762
rect 15962 64710 15974 64762
rect 16026 64710 16038 64762
rect 16090 64710 16102 64762
rect 16154 64710 25776 64762
rect 25828 64710 25840 64762
rect 25892 64710 25904 64762
rect 25956 64710 25968 64762
rect 26020 64710 26032 64762
rect 26084 64710 30820 64762
rect 1104 64688 30820 64710
rect 19429 64651 19487 64657
rect 19429 64617 19441 64651
rect 19475 64648 19487 64651
rect 19978 64648 19984 64660
rect 19475 64620 19984 64648
rect 19475 64617 19487 64620
rect 19429 64611 19487 64617
rect 19978 64608 19984 64620
rect 20036 64608 20042 64660
rect 20070 64608 20076 64660
rect 20128 64648 20134 64660
rect 21174 64648 21180 64660
rect 20128 64620 20173 64648
rect 21135 64620 21180 64648
rect 20128 64608 20134 64620
rect 21174 64608 21180 64620
rect 21232 64608 21238 64660
rect 24854 64608 24860 64660
rect 24912 64648 24918 64660
rect 25222 64648 25228 64660
rect 24912 64620 25228 64648
rect 24912 64608 24918 64620
rect 25222 64608 25228 64620
rect 25280 64608 25286 64660
rect 26326 64608 26332 64660
rect 26384 64648 26390 64660
rect 27341 64651 27399 64657
rect 27341 64648 27353 64651
rect 26384 64620 27353 64648
rect 26384 64608 26390 64620
rect 27341 64617 27353 64620
rect 27387 64617 27399 64651
rect 31294 64648 31300 64660
rect 27341 64611 27399 64617
rect 28966 64620 31300 64648
rect 21634 64540 21640 64592
rect 21692 64580 21698 64592
rect 22370 64580 22376 64592
rect 21692 64552 22376 64580
rect 21692 64540 21698 64552
rect 22370 64540 22376 64552
rect 22428 64540 22434 64592
rect 28966 64580 28994 64620
rect 31294 64608 31300 64620
rect 31352 64608 31358 64660
rect 26804 64552 28994 64580
rect 20346 64472 20352 64524
rect 20404 64512 20410 64524
rect 20404 64484 21864 64512
rect 20404 64472 20410 64484
rect 1578 64444 1584 64456
rect 1539 64416 1584 64444
rect 1578 64404 1584 64416
rect 1636 64404 1642 64456
rect 11238 64404 11244 64456
rect 11296 64444 11302 64456
rect 12897 64447 12955 64453
rect 12897 64444 12909 64447
rect 11296 64416 12909 64444
rect 11296 64404 11302 64416
rect 12897 64413 12909 64416
rect 12943 64413 12955 64447
rect 12897 64407 12955 64413
rect 19245 64447 19303 64453
rect 19245 64413 19257 64447
rect 19291 64444 19303 64447
rect 19334 64444 19340 64456
rect 19291 64416 19340 64444
rect 19291 64413 19303 64416
rect 19245 64407 19303 64413
rect 19334 64404 19340 64416
rect 19392 64404 19398 64456
rect 21453 64447 21511 64453
rect 21453 64413 21465 64447
rect 21499 64413 21511 64447
rect 21453 64407 21511 64413
rect 21545 64447 21603 64453
rect 21545 64413 21557 64447
rect 21591 64413 21603 64447
rect 21545 64407 21603 64413
rect 12710 64376 12716 64388
rect 12671 64348 12716 64376
rect 12710 64336 12716 64348
rect 12768 64336 12774 64388
rect 19981 64379 20039 64385
rect 19981 64345 19993 64379
rect 20027 64376 20039 64379
rect 20530 64376 20536 64388
rect 20027 64348 20536 64376
rect 20027 64345 20039 64348
rect 19981 64339 20039 64345
rect 20530 64336 20536 64348
rect 20588 64336 20594 64388
rect 1397 64311 1455 64317
rect 1397 64277 1409 64311
rect 1443 64308 1455 64311
rect 12158 64308 12164 64320
rect 1443 64280 12164 64308
rect 1443 64277 1455 64280
rect 1397 64271 1455 64277
rect 12158 64268 12164 64280
rect 12216 64268 12222 64320
rect 13081 64311 13139 64317
rect 13081 64277 13093 64311
rect 13127 64308 13139 64311
rect 15102 64308 15108 64320
rect 13127 64280 15108 64308
rect 13127 64277 13139 64280
rect 13081 64271 13139 64277
rect 15102 64268 15108 64280
rect 15160 64268 15166 64320
rect 21468 64308 21496 64407
rect 21560 64376 21588 64407
rect 21634 64404 21640 64456
rect 21692 64444 21698 64456
rect 21836 64453 21864 64484
rect 24394 64472 24400 64524
rect 24452 64512 24458 64524
rect 26804 64512 26832 64552
rect 24452 64484 26924 64512
rect 24452 64472 24458 64484
rect 21821 64447 21879 64453
rect 21692 64416 21737 64444
rect 21692 64404 21698 64416
rect 21821 64413 21833 64447
rect 21867 64413 21879 64447
rect 22738 64444 22744 64456
rect 21821 64407 21879 64413
rect 22066 64416 22744 64444
rect 21910 64376 21916 64388
rect 21560 64348 21916 64376
rect 21910 64336 21916 64348
rect 21968 64336 21974 64388
rect 22066 64308 22094 64416
rect 22738 64404 22744 64416
rect 22796 64444 22802 64456
rect 23385 64447 23443 64453
rect 23385 64444 23397 64447
rect 22796 64416 23397 64444
rect 22796 64404 22802 64416
rect 23385 64413 23397 64416
rect 23431 64413 23443 64447
rect 23385 64407 23443 64413
rect 23474 64404 23480 64456
rect 23532 64444 23538 64456
rect 23569 64447 23627 64453
rect 23569 64444 23581 64447
rect 23532 64416 23581 64444
rect 23532 64404 23538 64416
rect 23569 64413 23581 64416
rect 23615 64413 23627 64447
rect 23569 64407 23627 64413
rect 24857 64447 24915 64453
rect 24857 64413 24869 64447
rect 24903 64444 24915 64447
rect 24946 64444 24952 64456
rect 24903 64416 24952 64444
rect 24903 64413 24915 64416
rect 24857 64407 24915 64413
rect 24946 64404 24952 64416
rect 25004 64404 25010 64456
rect 25130 64444 25136 64456
rect 25091 64416 25136 64444
rect 25130 64404 25136 64416
rect 25188 64404 25194 64456
rect 25498 64404 25504 64456
rect 25556 64444 25562 64456
rect 25869 64447 25927 64453
rect 25869 64444 25881 64447
rect 25556 64416 25881 64444
rect 25556 64404 25562 64416
rect 25869 64413 25881 64416
rect 25915 64413 25927 64447
rect 26142 64444 26148 64456
rect 26103 64416 26148 64444
rect 25869 64407 25927 64413
rect 26142 64404 26148 64416
rect 26200 64404 26206 64456
rect 26326 64404 26332 64456
rect 26384 64444 26390 64456
rect 26896 64453 26924 64484
rect 27062 64472 27068 64524
rect 27120 64512 27126 64524
rect 27614 64512 27620 64524
rect 27120 64484 27620 64512
rect 27120 64472 27126 64484
rect 27614 64472 27620 64484
rect 27672 64512 27678 64524
rect 28077 64515 28135 64521
rect 28077 64512 28089 64515
rect 27672 64484 28089 64512
rect 27672 64472 27678 64484
rect 28077 64481 28089 64484
rect 28123 64481 28135 64515
rect 28077 64475 28135 64481
rect 26605 64447 26663 64453
rect 26605 64444 26617 64447
rect 26384 64416 26617 64444
rect 26384 64404 26390 64416
rect 26605 64413 26617 64416
rect 26651 64413 26663 64447
rect 26605 64407 26663 64413
rect 26789 64447 26847 64453
rect 26789 64413 26801 64447
rect 26835 64413 26847 64447
rect 26789 64407 26847 64413
rect 26881 64447 26939 64453
rect 26881 64413 26893 64447
rect 26927 64413 26939 64447
rect 26881 64407 26939 64413
rect 24486 64336 24492 64388
rect 24544 64376 24550 64388
rect 24762 64376 24768 64388
rect 24544 64348 24768 64376
rect 24544 64336 24550 64348
rect 24762 64336 24768 64348
rect 24820 64376 24826 64388
rect 25041 64379 25099 64385
rect 25041 64376 25053 64379
rect 24820 64348 25053 64376
rect 24820 64336 24826 64348
rect 25041 64345 25053 64348
rect 25087 64345 25099 64379
rect 25041 64339 25099 64345
rect 25685 64379 25743 64385
rect 25685 64345 25697 64379
rect 25731 64376 25743 64379
rect 26510 64376 26516 64388
rect 25731 64348 26516 64376
rect 25731 64345 25743 64348
rect 25685 64339 25743 64345
rect 26510 64336 26516 64348
rect 26568 64336 26574 64388
rect 21468 64280 22094 64308
rect 23753 64311 23811 64317
rect 23753 64277 23765 64311
rect 23799 64308 23811 64311
rect 24118 64308 24124 64320
rect 23799 64280 24124 64308
rect 23799 64277 23811 64280
rect 23753 64271 23811 64277
rect 24118 64268 24124 64280
rect 24176 64268 24182 64320
rect 24670 64308 24676 64320
rect 24631 64280 24676 64308
rect 24670 64268 24676 64280
rect 24728 64268 24734 64320
rect 25222 64268 25228 64320
rect 25280 64308 25286 64320
rect 26053 64311 26111 64317
rect 26053 64308 26065 64311
rect 25280 64280 26065 64308
rect 25280 64268 25286 64280
rect 26053 64277 26065 64280
rect 26099 64277 26111 64311
rect 26804 64308 26832 64407
rect 26970 64404 26976 64456
rect 27028 64444 27034 64456
rect 27157 64447 27215 64453
rect 27028 64416 27073 64444
rect 27028 64404 27034 64416
rect 27157 64413 27169 64447
rect 27203 64444 27215 64447
rect 27798 64444 27804 64456
rect 27203 64416 27804 64444
rect 27203 64413 27215 64416
rect 27157 64407 27215 64413
rect 27798 64404 27804 64416
rect 27856 64404 27862 64456
rect 27890 64404 27896 64456
rect 27948 64444 27954 64456
rect 31110 64444 31116 64456
rect 27948 64416 31116 64444
rect 27948 64404 27954 64416
rect 31110 64404 31116 64416
rect 31168 64404 31174 64456
rect 28902 64336 28908 64388
rect 28960 64376 28966 64388
rect 28960 64348 29224 64376
rect 28960 64336 28966 64348
rect 28350 64308 28356 64320
rect 26804 64280 28356 64308
rect 26053 64271 26111 64277
rect 28350 64268 28356 64280
rect 28408 64268 28414 64320
rect 28626 64268 28632 64320
rect 28684 64308 28690 64320
rect 29086 64308 29092 64320
rect 28684 64280 29092 64308
rect 28684 64268 28690 64280
rect 29086 64268 29092 64280
rect 29144 64268 29150 64320
rect 29196 64308 29224 64348
rect 29822 64336 29828 64388
rect 29880 64376 29886 64388
rect 29917 64379 29975 64385
rect 29917 64376 29929 64379
rect 29880 64348 29929 64376
rect 29880 64336 29886 64348
rect 29917 64345 29929 64348
rect 29963 64376 29975 64379
rect 30374 64376 30380 64388
rect 29963 64348 30380 64376
rect 29963 64345 29975 64348
rect 29917 64339 29975 64345
rect 30374 64336 30380 64348
rect 30432 64336 30438 64388
rect 30009 64311 30067 64317
rect 30009 64308 30021 64311
rect 29196 64280 30021 64308
rect 30009 64277 30021 64280
rect 30055 64277 30067 64311
rect 30009 64271 30067 64277
rect 1104 64218 30820 64240
rect 1104 64166 10880 64218
rect 10932 64166 10944 64218
rect 10996 64166 11008 64218
rect 11060 64166 11072 64218
rect 11124 64166 11136 64218
rect 11188 64166 20811 64218
rect 20863 64166 20875 64218
rect 20927 64166 20939 64218
rect 20991 64166 21003 64218
rect 21055 64166 21067 64218
rect 21119 64166 30820 64218
rect 1104 64144 30820 64166
rect 11330 64064 11336 64116
rect 11388 64104 11394 64116
rect 20622 64104 20628 64116
rect 11388 64076 12434 64104
rect 11388 64064 11394 64076
rect 12158 64036 12164 64048
rect 12119 64008 12164 64036
rect 12158 63996 12164 64008
rect 12216 63996 12222 64048
rect 12406 64036 12434 64076
rect 19812 64076 20628 64104
rect 12989 64039 13047 64045
rect 12989 64036 13001 64039
rect 12406 64008 13001 64036
rect 12989 64005 13001 64008
rect 13035 64005 13047 64039
rect 12989 63999 13047 64005
rect 14461 64039 14519 64045
rect 14461 64005 14473 64039
rect 14507 64036 14519 64039
rect 14642 64036 14648 64048
rect 14507 64008 14648 64036
rect 14507 64005 14519 64008
rect 14461 63999 14519 64005
rect 14642 63996 14648 64008
rect 14700 63996 14706 64048
rect 19812 64045 19840 64076
rect 20622 64064 20628 64076
rect 20680 64064 20686 64116
rect 25498 64064 25504 64116
rect 25556 64104 25562 64116
rect 25682 64104 25688 64116
rect 25556 64076 25688 64104
rect 25556 64064 25562 64076
rect 25682 64064 25688 64076
rect 25740 64064 25746 64116
rect 26786 64064 26792 64116
rect 26844 64104 26850 64116
rect 26973 64107 27031 64113
rect 26973 64104 26985 64107
rect 26844 64076 26985 64104
rect 26844 64064 26850 64076
rect 26973 64073 26985 64076
rect 27019 64073 27031 64107
rect 26973 64067 27031 64073
rect 27264 64076 27660 64104
rect 19797 64039 19855 64045
rect 19797 64005 19809 64039
rect 19843 64005 19855 64039
rect 19797 63999 19855 64005
rect 19981 64039 20039 64045
rect 19981 64005 19993 64039
rect 20027 64036 20039 64039
rect 20254 64036 20260 64048
rect 20027 64008 20260 64036
rect 20027 64005 20039 64008
rect 19981 63999 20039 64005
rect 20254 63996 20260 64008
rect 20312 63996 20318 64048
rect 20714 64036 20720 64048
rect 20675 64008 20720 64036
rect 20714 63996 20720 64008
rect 20772 63996 20778 64048
rect 24670 63996 24676 64048
rect 24728 64036 24734 64048
rect 27264 64036 27292 64076
rect 27522 64036 27528 64048
rect 24728 64008 27292 64036
rect 27377 64008 27528 64036
rect 24728 63996 24734 64008
rect 1578 63968 1584 63980
rect 1539 63940 1584 63968
rect 1578 63928 1584 63940
rect 1636 63928 1642 63980
rect 11977 63971 12035 63977
rect 11977 63937 11989 63971
rect 12023 63968 12035 63971
rect 12710 63968 12716 63980
rect 12023 63940 12716 63968
rect 12023 63937 12035 63940
rect 11977 63931 12035 63937
rect 12710 63928 12716 63940
rect 12768 63968 12774 63980
rect 12805 63971 12863 63977
rect 12805 63968 12817 63971
rect 12768 63940 12817 63968
rect 12768 63928 12774 63940
rect 12805 63937 12817 63940
rect 12851 63937 12863 63971
rect 12805 63931 12863 63937
rect 14277 63971 14335 63977
rect 14277 63937 14289 63971
rect 14323 63968 14335 63971
rect 15562 63968 15568 63980
rect 14323 63940 15568 63968
rect 14323 63937 14335 63940
rect 14277 63931 14335 63937
rect 15562 63928 15568 63940
rect 15620 63928 15626 63980
rect 17126 63968 17132 63980
rect 17087 63940 17132 63968
rect 17126 63928 17132 63940
rect 17184 63928 17190 63980
rect 20530 63968 20536 63980
rect 20443 63940 20536 63968
rect 20530 63928 20536 63940
rect 20588 63968 20594 63980
rect 22922 63968 22928 63980
rect 20588 63940 22928 63968
rect 20588 63928 20594 63940
rect 22922 63928 22928 63940
rect 22980 63928 22986 63980
rect 23198 63928 23204 63980
rect 23256 63968 23262 63980
rect 23385 63971 23443 63977
rect 23385 63968 23397 63971
rect 23256 63940 23397 63968
rect 23256 63928 23262 63940
rect 23385 63937 23397 63940
rect 23431 63937 23443 63971
rect 23385 63931 23443 63937
rect 23474 63928 23480 63980
rect 23532 63968 23538 63980
rect 23569 63971 23627 63977
rect 23569 63968 23581 63971
rect 23532 63940 23581 63968
rect 23532 63928 23538 63940
rect 23569 63937 23581 63940
rect 23615 63937 23627 63971
rect 23569 63931 23627 63937
rect 25130 63928 25136 63980
rect 25188 63968 25194 63980
rect 25225 63971 25283 63977
rect 25225 63968 25237 63971
rect 25188 63940 25237 63968
rect 25188 63928 25194 63940
rect 25225 63937 25237 63940
rect 25271 63937 25283 63971
rect 25225 63931 25283 63937
rect 27062 63928 27068 63980
rect 27120 63968 27126 63980
rect 27377 63977 27405 64008
rect 27522 63996 27528 64008
rect 27580 63996 27586 64048
rect 27632 63977 27660 64076
rect 27706 64064 27712 64116
rect 27764 64104 27770 64116
rect 28905 64107 28963 64113
rect 28905 64104 28917 64107
rect 27764 64076 28917 64104
rect 27764 64064 27770 64076
rect 28905 64073 28917 64076
rect 28951 64073 28963 64107
rect 28905 64067 28963 64073
rect 29454 64064 29460 64116
rect 29512 64104 29518 64116
rect 30101 64107 30159 64113
rect 30101 64104 30113 64107
rect 29512 64076 30113 64104
rect 29512 64064 29518 64076
rect 30101 64073 30113 64076
rect 30147 64073 30159 64107
rect 30101 64067 30159 64073
rect 29086 64036 29092 64048
rect 28736 64008 29092 64036
rect 27249 63971 27307 63977
rect 27249 63968 27261 63971
rect 27120 63940 27261 63968
rect 27120 63928 27126 63940
rect 27249 63937 27261 63940
rect 27295 63937 27307 63971
rect 27249 63931 27307 63937
rect 27338 63971 27405 63977
rect 27338 63937 27350 63971
rect 27384 63940 27405 63971
rect 27433 63971 27491 63977
rect 27384 63937 27396 63940
rect 27338 63931 27396 63937
rect 27433 63937 27445 63971
rect 27479 63937 27491 63971
rect 27433 63931 27491 63937
rect 27617 63971 27675 63977
rect 27617 63937 27629 63971
rect 27663 63937 27675 63971
rect 28166 63968 28172 63980
rect 28127 63940 28172 63968
rect 27617 63931 27675 63937
rect 12345 63903 12403 63909
rect 12345 63869 12357 63903
rect 12391 63900 12403 63903
rect 14550 63900 14556 63912
rect 12391 63872 14412 63900
rect 14511 63872 14556 63900
rect 12391 63869 12403 63872
rect 12345 63863 12403 63869
rect 13998 63832 14004 63844
rect 13959 63804 14004 63832
rect 13998 63792 14004 63804
rect 14056 63792 14062 63844
rect 14384 63832 14412 63872
rect 14550 63860 14556 63872
rect 14608 63900 14614 63912
rect 17313 63903 17371 63909
rect 17313 63900 17325 63903
rect 14608 63872 17325 63900
rect 14608 63860 14614 63872
rect 17313 63869 17325 63872
rect 17359 63869 17371 63903
rect 17313 63863 17371 63869
rect 24026 63860 24032 63912
rect 24084 63900 24090 63912
rect 24949 63903 25007 63909
rect 24949 63900 24961 63903
rect 24084 63872 24961 63900
rect 24084 63860 24090 63872
rect 24949 63869 24961 63872
rect 24995 63900 25007 63903
rect 25406 63900 25412 63912
rect 24995 63872 25412 63900
rect 24995 63869 25007 63872
rect 24949 63863 25007 63869
rect 25406 63860 25412 63872
rect 25464 63860 25470 63912
rect 25682 63860 25688 63912
rect 25740 63900 25746 63912
rect 27448 63900 27476 63931
rect 28166 63928 28172 63940
rect 28224 63928 28230 63980
rect 28350 63968 28356 63980
rect 28311 63940 28356 63968
rect 28350 63928 28356 63940
rect 28408 63968 28414 63980
rect 28736 63977 28764 64008
rect 29086 63996 29092 64008
rect 29144 64036 29150 64048
rect 29144 64008 29960 64036
rect 29144 63996 29150 64008
rect 28721 63971 28779 63977
rect 28408 63940 28672 63968
rect 28408 63928 28414 63940
rect 25740 63872 27476 63900
rect 25740 63860 25746 63872
rect 28074 63860 28080 63912
rect 28132 63900 28138 63912
rect 28445 63903 28503 63909
rect 28445 63900 28457 63903
rect 28132 63872 28457 63900
rect 28132 63860 28138 63872
rect 28445 63869 28457 63872
rect 28491 63869 28503 63903
rect 28445 63863 28503 63869
rect 28537 63903 28595 63909
rect 28537 63869 28549 63903
rect 28583 63869 28595 63903
rect 28644 63900 28672 63940
rect 28721 63937 28733 63971
rect 28767 63937 28779 63971
rect 28721 63931 28779 63937
rect 29365 63971 29423 63977
rect 29365 63937 29377 63971
rect 29411 63968 29423 63971
rect 29454 63968 29460 63980
rect 29411 63940 29460 63968
rect 29411 63937 29423 63940
rect 29365 63931 29423 63937
rect 29454 63928 29460 63940
rect 29512 63928 29518 63980
rect 29932 63977 29960 64008
rect 29549 63971 29607 63977
rect 29549 63937 29561 63971
rect 29595 63937 29607 63971
rect 29549 63931 29607 63937
rect 29641 63971 29699 63977
rect 29641 63937 29653 63971
rect 29687 63968 29699 63971
rect 29917 63971 29975 63977
rect 29687 63940 29868 63968
rect 29687 63937 29699 63940
rect 29641 63931 29699 63937
rect 29564 63900 29592 63931
rect 28644 63872 29592 63900
rect 29733 63903 29791 63909
rect 28537 63863 28595 63869
rect 29733 63869 29745 63903
rect 29779 63869 29791 63903
rect 29840 63900 29868 63940
rect 29917 63937 29929 63971
rect 29963 63968 29975 63971
rect 30006 63968 30012 63980
rect 29963 63940 30012 63968
rect 29963 63937 29975 63940
rect 29917 63931 29975 63937
rect 30006 63928 30012 63940
rect 30064 63928 30070 63980
rect 30742 63900 30748 63912
rect 29840 63872 30748 63900
rect 29733 63863 29791 63869
rect 17954 63832 17960 63844
rect 14384 63804 17960 63832
rect 17954 63792 17960 63804
rect 18012 63792 18018 63844
rect 23753 63835 23811 63841
rect 23753 63801 23765 63835
rect 23799 63832 23811 63835
rect 27706 63832 27712 63844
rect 23799 63804 27712 63832
rect 23799 63801 23811 63804
rect 23753 63795 23811 63801
rect 27706 63792 27712 63804
rect 27764 63792 27770 63844
rect 1397 63767 1455 63773
rect 1397 63733 1409 63767
rect 1443 63764 1455 63767
rect 11330 63764 11336 63776
rect 1443 63736 11336 63764
rect 1443 63733 1455 63736
rect 1397 63727 1455 63733
rect 11330 63724 11336 63736
rect 11388 63724 11394 63776
rect 13173 63767 13231 63773
rect 13173 63733 13185 63767
rect 13219 63764 13231 63767
rect 13906 63764 13912 63776
rect 13219 63736 13912 63764
rect 13219 63733 13231 63736
rect 13173 63727 13231 63733
rect 13906 63724 13912 63736
rect 13964 63724 13970 63776
rect 24118 63724 24124 63776
rect 24176 63764 24182 63776
rect 28092 63764 28120 63860
rect 28258 63792 28264 63844
rect 28316 63832 28322 63844
rect 28552 63832 28580 63863
rect 28316 63804 28580 63832
rect 28316 63792 28322 63804
rect 28810 63792 28816 63844
rect 28868 63832 28874 63844
rect 29748 63832 29776 63863
rect 30742 63860 30748 63872
rect 30800 63900 30806 63912
rect 31662 63900 31668 63912
rect 30800 63872 31668 63900
rect 30800 63860 30806 63872
rect 31662 63860 31668 63872
rect 31720 63860 31726 63912
rect 28868 63804 29776 63832
rect 28868 63792 28874 63804
rect 24176 63736 28120 63764
rect 24176 63724 24182 63736
rect 1104 63674 30820 63696
rect 1104 63622 5915 63674
rect 5967 63622 5979 63674
rect 6031 63622 6043 63674
rect 6095 63622 6107 63674
rect 6159 63622 6171 63674
rect 6223 63622 15846 63674
rect 15898 63622 15910 63674
rect 15962 63622 15974 63674
rect 16026 63622 16038 63674
rect 16090 63622 16102 63674
rect 16154 63622 25776 63674
rect 25828 63622 25840 63674
rect 25892 63622 25904 63674
rect 25956 63622 25968 63674
rect 26020 63622 26032 63674
rect 26084 63622 30820 63674
rect 1104 63600 30820 63622
rect 23382 63520 23388 63572
rect 23440 63560 23446 63572
rect 23658 63560 23664 63572
rect 23440 63532 23664 63560
rect 23440 63520 23446 63532
rect 23658 63520 23664 63532
rect 23716 63520 23722 63572
rect 27706 63520 27712 63572
rect 27764 63560 27770 63572
rect 27764 63532 28396 63560
rect 27764 63520 27770 63532
rect 13814 63452 13820 63504
rect 13872 63492 13878 63504
rect 14185 63495 14243 63501
rect 14185 63492 14197 63495
rect 13872 63464 14197 63492
rect 13872 63452 13878 63464
rect 14185 63461 14197 63464
rect 14231 63461 14243 63495
rect 15562 63492 15568 63504
rect 14185 63455 14243 63461
rect 14660 63464 15568 63492
rect 14660 63433 14688 63464
rect 15562 63452 15568 63464
rect 15620 63452 15626 63504
rect 16761 63495 16819 63501
rect 16761 63461 16773 63495
rect 16807 63492 16819 63495
rect 17770 63492 17776 63504
rect 16807 63464 17776 63492
rect 16807 63461 16819 63464
rect 16761 63455 16819 63461
rect 17770 63452 17776 63464
rect 17828 63452 17834 63504
rect 19889 63495 19947 63501
rect 19889 63461 19901 63495
rect 19935 63492 19947 63495
rect 20346 63492 20352 63504
rect 19935 63464 20352 63492
rect 19935 63461 19947 63464
rect 19889 63455 19947 63461
rect 20346 63452 20352 63464
rect 20404 63452 20410 63504
rect 23293 63495 23351 63501
rect 23293 63461 23305 63495
rect 23339 63492 23351 63495
rect 23566 63492 23572 63504
rect 23339 63464 23572 63492
rect 23339 63461 23351 63464
rect 23293 63455 23351 63461
rect 23566 63452 23572 63464
rect 23624 63452 23630 63504
rect 27525 63495 27583 63501
rect 27525 63461 27537 63495
rect 27571 63492 27583 63495
rect 28074 63492 28080 63504
rect 27571 63464 28080 63492
rect 27571 63461 27583 63464
rect 27525 63455 27583 63461
rect 28074 63452 28080 63464
rect 28132 63452 28138 63504
rect 28258 63452 28264 63504
rect 28316 63452 28322 63504
rect 13173 63427 13231 63433
rect 13173 63393 13185 63427
rect 13219 63424 13231 63427
rect 14645 63427 14703 63433
rect 13219 63396 14596 63424
rect 13219 63393 13231 63396
rect 13173 63387 13231 63393
rect 1578 63356 1584 63368
rect 1539 63328 1584 63356
rect 1578 63316 1584 63328
rect 1636 63316 1642 63368
rect 12989 63359 13047 63365
rect 12989 63356 13001 63359
rect 12406 63328 13001 63356
rect 11422 63248 11428 63300
rect 11480 63288 11486 63300
rect 12406 63288 12434 63328
rect 12989 63325 13001 63328
rect 13035 63325 13047 63359
rect 12989 63319 13047 63325
rect 13814 63316 13820 63368
rect 13872 63356 13878 63368
rect 14182 63356 14188 63368
rect 13872 63328 14188 63356
rect 13872 63316 13878 63328
rect 14182 63316 14188 63328
rect 14240 63316 14246 63368
rect 14568 63356 14596 63396
rect 14645 63393 14657 63427
rect 14691 63393 14703 63427
rect 20254 63424 20260 63436
rect 20215 63396 20260 63424
rect 14645 63387 14703 63393
rect 20254 63384 20260 63396
rect 20312 63384 20318 63436
rect 20441 63427 20499 63433
rect 20441 63393 20453 63427
rect 20487 63424 20499 63427
rect 20714 63424 20720 63436
rect 20487 63396 20720 63424
rect 20487 63393 20499 63396
rect 20441 63387 20499 63393
rect 20714 63384 20720 63396
rect 20772 63384 20778 63436
rect 23658 63384 23664 63436
rect 23716 63424 23722 63436
rect 24578 63424 24584 63436
rect 23716 63396 24584 63424
rect 23716 63384 23722 63396
rect 24578 63384 24584 63396
rect 24636 63384 24642 63436
rect 28276 63424 28304 63452
rect 27816 63396 28304 63424
rect 28368 63424 28396 63532
rect 28534 63520 28540 63572
rect 28592 63520 28598 63572
rect 28552 63492 28580 63520
rect 28997 63495 29055 63501
rect 28997 63492 29009 63495
rect 28552 63464 29009 63492
rect 28997 63461 29009 63464
rect 29043 63461 29055 63495
rect 28997 63455 29055 63461
rect 28534 63433 28540 63436
rect 28531 63424 28540 63433
rect 28368 63396 28540 63424
rect 15562 63356 15568 63368
rect 14568 63328 15568 63356
rect 15562 63316 15568 63328
rect 15620 63316 15626 63368
rect 23477 63359 23535 63365
rect 23477 63325 23489 63359
rect 23523 63356 23535 63359
rect 23842 63356 23848 63368
rect 23523 63328 23848 63356
rect 23523 63325 23535 63328
rect 23477 63319 23535 63325
rect 23842 63316 23848 63328
rect 23900 63316 23906 63368
rect 24857 63359 24915 63365
rect 24857 63325 24869 63359
rect 24903 63356 24915 63359
rect 24946 63356 24952 63368
rect 24903 63328 24952 63356
rect 24903 63325 24915 63328
rect 24857 63319 24915 63325
rect 24946 63316 24952 63328
rect 25004 63316 25010 63368
rect 25406 63316 25412 63368
rect 25464 63356 25470 63368
rect 25961 63359 26019 63365
rect 25961 63356 25973 63359
rect 25464 63328 25973 63356
rect 25464 63316 25470 63328
rect 25961 63325 25973 63328
rect 26007 63325 26019 63359
rect 25961 63319 26019 63325
rect 26789 63359 26847 63365
rect 26789 63325 26801 63359
rect 26835 63325 26847 63359
rect 26789 63319 26847 63325
rect 27341 63359 27399 63365
rect 27341 63325 27353 63359
rect 27387 63356 27399 63359
rect 27706 63356 27712 63368
rect 27387 63328 27712 63356
rect 27387 63325 27399 63328
rect 27341 63319 27399 63325
rect 11480 63260 12434 63288
rect 11480 63248 11486 63260
rect 12710 63248 12716 63300
rect 12768 63288 12774 63300
rect 12805 63291 12863 63297
rect 12805 63288 12817 63291
rect 12768 63260 12817 63288
rect 12768 63248 12774 63260
rect 12805 63257 12817 63260
rect 12851 63257 12863 63291
rect 12805 63251 12863 63257
rect 14550 63248 14556 63300
rect 14608 63288 14614 63300
rect 14737 63291 14795 63297
rect 14737 63288 14749 63291
rect 14608 63260 14749 63288
rect 14608 63248 14614 63260
rect 14737 63257 14749 63260
rect 14783 63257 14795 63291
rect 15378 63288 15384 63300
rect 15339 63260 15384 63288
rect 14737 63251 14795 63257
rect 15378 63248 15384 63260
rect 15436 63248 15442 63300
rect 16574 63288 16580 63300
rect 16535 63260 16580 63288
rect 16574 63248 16580 63260
rect 16632 63248 16638 63300
rect 23934 63288 23940 63300
rect 16684 63260 23940 63288
rect 1397 63223 1455 63229
rect 1397 63189 1409 63223
rect 1443 63220 1455 63223
rect 11238 63220 11244 63232
rect 1443 63192 11244 63220
rect 1443 63189 1455 63192
rect 1397 63183 1455 63189
rect 11238 63180 11244 63192
rect 11296 63180 11302 63232
rect 14642 63220 14648 63232
rect 14603 63192 14648 63220
rect 14642 63180 14648 63192
rect 14700 63180 14706 63232
rect 15010 63180 15016 63232
rect 15068 63220 15074 63232
rect 16684 63220 16712 63260
rect 23934 63248 23940 63260
rect 23992 63288 23998 63300
rect 24578 63288 24584 63300
rect 23992 63260 24584 63288
rect 23992 63248 23998 63260
rect 24578 63248 24584 63260
rect 24636 63248 24642 63300
rect 26804 63288 26832 63319
rect 27706 63316 27712 63328
rect 27764 63316 27770 63368
rect 27614 63288 27620 63300
rect 26804 63260 27620 63288
rect 27614 63248 27620 63260
rect 27672 63248 27678 63300
rect 15068 63192 16712 63220
rect 20349 63223 20407 63229
rect 15068 63180 15074 63192
rect 20349 63189 20361 63223
rect 20395 63220 20407 63223
rect 21266 63220 21272 63232
rect 20395 63192 21272 63220
rect 20395 63189 20407 63192
rect 20349 63183 20407 63189
rect 21266 63180 21272 63192
rect 21324 63180 21330 63232
rect 25406 63180 25412 63232
rect 25464 63220 25470 63232
rect 26053 63223 26111 63229
rect 26053 63220 26065 63223
rect 25464 63192 26065 63220
rect 25464 63180 25470 63192
rect 26053 63189 26065 63192
rect 26099 63220 26111 63223
rect 26142 63220 26148 63232
rect 26099 63192 26148 63220
rect 26099 63189 26111 63192
rect 26053 63183 26111 63189
rect 26142 63180 26148 63192
rect 26200 63180 26206 63232
rect 26786 63180 26792 63232
rect 26844 63220 26850 63232
rect 26973 63223 27031 63229
rect 26973 63220 26985 63223
rect 26844 63192 26985 63220
rect 26844 63180 26850 63192
rect 26973 63189 26985 63192
rect 27019 63220 27031 63223
rect 27816 63220 27844 63396
rect 28531 63387 28540 63396
rect 28534 63384 28540 63387
rect 28592 63384 28598 63436
rect 30558 63424 30564 63436
rect 28644 63396 30564 63424
rect 28258 63356 28264 63368
rect 28219 63328 28264 63356
rect 28258 63316 28264 63328
rect 28316 63316 28322 63368
rect 28350 63316 28356 63368
rect 28408 63356 28414 63368
rect 28644 63365 28672 63396
rect 30558 63384 30564 63396
rect 30616 63384 30622 63436
rect 28445 63359 28503 63365
rect 28445 63356 28457 63359
rect 28408 63328 28457 63356
rect 28408 63316 28414 63328
rect 28445 63325 28457 63328
rect 28491 63325 28503 63359
rect 28445 63319 28503 63325
rect 28629 63359 28687 63365
rect 28629 63325 28641 63359
rect 28675 63325 28687 63359
rect 28629 63319 28687 63325
rect 28813 63359 28871 63365
rect 28813 63325 28825 63359
rect 28859 63358 28871 63359
rect 28859 63356 28948 63358
rect 29086 63356 29092 63368
rect 28859 63330 29092 63356
rect 28859 63325 28871 63330
rect 28920 63328 29092 63330
rect 28813 63319 28871 63325
rect 27985 63291 28043 63297
rect 27985 63257 27997 63291
rect 28031 63288 28043 63291
rect 28534 63288 28540 63300
rect 28031 63260 28540 63288
rect 28031 63257 28043 63260
rect 27985 63251 28043 63257
rect 28534 63248 28540 63260
rect 28592 63288 28598 63300
rect 28644 63288 28672 63319
rect 29086 63316 29092 63328
rect 29144 63316 29150 63368
rect 29822 63356 29828 63368
rect 29783 63328 29828 63356
rect 29822 63316 29828 63328
rect 29880 63316 29886 63368
rect 28592 63260 28672 63288
rect 28592 63248 28598 63260
rect 29270 63248 29276 63300
rect 29328 63288 29334 63300
rect 29730 63288 29736 63300
rect 29328 63260 29736 63288
rect 29328 63248 29334 63260
rect 29730 63248 29736 63260
rect 29788 63248 29794 63300
rect 30374 63248 30380 63300
rect 30432 63288 30438 63300
rect 30558 63288 30564 63300
rect 30432 63260 30564 63288
rect 30432 63248 30438 63260
rect 30558 63248 30564 63260
rect 30616 63248 30622 63300
rect 27019 63192 27844 63220
rect 27019 63189 27031 63192
rect 26973 63183 27031 63189
rect 29546 63180 29552 63232
rect 29604 63220 29610 63232
rect 30009 63223 30067 63229
rect 30009 63220 30021 63223
rect 29604 63192 30021 63220
rect 29604 63180 29610 63192
rect 30009 63189 30021 63192
rect 30055 63189 30067 63223
rect 30009 63183 30067 63189
rect 1104 63130 30820 63152
rect 1104 63078 10880 63130
rect 10932 63078 10944 63130
rect 10996 63078 11008 63130
rect 11060 63078 11072 63130
rect 11124 63078 11136 63130
rect 11188 63078 20811 63130
rect 20863 63078 20875 63130
rect 20927 63078 20939 63130
rect 20991 63078 21003 63130
rect 21055 63078 21067 63130
rect 21119 63078 30820 63130
rect 1104 63056 30820 63078
rect 17862 63016 17868 63028
rect 13004 62988 17868 63016
rect 11330 62908 11336 62960
rect 11388 62948 11394 62960
rect 13004 62957 13032 62988
rect 17862 62976 17868 62988
rect 17920 62976 17926 63028
rect 26970 63016 26976 63028
rect 26436 62988 26976 63016
rect 12805 62951 12863 62957
rect 12805 62948 12817 62951
rect 11388 62920 12817 62948
rect 11388 62908 11394 62920
rect 12805 62917 12817 62920
rect 12851 62917 12863 62951
rect 12805 62911 12863 62917
rect 12989 62951 13047 62957
rect 12989 62917 13001 62951
rect 13035 62917 13047 62951
rect 12989 62911 13047 62917
rect 1578 62880 1584 62892
rect 1539 62852 1584 62880
rect 1578 62840 1584 62852
rect 1636 62840 1642 62892
rect 12621 62883 12679 62889
rect 12621 62849 12633 62883
rect 12667 62880 12679 62883
rect 12710 62880 12716 62892
rect 12667 62852 12716 62880
rect 12667 62849 12679 62852
rect 12621 62843 12679 62849
rect 12710 62840 12716 62852
rect 12768 62840 12774 62892
rect 17402 62840 17408 62892
rect 17460 62889 17466 62892
rect 17460 62883 17509 62889
rect 17460 62849 17463 62883
rect 17497 62849 17509 62883
rect 17460 62843 17509 62849
rect 17570 62886 17628 62892
rect 17570 62852 17582 62886
rect 17616 62852 17628 62886
rect 17570 62846 17628 62852
rect 17702 62886 17760 62892
rect 17702 62852 17714 62886
rect 17748 62852 17760 62886
rect 17702 62846 17760 62852
rect 17460 62840 17466 62843
rect 17218 62772 17224 62824
rect 17276 62812 17282 62824
rect 17584 62812 17612 62846
rect 17276 62784 17612 62812
rect 17717 62812 17745 62846
rect 17862 62840 17868 62892
rect 17920 62880 17926 62892
rect 19337 62883 19395 62889
rect 17920 62852 17965 62880
rect 17920 62840 17926 62852
rect 19337 62849 19349 62883
rect 19383 62880 19395 62883
rect 19426 62880 19432 62892
rect 19383 62852 19432 62880
rect 19383 62849 19395 62852
rect 19337 62843 19395 62849
rect 19426 62840 19432 62852
rect 19484 62840 19490 62892
rect 20346 62880 20352 62892
rect 20307 62852 20352 62880
rect 20346 62840 20352 62852
rect 20404 62840 20410 62892
rect 23569 62883 23627 62889
rect 23569 62849 23581 62883
rect 23615 62880 23627 62883
rect 23842 62880 23848 62892
rect 23615 62852 23848 62880
rect 23615 62849 23627 62852
rect 23569 62843 23627 62849
rect 23842 62840 23848 62852
rect 23900 62840 23906 62892
rect 18414 62812 18420 62824
rect 17717 62784 18420 62812
rect 17276 62772 17282 62784
rect 18414 62772 18420 62784
rect 18472 62772 18478 62824
rect 24578 62772 24584 62824
rect 24636 62812 24642 62824
rect 26436 62812 26464 62988
rect 26970 62976 26976 62988
rect 27028 62976 27034 63028
rect 27709 63019 27767 63025
rect 27709 62985 27721 63019
rect 27755 63016 27767 63019
rect 28626 63016 28632 63028
rect 27755 62988 28632 63016
rect 27755 62985 27767 62988
rect 27709 62979 27767 62985
rect 28626 62976 28632 62988
rect 28684 62976 28690 63028
rect 29178 62976 29184 63028
rect 29236 63016 29242 63028
rect 30101 63019 30159 63025
rect 30101 63016 30113 63019
rect 29236 62988 30113 63016
rect 29236 62976 29242 62988
rect 30101 62985 30113 62988
rect 30147 62985 30159 63019
rect 30101 62979 30159 62985
rect 28902 62948 28908 62960
rect 27920 62920 28908 62948
rect 26973 62883 27031 62889
rect 26973 62849 26985 62883
rect 27019 62880 27031 62883
rect 27614 62880 27620 62892
rect 27019 62852 27620 62880
rect 27019 62849 27031 62852
rect 26973 62843 27031 62849
rect 27614 62840 27620 62852
rect 27672 62840 27678 62892
rect 27920 62889 27948 62920
rect 28902 62908 28908 62920
rect 28960 62908 28966 62960
rect 29012 62920 29776 62948
rect 27920 62883 27997 62889
rect 27920 62852 27951 62883
rect 27939 62849 27951 62852
rect 27985 62849 27997 62883
rect 27939 62843 27997 62849
rect 28058 62883 28116 62889
rect 28058 62849 28070 62883
rect 28104 62880 28116 62883
rect 28190 62883 28248 62889
rect 28104 62849 28120 62880
rect 28058 62843 28120 62849
rect 28190 62849 28202 62883
rect 28236 62849 28248 62883
rect 28190 62843 28248 62849
rect 28353 62883 28411 62889
rect 28353 62849 28365 62883
rect 28399 62880 28411 62883
rect 28534 62880 28540 62892
rect 28399 62852 28540 62880
rect 28399 62849 28411 62852
rect 28353 62843 28411 62849
rect 26510 62812 26516 62824
rect 24636 62784 24992 62812
rect 26436 62784 26516 62812
rect 24636 62772 24642 62784
rect 15194 62704 15200 62756
rect 15252 62744 15258 62756
rect 17310 62744 17316 62756
rect 15252 62716 17316 62744
rect 15252 62704 15258 62716
rect 17310 62704 17316 62716
rect 17368 62704 17374 62756
rect 24964 62744 24992 62784
rect 26510 62772 26516 62784
rect 26568 62772 26574 62824
rect 28092 62812 28120 62843
rect 28205 62812 28233 62843
rect 28534 62840 28540 62852
rect 28592 62840 28598 62892
rect 28626 62812 28632 62824
rect 28092 62784 28133 62812
rect 28205 62784 28632 62812
rect 28105 62756 28133 62784
rect 28626 62772 28632 62784
rect 28684 62772 28690 62824
rect 24964 62716 27844 62744
rect 1397 62679 1455 62685
rect 1397 62645 1409 62679
rect 1443 62676 1455 62679
rect 11330 62676 11336 62688
rect 1443 62648 11336 62676
rect 1443 62645 1455 62648
rect 1397 62639 1455 62645
rect 11330 62636 11336 62648
rect 11388 62636 11394 62688
rect 15102 62636 15108 62688
rect 15160 62676 15166 62688
rect 16482 62676 16488 62688
rect 15160 62648 16488 62676
rect 15160 62636 15166 62648
rect 16482 62636 16488 62648
rect 16540 62636 16546 62688
rect 17221 62679 17279 62685
rect 17221 62645 17233 62679
rect 17267 62676 17279 62679
rect 17402 62676 17408 62688
rect 17267 62648 17408 62676
rect 17267 62645 17279 62648
rect 17221 62639 17279 62645
rect 17402 62636 17408 62648
rect 17460 62636 17466 62688
rect 19521 62679 19579 62685
rect 19521 62645 19533 62679
rect 19567 62676 19579 62679
rect 19978 62676 19984 62688
rect 19567 62648 19984 62676
rect 19567 62645 19579 62648
rect 19521 62639 19579 62645
rect 19978 62636 19984 62648
rect 20036 62636 20042 62688
rect 20533 62679 20591 62685
rect 20533 62645 20545 62679
rect 20579 62676 20591 62679
rect 21082 62676 21088 62688
rect 20579 62648 21088 62676
rect 20579 62645 20591 62648
rect 20533 62639 20591 62645
rect 21082 62636 21088 62648
rect 21140 62636 21146 62688
rect 23753 62679 23811 62685
rect 23753 62645 23765 62679
rect 23799 62676 23811 62679
rect 24026 62676 24032 62688
rect 23799 62648 24032 62676
rect 23799 62645 23811 62648
rect 23753 62639 23811 62645
rect 24026 62636 24032 62648
rect 24084 62636 24090 62688
rect 27154 62676 27160 62688
rect 27067 62648 27160 62676
rect 27154 62636 27160 62648
rect 27212 62676 27218 62688
rect 27338 62676 27344 62688
rect 27212 62648 27344 62676
rect 27212 62636 27218 62648
rect 27338 62636 27344 62648
rect 27396 62636 27402 62688
rect 27816 62676 27844 62716
rect 28074 62704 28080 62756
rect 28132 62704 28138 62756
rect 28534 62704 28540 62756
rect 28592 62744 28598 62756
rect 29012 62744 29040 62920
rect 29362 62880 29368 62892
rect 29323 62852 29368 62880
rect 29362 62840 29368 62852
rect 29420 62840 29426 62892
rect 29549 62883 29607 62889
rect 29549 62849 29561 62883
rect 29595 62849 29607 62883
rect 29549 62843 29607 62849
rect 29178 62772 29184 62824
rect 29236 62812 29242 62824
rect 29564 62812 29592 62843
rect 29748 62821 29776 62920
rect 29917 62883 29975 62889
rect 29917 62849 29929 62883
rect 29963 62880 29975 62883
rect 30006 62880 30012 62892
rect 29963 62852 30012 62880
rect 29963 62849 29975 62852
rect 29917 62843 29975 62849
rect 30006 62840 30012 62852
rect 30064 62840 30070 62892
rect 29236 62784 29592 62812
rect 29641 62815 29699 62821
rect 29236 62772 29242 62784
rect 29641 62781 29653 62815
rect 29687 62781 29699 62815
rect 29641 62775 29699 62781
rect 29733 62815 29791 62821
rect 29733 62781 29745 62815
rect 29779 62781 29791 62815
rect 29733 62775 29791 62781
rect 28592 62716 29040 62744
rect 28592 62704 28598 62716
rect 29656 62676 29684 62775
rect 27816 62648 29684 62676
rect 1104 62586 30820 62608
rect 1104 62534 5915 62586
rect 5967 62534 5979 62586
rect 6031 62534 6043 62586
rect 6095 62534 6107 62586
rect 6159 62534 6171 62586
rect 6223 62534 15846 62586
rect 15898 62534 15910 62586
rect 15962 62534 15974 62586
rect 16026 62534 16038 62586
rect 16090 62534 16102 62586
rect 16154 62534 25776 62586
rect 25828 62534 25840 62586
rect 25892 62534 25904 62586
rect 25956 62534 25968 62586
rect 26020 62534 26032 62586
rect 26084 62534 30820 62586
rect 1104 62512 30820 62534
rect 18322 62472 18328 62484
rect 16040 62444 18328 62472
rect 16040 62416 16068 62444
rect 18322 62432 18328 62444
rect 18380 62432 18386 62484
rect 23661 62475 23719 62481
rect 23661 62441 23673 62475
rect 23707 62472 23719 62475
rect 24394 62472 24400 62484
rect 23707 62444 24400 62472
rect 23707 62441 23719 62444
rect 23661 62435 23719 62441
rect 24394 62432 24400 62444
rect 24452 62432 24458 62484
rect 26881 62475 26939 62481
rect 26881 62441 26893 62475
rect 26927 62472 26939 62475
rect 28350 62472 28356 62484
rect 26927 62444 28356 62472
rect 26927 62441 26939 62444
rect 26881 62435 26939 62441
rect 28350 62432 28356 62444
rect 28408 62432 28414 62484
rect 29454 62432 29460 62484
rect 29512 62472 29518 62484
rect 29549 62475 29607 62481
rect 29549 62472 29561 62475
rect 29512 62444 29561 62472
rect 29512 62432 29518 62444
rect 29549 62441 29561 62444
rect 29595 62441 29607 62475
rect 29549 62435 29607 62441
rect 16022 62364 16028 62416
rect 16080 62364 16086 62416
rect 22465 62407 22523 62413
rect 22465 62373 22477 62407
rect 22511 62373 22523 62407
rect 22465 62367 22523 62373
rect 16850 62336 16856 62348
rect 16316 62308 16856 62336
rect 16022 62228 16028 62280
rect 16080 62277 16086 62280
rect 16080 62271 16129 62277
rect 16080 62237 16083 62271
rect 16117 62237 16129 62271
rect 16206 62268 16212 62280
rect 16167 62240 16212 62268
rect 16080 62231 16129 62237
rect 16080 62228 16086 62231
rect 16206 62228 16212 62240
rect 16264 62228 16270 62280
rect 16316 62277 16344 62308
rect 16850 62296 16856 62308
rect 16908 62296 16914 62348
rect 21082 62336 21088 62348
rect 21043 62308 21088 62336
rect 21082 62296 21088 62308
rect 21140 62296 21146 62348
rect 22094 62296 22100 62348
rect 22152 62336 22158 62348
rect 22480 62336 22508 62367
rect 24946 62364 24952 62416
rect 25004 62364 25010 62416
rect 23293 62339 23351 62345
rect 23293 62336 23305 62339
rect 22152 62308 23305 62336
rect 22152 62296 22158 62308
rect 23293 62305 23305 62308
rect 23339 62305 23351 62339
rect 24964 62336 24992 62364
rect 23293 62299 23351 62305
rect 24688 62308 24992 62336
rect 16301 62271 16359 62277
rect 16301 62237 16313 62271
rect 16347 62237 16359 62271
rect 16301 62231 16359 62237
rect 16482 62228 16488 62280
rect 16540 62268 16546 62280
rect 17310 62268 17316 62280
rect 16540 62240 16585 62268
rect 17271 62240 17316 62268
rect 16540 62228 16546 62240
rect 17310 62228 17316 62240
rect 17368 62228 17374 62280
rect 17402 62228 17408 62280
rect 17460 62268 17466 62280
rect 17569 62271 17627 62277
rect 17569 62268 17581 62271
rect 17460 62240 17581 62268
rect 17460 62228 17466 62240
rect 17569 62237 17581 62240
rect 17615 62237 17627 62271
rect 23474 62268 23480 62280
rect 23435 62240 23480 62268
rect 17569 62231 17627 62237
rect 23474 62228 23480 62240
rect 23532 62228 23538 62280
rect 24688 62277 24716 62308
rect 26142 62296 26148 62348
rect 26200 62336 26206 62348
rect 26200 62308 27384 62336
rect 26200 62296 26206 62308
rect 24673 62271 24731 62277
rect 24673 62237 24685 62271
rect 24719 62237 24731 62271
rect 24854 62268 24860 62280
rect 24815 62240 24860 62268
rect 24673 62231 24731 62237
rect 24854 62228 24860 62240
rect 24912 62228 24918 62280
rect 24949 62271 25007 62277
rect 24949 62237 24961 62271
rect 24995 62268 25007 62271
rect 25222 62268 25228 62280
rect 24995 62240 25228 62268
rect 24995 62237 25007 62240
rect 24949 62231 25007 62237
rect 25222 62228 25228 62240
rect 25280 62228 25286 62280
rect 26970 62228 26976 62280
rect 27028 62268 27034 62280
rect 27111 62271 27169 62277
rect 27111 62268 27123 62271
rect 27028 62240 27123 62268
rect 27028 62228 27034 62240
rect 27111 62237 27123 62240
rect 27157 62237 27169 62271
rect 27246 62268 27252 62280
rect 27207 62240 27252 62268
rect 27111 62231 27169 62237
rect 27246 62228 27252 62240
rect 27304 62228 27310 62280
rect 27356 62277 27384 62308
rect 27706 62296 27712 62348
rect 27764 62336 27770 62348
rect 28626 62336 28632 62348
rect 27764 62308 28632 62336
rect 27764 62296 27770 62308
rect 28626 62296 28632 62308
rect 28684 62296 28690 62348
rect 29270 62296 29276 62348
rect 29328 62336 29334 62348
rect 29454 62336 29460 62348
rect 29328 62308 29460 62336
rect 29328 62296 29334 62308
rect 29454 62296 29460 62308
rect 29512 62296 29518 62348
rect 27341 62271 27399 62277
rect 27341 62237 27353 62271
rect 27387 62237 27399 62271
rect 27341 62231 27399 62237
rect 27430 62228 27436 62280
rect 27488 62268 27494 62280
rect 27525 62271 27583 62277
rect 27525 62268 27537 62271
rect 27488 62240 27537 62268
rect 27488 62228 27494 62240
rect 27525 62237 27537 62240
rect 27571 62237 27583 62271
rect 27525 62231 27583 62237
rect 27632 62240 28764 62268
rect 14829 62203 14887 62209
rect 14829 62169 14841 62203
rect 14875 62200 14887 62203
rect 16758 62200 16764 62212
rect 14875 62172 16764 62200
rect 14875 62169 14887 62172
rect 14829 62163 14887 62169
rect 16758 62160 16764 62172
rect 16816 62160 16822 62212
rect 21352 62203 21410 62209
rect 21352 62169 21364 62203
rect 21398 62200 21410 62203
rect 21818 62200 21824 62212
rect 21398 62172 21824 62200
rect 21398 62169 21410 62172
rect 21352 62163 21410 62169
rect 21818 62160 21824 62172
rect 21876 62160 21882 62212
rect 27632 62200 27660 62240
rect 28626 62200 28632 62212
rect 22066 62172 27660 62200
rect 28587 62172 28632 62200
rect 14642 62092 14648 62144
rect 14700 62132 14706 62144
rect 14921 62135 14979 62141
rect 14921 62132 14933 62135
rect 14700 62104 14933 62132
rect 14700 62092 14706 62104
rect 14921 62101 14933 62104
rect 14967 62101 14979 62135
rect 14921 62095 14979 62101
rect 15841 62135 15899 62141
rect 15841 62101 15853 62135
rect 15887 62132 15899 62135
rect 16666 62132 16672 62144
rect 15887 62104 16672 62132
rect 15887 62101 15899 62104
rect 15841 62095 15899 62101
rect 16666 62092 16672 62104
rect 16724 62092 16730 62144
rect 17494 62092 17500 62144
rect 17552 62132 17558 62144
rect 18690 62132 18696 62144
rect 17552 62104 18696 62132
rect 17552 62092 17558 62104
rect 18690 62092 18696 62104
rect 18748 62092 18754 62144
rect 18874 62092 18880 62144
rect 18932 62132 18938 62144
rect 22066 62132 22094 62172
rect 28626 62160 28632 62172
rect 28684 62160 28690 62212
rect 28736 62200 28764 62240
rect 29086 62228 29092 62280
rect 29144 62268 29150 62280
rect 29733 62271 29791 62277
rect 29733 62268 29745 62271
rect 29144 62240 29745 62268
rect 29144 62228 29150 62240
rect 29733 62237 29745 62240
rect 29779 62237 29791 62271
rect 30006 62268 30012 62280
rect 29967 62240 30012 62268
rect 29733 62231 29791 62237
rect 30006 62228 30012 62240
rect 30064 62228 30070 62280
rect 29917 62203 29975 62209
rect 29917 62200 29929 62203
rect 28736 62172 29929 62200
rect 29917 62169 29929 62172
rect 29963 62169 29975 62203
rect 29917 62163 29975 62169
rect 18932 62104 22094 62132
rect 24489 62135 24547 62141
rect 18932 62092 18938 62104
rect 24489 62101 24501 62135
rect 24535 62132 24547 62135
rect 25958 62132 25964 62144
rect 24535 62104 25964 62132
rect 24535 62101 24547 62104
rect 24489 62095 24547 62101
rect 25958 62092 25964 62104
rect 26016 62092 26022 62144
rect 26418 62092 26424 62144
rect 26476 62132 26482 62144
rect 27890 62132 27896 62144
rect 26476 62104 27896 62132
rect 26476 62092 26482 62104
rect 27890 62092 27896 62104
rect 27948 62132 27954 62144
rect 28721 62135 28779 62141
rect 28721 62132 28733 62135
rect 27948 62104 28733 62132
rect 27948 62092 27954 62104
rect 28721 62101 28733 62104
rect 28767 62101 28779 62135
rect 28721 62095 28779 62101
rect 1104 62042 30820 62064
rect 1104 61990 10880 62042
rect 10932 61990 10944 62042
rect 10996 61990 11008 62042
rect 11060 61990 11072 62042
rect 11124 61990 11136 62042
rect 11188 61990 20811 62042
rect 20863 61990 20875 62042
rect 20927 61990 20939 62042
rect 20991 61990 21003 62042
rect 21055 61990 21067 62042
rect 21119 61990 30820 62042
rect 1104 61968 30820 61990
rect 14090 61888 14096 61940
rect 14148 61928 14154 61940
rect 16850 61928 16856 61940
rect 14148 61900 16856 61928
rect 14148 61888 14154 61900
rect 11238 61820 11244 61872
rect 11296 61860 11302 61872
rect 12713 61863 12771 61869
rect 12713 61860 12725 61863
rect 11296 61832 12725 61860
rect 11296 61820 11302 61832
rect 12713 61829 12725 61832
rect 12759 61829 12771 61863
rect 12713 61823 12771 61829
rect 1578 61792 1584 61804
rect 1539 61764 1584 61792
rect 1578 61752 1584 61764
rect 1636 61752 1642 61804
rect 12526 61792 12532 61804
rect 12487 61764 12532 61792
rect 12526 61752 12532 61764
rect 12584 61752 12590 61804
rect 15194 61792 15200 61804
rect 15155 61764 15200 61792
rect 15194 61752 15200 61764
rect 15252 61752 15258 61804
rect 15396 61801 15424 61900
rect 16850 61888 16856 61900
rect 16908 61888 16914 61940
rect 21818 61928 21824 61940
rect 21779 61900 21824 61928
rect 21818 61888 21824 61900
rect 21876 61888 21882 61940
rect 24673 61931 24731 61937
rect 24673 61897 24685 61931
rect 24719 61928 24731 61931
rect 24762 61928 24768 61940
rect 24719 61900 24768 61928
rect 24719 61897 24731 61900
rect 24673 61891 24731 61897
rect 24762 61888 24768 61900
rect 24820 61888 24826 61940
rect 25038 61928 25044 61940
rect 24999 61900 25044 61928
rect 25038 61888 25044 61900
rect 25096 61888 25102 61940
rect 25682 61928 25688 61940
rect 25643 61900 25688 61928
rect 25682 61888 25688 61900
rect 25740 61888 25746 61940
rect 26973 61931 27031 61937
rect 26973 61897 26985 61931
rect 27019 61928 27031 61931
rect 27019 61900 28304 61928
rect 27019 61897 27031 61900
rect 26973 61891 27031 61897
rect 19702 61860 19708 61872
rect 16684 61832 19708 61860
rect 15286 61795 15344 61801
rect 15286 61761 15298 61795
rect 15332 61761 15344 61795
rect 15286 61755 15344 61761
rect 15381 61795 15439 61801
rect 15381 61761 15393 61795
rect 15427 61761 15439 61795
rect 15381 61755 15439 61761
rect 15304 61724 15332 61755
rect 15562 61752 15568 61804
rect 15620 61792 15626 61804
rect 15620 61764 15665 61792
rect 15620 61752 15626 61764
rect 16574 61752 16580 61804
rect 16632 61792 16638 61804
rect 16684 61801 16712 61832
rect 19702 61820 19708 61832
rect 19760 61820 19766 61872
rect 21174 61820 21180 61872
rect 21232 61860 21238 61872
rect 22370 61860 22376 61872
rect 21232 61832 22376 61860
rect 21232 61820 21238 61832
rect 18782 61801 18788 61804
rect 16669 61795 16727 61801
rect 16669 61792 16681 61795
rect 16632 61764 16681 61792
rect 16632 61752 16638 61764
rect 16669 61761 16681 61764
rect 16715 61761 16727 61795
rect 16669 61755 16727 61761
rect 18776 61755 18788 61801
rect 18840 61792 18846 61804
rect 22094 61792 22100 61804
rect 18840 61764 18876 61792
rect 22055 61764 22100 61792
rect 18782 61752 18788 61755
rect 18840 61752 18846 61764
rect 22094 61752 22100 61764
rect 22152 61752 22158 61804
rect 22296 61801 22324 61832
rect 22370 61820 22376 61832
rect 22428 61820 22434 61872
rect 24228 61832 25084 61860
rect 22186 61795 22244 61801
rect 22186 61761 22198 61795
rect 22232 61761 22244 61795
rect 22186 61755 22244 61761
rect 22286 61795 22344 61801
rect 22286 61761 22298 61795
rect 22332 61761 22344 61795
rect 22462 61792 22468 61804
rect 22423 61764 22468 61792
rect 22286 61755 22344 61761
rect 16206 61724 16212 61736
rect 15304 61696 16212 61724
rect 16206 61684 16212 61696
rect 16264 61724 16270 61736
rect 16945 61727 17003 61733
rect 16945 61724 16957 61727
rect 16264 61696 16957 61724
rect 16264 61684 16270 61696
rect 16945 61693 16957 61696
rect 16991 61724 17003 61727
rect 17218 61724 17224 61736
rect 16991 61696 17224 61724
rect 16991 61693 17003 61696
rect 16945 61687 17003 61693
rect 17218 61684 17224 61696
rect 17276 61724 17282 61736
rect 17494 61724 17500 61736
rect 17276 61696 17500 61724
rect 17276 61684 17282 61696
rect 17494 61684 17500 61696
rect 17552 61684 17558 61736
rect 18506 61724 18512 61736
rect 18467 61696 18512 61724
rect 18506 61684 18512 61696
rect 18564 61684 18570 61736
rect 22002 61684 22008 61736
rect 22060 61724 22066 61736
rect 22201 61724 22229 61755
rect 22462 61752 22468 61764
rect 22520 61752 22526 61804
rect 23293 61795 23351 61801
rect 23293 61761 23305 61795
rect 23339 61792 23351 61795
rect 23842 61792 23848 61804
rect 23339 61764 23848 61792
rect 23339 61761 23351 61764
rect 23293 61755 23351 61761
rect 23842 61752 23848 61764
rect 23900 61752 23906 61804
rect 23937 61795 23995 61801
rect 23937 61761 23949 61795
rect 23983 61761 23995 61795
rect 24118 61792 24124 61804
rect 24079 61764 24124 61792
rect 23937 61755 23995 61761
rect 23952 61724 23980 61755
rect 24118 61752 24124 61764
rect 24176 61752 24182 61804
rect 24228 61801 24256 61832
rect 24213 61795 24271 61801
rect 24213 61761 24225 61795
rect 24259 61761 24271 61795
rect 24213 61755 24271 61761
rect 24486 61752 24492 61804
rect 24544 61792 24550 61804
rect 24544 61764 24808 61792
rect 24544 61752 24550 61764
rect 22060 61696 22229 61724
rect 23676 61696 23980 61724
rect 24780 61724 24808 61764
rect 24854 61752 24860 61804
rect 24912 61792 24918 61804
rect 25056 61792 25084 61832
rect 25958 61820 25964 61872
rect 26016 61860 26022 61872
rect 28276 61860 28304 61900
rect 30650 61860 30656 61872
rect 26016 61832 27660 61860
rect 28276 61832 30656 61860
rect 26016 61820 26022 61832
rect 25133 61795 25191 61801
rect 25133 61792 25145 61795
rect 24912 61764 24957 61792
rect 25056 61764 25145 61792
rect 24912 61752 24918 61764
rect 25133 61761 25145 61764
rect 25179 61792 25191 61795
rect 25222 61792 25228 61804
rect 25179 61764 25228 61792
rect 25179 61761 25191 61764
rect 25133 61755 25191 61761
rect 25222 61752 25228 61764
rect 25280 61752 25286 61804
rect 25682 61752 25688 61804
rect 25740 61792 25746 61804
rect 25869 61795 25927 61801
rect 25869 61792 25881 61795
rect 25740 61764 25881 61792
rect 25740 61752 25746 61764
rect 25869 61761 25881 61764
rect 25915 61761 25927 61795
rect 25869 61755 25927 61761
rect 26053 61795 26111 61801
rect 26053 61761 26065 61795
rect 26099 61761 26111 61795
rect 26053 61755 26111 61761
rect 26145 61795 26203 61801
rect 26145 61761 26157 61795
rect 26191 61792 26203 61795
rect 26326 61792 26332 61804
rect 26191 61764 26332 61792
rect 26191 61761 26203 61764
rect 26145 61755 26203 61761
rect 26068 61724 26096 61755
rect 26326 61752 26332 61764
rect 26384 61752 26390 61804
rect 26970 61752 26976 61804
rect 27028 61792 27034 61804
rect 27249 61795 27307 61801
rect 27249 61792 27261 61795
rect 27028 61764 27261 61792
rect 27028 61752 27034 61764
rect 27249 61761 27261 61764
rect 27295 61761 27307 61795
rect 27341 61795 27399 61801
rect 27341 61788 27353 61795
rect 27387 61788 27399 61795
rect 27433 61795 27491 61801
rect 27249 61755 27307 61761
rect 27338 61736 27344 61788
rect 27396 61736 27402 61788
rect 27433 61761 27445 61795
rect 27479 61792 27491 61795
rect 27522 61792 27528 61804
rect 27479 61764 27528 61792
rect 27479 61761 27491 61764
rect 27433 61755 27491 61761
rect 27522 61752 27528 61764
rect 27580 61752 27586 61804
rect 27632 61801 27660 61832
rect 30650 61820 30656 61832
rect 30708 61820 30714 61872
rect 27617 61795 27675 61801
rect 27617 61761 27629 61795
rect 27663 61761 27675 61795
rect 27617 61755 27675 61761
rect 28169 61795 28227 61801
rect 28169 61761 28181 61795
rect 28215 61792 28227 61795
rect 28350 61792 28356 61804
rect 28215 61764 28356 61792
rect 28215 61761 28227 61764
rect 28169 61755 28227 61761
rect 28350 61752 28356 61764
rect 28408 61752 28414 61804
rect 28718 61752 28724 61804
rect 28776 61752 28782 61804
rect 29178 61792 29184 61804
rect 29139 61764 29184 61792
rect 29178 61752 29184 61764
rect 29236 61752 29242 61804
rect 28736 61724 28764 61752
rect 24780 61696 26096 61724
rect 28000 61696 28764 61724
rect 28905 61727 28963 61733
rect 22060 61684 22066 61696
rect 1397 61591 1455 61597
rect 1397 61557 1409 61591
rect 1443 61588 1455 61591
rect 7558 61588 7564 61600
rect 1443 61560 7564 61588
rect 1443 61557 1455 61560
rect 1397 61551 1455 61557
rect 7558 61548 7564 61560
rect 7616 61548 7622 61600
rect 12897 61591 12955 61597
rect 12897 61557 12909 61591
rect 12943 61588 12955 61591
rect 14734 61588 14740 61600
rect 12943 61560 14740 61588
rect 12943 61557 12955 61560
rect 12897 61551 12955 61557
rect 14734 61548 14740 61560
rect 14792 61548 14798 61600
rect 14918 61588 14924 61600
rect 14879 61560 14924 61588
rect 14918 61548 14924 61560
rect 14976 61548 14982 61600
rect 19150 61548 19156 61600
rect 19208 61588 19214 61600
rect 19889 61591 19947 61597
rect 19889 61588 19901 61591
rect 19208 61560 19901 61588
rect 19208 61548 19214 61560
rect 19889 61557 19901 61560
rect 19935 61588 19947 61591
rect 22830 61588 22836 61600
rect 19935 61560 22836 61588
rect 19935 61557 19947 61560
rect 19889 61551 19947 61557
rect 22830 61548 22836 61560
rect 22888 61548 22894 61600
rect 23109 61591 23167 61597
rect 23109 61557 23121 61591
rect 23155 61588 23167 61591
rect 23474 61588 23480 61600
rect 23155 61560 23480 61588
rect 23155 61557 23167 61560
rect 23109 61551 23167 61557
rect 23474 61548 23480 61560
rect 23532 61548 23538 61600
rect 23676 61588 23704 61696
rect 23753 61659 23811 61665
rect 23753 61625 23765 61659
rect 23799 61656 23811 61659
rect 27890 61656 27896 61668
rect 23799 61628 27896 61656
rect 23799 61625 23811 61628
rect 23753 61619 23811 61625
rect 27890 61616 27896 61628
rect 27948 61616 27954 61668
rect 24946 61588 24952 61600
rect 23676 61560 24952 61588
rect 24946 61548 24952 61560
rect 25004 61548 25010 61600
rect 25038 61548 25044 61600
rect 25096 61588 25102 61600
rect 25406 61588 25412 61600
rect 25096 61560 25412 61588
rect 25096 61548 25102 61560
rect 25406 61548 25412 61560
rect 25464 61548 25470 61600
rect 27430 61548 27436 61600
rect 27488 61588 27494 61600
rect 28000 61588 28028 61696
rect 28905 61693 28917 61727
rect 28951 61693 28963 61727
rect 28905 61687 28963 61693
rect 28718 61616 28724 61668
rect 28776 61656 28782 61668
rect 28920 61656 28948 61687
rect 28776 61628 28948 61656
rect 28776 61616 28782 61628
rect 27488 61560 28028 61588
rect 28353 61591 28411 61597
rect 27488 61548 27494 61560
rect 28353 61557 28365 61591
rect 28399 61588 28411 61591
rect 28810 61588 28816 61600
rect 28399 61560 28816 61588
rect 28399 61557 28411 61560
rect 28353 61551 28411 61557
rect 28810 61548 28816 61560
rect 28868 61548 28874 61600
rect 1104 61498 30820 61520
rect 1104 61446 5915 61498
rect 5967 61446 5979 61498
rect 6031 61446 6043 61498
rect 6095 61446 6107 61498
rect 6159 61446 6171 61498
rect 6223 61446 15846 61498
rect 15898 61446 15910 61498
rect 15962 61446 15974 61498
rect 16026 61446 16038 61498
rect 16090 61446 16102 61498
rect 16154 61446 25776 61498
rect 25828 61446 25840 61498
rect 25892 61446 25904 61498
rect 25956 61446 25968 61498
rect 26020 61446 26032 61498
rect 26084 61446 30820 61498
rect 1104 61424 30820 61446
rect 15378 61344 15384 61396
rect 15436 61384 15442 61396
rect 16390 61384 16396 61396
rect 15436 61356 16396 61384
rect 15436 61344 15442 61356
rect 16390 61344 16396 61356
rect 16448 61344 16454 61396
rect 18506 61344 18512 61396
rect 18564 61384 18570 61396
rect 18693 61387 18751 61393
rect 18693 61384 18705 61387
rect 18564 61356 18705 61384
rect 18564 61344 18570 61356
rect 18693 61353 18705 61356
rect 18739 61353 18751 61387
rect 18693 61347 18751 61353
rect 24670 61344 24676 61396
rect 24728 61384 24734 61396
rect 25406 61384 25412 61396
rect 24728 61356 25412 61384
rect 24728 61344 24734 61356
rect 25406 61344 25412 61356
rect 25464 61344 25470 61396
rect 27249 61387 27307 61393
rect 27249 61353 27261 61387
rect 27295 61353 27307 61387
rect 27249 61347 27307 61353
rect 14461 61319 14519 61325
rect 14461 61285 14473 61319
rect 14507 61316 14519 61319
rect 20162 61316 20168 61328
rect 14507 61288 20168 61316
rect 14507 61285 14519 61288
rect 14461 61279 14519 61285
rect 20162 61276 20168 61288
rect 20220 61276 20226 61328
rect 27264 61316 27292 61347
rect 27430 61344 27436 61396
rect 27488 61384 27494 61396
rect 28537 61387 28595 61393
rect 28537 61384 28549 61387
rect 27488 61356 28549 61384
rect 27488 61344 27494 61356
rect 28537 61353 28549 61356
rect 28583 61353 28595 61387
rect 29549 61387 29607 61393
rect 29549 61384 29561 61387
rect 28537 61347 28595 61353
rect 29288 61356 29561 61384
rect 29288 61328 29316 61356
rect 29549 61353 29561 61356
rect 29595 61353 29607 61387
rect 29549 61347 29607 61353
rect 29730 61344 29736 61396
rect 29788 61344 29794 61396
rect 28810 61316 28816 61328
rect 27264 61288 28816 61316
rect 28810 61276 28816 61288
rect 28868 61276 28874 61328
rect 29086 61276 29092 61328
rect 29144 61276 29150 61328
rect 29270 61276 29276 61328
rect 29328 61276 29334 61328
rect 29362 61276 29368 61328
rect 29420 61316 29426 61328
rect 29748 61316 29776 61344
rect 29420 61288 29776 61316
rect 29420 61276 29426 61288
rect 7558 61208 7564 61260
rect 7616 61248 7622 61260
rect 7616 61220 14320 61248
rect 7616 61208 7622 61220
rect 1578 61180 1584 61192
rect 1539 61152 1584 61180
rect 1578 61140 1584 61152
rect 1636 61140 1642 61192
rect 12894 61180 12900 61192
rect 12807 61152 12900 61180
rect 12894 61140 12900 61152
rect 12952 61180 12958 61192
rect 13446 61180 13452 61192
rect 12952 61152 13452 61180
rect 12952 61140 12958 61152
rect 13446 61140 13452 61152
rect 13504 61140 13510 61192
rect 14292 61189 14320 61220
rect 15194 61208 15200 61260
rect 15252 61248 15258 61260
rect 15654 61248 15660 61260
rect 15252 61220 15660 61248
rect 15252 61208 15258 61220
rect 15654 61208 15660 61220
rect 15712 61208 15718 61260
rect 16850 61208 16856 61260
rect 16908 61248 16914 61260
rect 16908 61220 17908 61248
rect 16908 61208 16914 61220
rect 14277 61183 14335 61189
rect 14277 61149 14289 61183
rect 14323 61149 14335 61183
rect 14277 61143 14335 61149
rect 17402 61140 17408 61192
rect 17460 61180 17466 61192
rect 17589 61183 17647 61189
rect 17589 61180 17601 61183
rect 17460 61152 17601 61180
rect 17460 61140 17466 61152
rect 17589 61149 17601 61152
rect 17635 61149 17647 61183
rect 17694 61183 17752 61189
rect 17694 61156 17706 61183
rect 17589 61143 17647 61149
rect 17677 61149 17706 61156
rect 17740 61149 17752 61183
rect 17677 61143 17752 61149
rect 17794 61180 17852 61186
rect 17794 61146 17806 61180
rect 17840 61177 17852 61180
rect 17880 61177 17908 61220
rect 18322 61208 18328 61260
rect 18380 61248 18386 61260
rect 23934 61248 23940 61260
rect 18380 61220 23940 61248
rect 18380 61208 18386 61220
rect 23934 61208 23940 61220
rect 23992 61248 23998 61260
rect 24854 61248 24860 61260
rect 23992 61220 24860 61248
rect 23992 61208 23998 61220
rect 24854 61208 24860 61220
rect 24912 61208 24918 61260
rect 25869 61251 25927 61257
rect 25869 61217 25881 61251
rect 25915 61248 25927 61251
rect 28626 61248 28632 61260
rect 25915 61220 27752 61248
rect 25915 61217 25927 61220
rect 25869 61211 25927 61217
rect 17840 61149 17908 61177
rect 17840 61146 17852 61149
rect 17677 61128 17724 61143
rect 17794 61140 17852 61146
rect 17954 61140 17960 61192
rect 18012 61180 18018 61192
rect 18506 61180 18512 61192
rect 18012 61152 18057 61180
rect 18467 61152 18512 61180
rect 18012 61140 18018 61152
rect 18506 61140 18512 61152
rect 18564 61140 18570 61192
rect 19702 61180 19708 61192
rect 19663 61152 19708 61180
rect 19702 61140 19708 61152
rect 19760 61180 19766 61192
rect 20254 61180 20260 61192
rect 19760 61152 20260 61180
rect 19760 61140 19766 61152
rect 20254 61140 20260 61152
rect 20312 61140 20318 61192
rect 22370 61140 22376 61192
rect 22428 61180 22434 61192
rect 23293 61183 23351 61189
rect 23293 61180 23305 61183
rect 22428 61152 23305 61180
rect 22428 61140 22434 61152
rect 23293 61149 23305 61152
rect 23339 61149 23351 61183
rect 23293 61143 23351 61149
rect 23474 61140 23480 61192
rect 23532 61180 23538 61192
rect 24397 61183 24455 61189
rect 24397 61180 24409 61183
rect 23532 61152 24409 61180
rect 23532 61140 23538 61152
rect 24397 61149 24409 61152
rect 24443 61149 24455 61183
rect 24397 61143 24455 61149
rect 24673 61183 24731 61189
rect 24673 61149 24685 61183
rect 24719 61180 24731 61183
rect 25222 61180 25228 61192
rect 24719 61152 25228 61180
rect 24719 61149 24731 61152
rect 24673 61143 24731 61149
rect 25222 61140 25228 61152
rect 25280 61140 25286 61192
rect 25682 61140 25688 61192
rect 25740 61180 25746 61192
rect 25958 61180 25964 61192
rect 25740 61152 25964 61180
rect 25740 61140 25746 61152
rect 25958 61140 25964 61152
rect 26016 61180 26022 61192
rect 26053 61183 26111 61189
rect 26053 61180 26065 61183
rect 26016 61152 26065 61180
rect 26016 61140 26022 61152
rect 26053 61149 26065 61152
rect 26099 61149 26111 61183
rect 26326 61180 26332 61192
rect 26287 61152 26332 61180
rect 26053 61143 26111 61149
rect 26326 61140 26332 61152
rect 26384 61140 26390 61192
rect 26970 61140 26976 61192
rect 27028 61180 27034 61192
rect 27724 61189 27752 61220
rect 27816 61220 28632 61248
rect 27525 61183 27583 61189
rect 27525 61180 27537 61183
rect 27028 61152 27537 61180
rect 27028 61140 27034 61152
rect 27525 61149 27537 61152
rect 27571 61149 27583 61183
rect 27525 61143 27583 61149
rect 27617 61183 27675 61189
rect 27617 61149 27629 61183
rect 27663 61149 27675 61183
rect 27617 61143 27675 61149
rect 27709 61183 27767 61189
rect 27709 61149 27721 61183
rect 27755 61149 27767 61183
rect 27709 61143 27767 61149
rect 14093 61115 14151 61121
rect 14093 61112 14105 61115
rect 12728 61084 14105 61112
rect 1397 61047 1455 61053
rect 1397 61013 1409 61047
rect 1443 61044 1455 61047
rect 11238 61044 11244 61056
rect 1443 61016 11244 61044
rect 1443 61013 1455 61016
rect 1397 61007 1455 61013
rect 11238 61004 11244 61016
rect 11296 61004 11302 61056
rect 12526 61004 12532 61056
rect 12584 61044 12590 61056
rect 12728 61053 12756 61084
rect 14093 61081 14105 61084
rect 14139 61081 14151 61115
rect 14093 61075 14151 61081
rect 15105 61115 15163 61121
rect 15105 61081 15117 61115
rect 15151 61112 15163 61115
rect 16206 61112 16212 61124
rect 15151 61084 16212 61112
rect 15151 61081 15163 61084
rect 15105 61075 15163 61081
rect 16206 61072 16212 61084
rect 16264 61072 16270 61124
rect 17494 61072 17500 61124
rect 17552 61112 17558 61124
rect 17677 61112 17705 61128
rect 17552 61084 17705 61112
rect 17552 61072 17558 61084
rect 24854 61072 24860 61124
rect 24912 61112 24918 61124
rect 25590 61112 25596 61124
rect 24912 61084 25596 61112
rect 24912 61072 24918 61084
rect 25590 61072 25596 61084
rect 25648 61072 25654 61124
rect 25774 61072 25780 61124
rect 25832 61112 25838 61124
rect 27632 61112 27660 61143
rect 27816 61112 27844 61220
rect 28626 61208 28632 61220
rect 28684 61208 28690 61260
rect 29104 61248 29132 61276
rect 28736 61220 29776 61248
rect 27890 61140 27896 61192
rect 27948 61180 27954 61192
rect 27948 61152 27993 61180
rect 27948 61140 27954 61152
rect 28442 61140 28448 61192
rect 28500 61180 28506 61192
rect 28736 61189 28764 61220
rect 28721 61183 28779 61189
rect 28721 61180 28733 61183
rect 28500 61152 28733 61180
rect 28500 61140 28506 61152
rect 28721 61149 28733 61152
rect 28767 61149 28779 61183
rect 28721 61143 28779 61149
rect 28810 61140 28816 61192
rect 28868 61180 28874 61192
rect 28905 61183 28963 61189
rect 28905 61180 28917 61183
rect 28868 61152 28917 61180
rect 28868 61140 28874 61152
rect 28905 61149 28917 61152
rect 28951 61149 28963 61183
rect 28905 61143 28963 61149
rect 28997 61183 29055 61189
rect 28997 61149 29009 61183
rect 29043 61180 29055 61183
rect 29086 61180 29092 61192
rect 29043 61152 29092 61180
rect 29043 61149 29055 61152
rect 28997 61143 29055 61149
rect 29086 61140 29092 61152
rect 29144 61140 29150 61192
rect 29748 61189 29776 61220
rect 29733 61183 29791 61189
rect 29733 61149 29745 61183
rect 29779 61149 29791 61183
rect 30006 61180 30012 61192
rect 29967 61152 30012 61180
rect 29733 61143 29791 61149
rect 30006 61140 30012 61152
rect 30064 61140 30070 61192
rect 29917 61115 29975 61121
rect 29917 61112 29929 61115
rect 25832 61084 26372 61112
rect 27632 61084 27844 61112
rect 28966 61084 29929 61112
rect 25832 61072 25838 61084
rect 12713 61047 12771 61053
rect 12713 61044 12725 61047
rect 12584 61016 12725 61044
rect 12584 61004 12590 61016
rect 12713 61013 12725 61016
rect 12759 61013 12771 61047
rect 12713 61007 12771 61013
rect 16942 61004 16948 61056
rect 17000 61044 17006 61056
rect 17313 61047 17371 61053
rect 17313 61044 17325 61047
rect 17000 61016 17325 61044
rect 17000 61004 17006 61016
rect 17313 61013 17325 61016
rect 17359 61013 17371 61047
rect 17313 61007 17371 61013
rect 19702 61004 19708 61056
rect 19760 61044 19766 61056
rect 19797 61047 19855 61053
rect 19797 61044 19809 61047
rect 19760 61016 19809 61044
rect 19760 61004 19766 61016
rect 19797 61013 19809 61016
rect 19843 61013 19855 61047
rect 19797 61007 19855 61013
rect 23474 61004 23480 61056
rect 23532 61044 23538 61056
rect 23661 61047 23719 61053
rect 23661 61044 23673 61047
rect 23532 61016 23673 61044
rect 23532 61004 23538 61016
rect 23661 61013 23673 61016
rect 23707 61013 23719 61047
rect 23661 61007 23719 61013
rect 24578 61004 24584 61056
rect 24636 61044 24642 61056
rect 25314 61044 25320 61056
rect 24636 61016 25320 61044
rect 24636 61004 24642 61016
rect 25314 61004 25320 61016
rect 25372 61004 25378 61056
rect 25498 61004 25504 61056
rect 25556 61044 25562 61056
rect 25682 61044 25688 61056
rect 25556 61016 25688 61044
rect 25556 61004 25562 61016
rect 25682 61004 25688 61016
rect 25740 61004 25746 61056
rect 26234 61044 26240 61056
rect 26195 61016 26240 61044
rect 26234 61004 26240 61016
rect 26292 61004 26298 61056
rect 26344 61044 26372 61084
rect 28966 61044 28994 61084
rect 29917 61081 29929 61084
rect 29963 61081 29975 61115
rect 29917 61075 29975 61081
rect 26344 61016 28994 61044
rect 29086 61004 29092 61056
rect 29144 61044 29150 61056
rect 30098 61044 30104 61056
rect 29144 61016 30104 61044
rect 29144 61004 29150 61016
rect 30098 61004 30104 61016
rect 30156 61004 30162 61056
rect 1104 60954 30820 60976
rect 1104 60902 10880 60954
rect 10932 60902 10944 60954
rect 10996 60902 11008 60954
rect 11060 60902 11072 60954
rect 11124 60902 11136 60954
rect 11188 60902 20811 60954
rect 20863 60902 20875 60954
rect 20927 60902 20939 60954
rect 20991 60902 21003 60954
rect 21055 60902 21067 60954
rect 21119 60902 30820 60954
rect 1104 60880 30820 60902
rect 16114 60840 16120 60852
rect 13740 60812 16120 60840
rect 12526 60772 12532 60784
rect 12487 60744 12532 60772
rect 12526 60732 12532 60744
rect 12584 60732 12590 60784
rect 1578 60704 1584 60716
rect 1539 60676 1584 60704
rect 1578 60664 1584 60676
rect 1636 60664 1642 60716
rect 12713 60707 12771 60713
rect 12713 60704 12725 60707
rect 12406 60676 12725 60704
rect 11330 60596 11336 60648
rect 11388 60636 11394 60648
rect 12406 60636 12434 60676
rect 12713 60673 12725 60676
rect 12759 60673 12771 60707
rect 13630 60704 13636 60716
rect 13591 60676 13636 60704
rect 12713 60667 12771 60673
rect 13630 60664 13636 60676
rect 13688 60664 13694 60716
rect 13740 60713 13768 60812
rect 16114 60800 16120 60812
rect 16172 60800 16178 60852
rect 18322 60840 18328 60852
rect 18283 60812 18328 60840
rect 18322 60800 18328 60812
rect 18380 60800 18386 60852
rect 18782 60800 18788 60852
rect 18840 60840 18846 60852
rect 18877 60843 18935 60849
rect 18877 60840 18889 60843
rect 18840 60812 18889 60840
rect 18840 60800 18846 60812
rect 18877 60809 18889 60812
rect 18923 60809 18935 60843
rect 19702 60840 19708 60852
rect 18877 60803 18935 60809
rect 19257 60812 19708 60840
rect 17862 60732 17868 60784
rect 17920 60772 17926 60784
rect 18966 60772 18972 60784
rect 17920 60744 18972 60772
rect 17920 60732 17926 60744
rect 18966 60732 18972 60744
rect 19024 60732 19030 60784
rect 13725 60707 13783 60713
rect 13725 60673 13737 60707
rect 13771 60673 13783 60707
rect 13725 60667 13783 60673
rect 13817 60707 13875 60713
rect 13817 60673 13829 60707
rect 13863 60673 13875 60707
rect 13817 60667 13875 60673
rect 11388 60608 12434 60636
rect 13832 60636 13860 60667
rect 13998 60664 14004 60716
rect 14056 60704 14062 60716
rect 14717 60707 14775 60713
rect 14717 60704 14729 60707
rect 14056 60676 14101 60704
rect 14200 60676 14729 60704
rect 14056 60664 14062 60676
rect 13832 60608 14044 60636
rect 11388 60596 11394 60608
rect 14016 60580 14044 60608
rect 13998 60528 14004 60580
rect 14056 60528 14062 60580
rect 1397 60503 1455 60509
rect 1397 60469 1409 60503
rect 1443 60500 1455 60503
rect 12710 60500 12716 60512
rect 1443 60472 12716 60500
rect 1443 60469 1455 60472
rect 1397 60463 1455 60469
rect 12710 60460 12716 60472
rect 12768 60460 12774 60512
rect 12894 60500 12900 60512
rect 12855 60472 12900 60500
rect 12894 60460 12900 60472
rect 12952 60460 12958 60512
rect 13357 60503 13415 60509
rect 13357 60469 13369 60503
rect 13403 60500 13415 60503
rect 14200 60500 14228 60676
rect 14717 60673 14729 60676
rect 14763 60673 14775 60707
rect 14717 60667 14775 60673
rect 16666 60664 16672 60716
rect 16724 60704 16730 60716
rect 17201 60707 17259 60713
rect 17201 60704 17213 60707
rect 16724 60676 17213 60704
rect 16724 60664 16730 60676
rect 17201 60673 17213 60676
rect 17247 60673 17259 60707
rect 17201 60667 17259 60673
rect 19058 60664 19064 60716
rect 19116 60704 19122 60716
rect 19257 60713 19285 60812
rect 19702 60800 19708 60812
rect 19760 60800 19766 60852
rect 24118 60800 24124 60852
rect 24176 60840 24182 60852
rect 24670 60840 24676 60852
rect 24176 60812 24676 60840
rect 24176 60800 24182 60812
rect 24670 60800 24676 60812
rect 24728 60800 24734 60852
rect 25866 60800 25872 60852
rect 25924 60840 25930 60852
rect 26973 60843 27031 60849
rect 25924 60812 26464 60840
rect 25924 60800 25930 60812
rect 22002 60772 22008 60784
rect 21008 60744 22008 60772
rect 19153 60707 19211 60713
rect 19153 60704 19165 60707
rect 19116 60676 19165 60704
rect 19116 60664 19122 60676
rect 19153 60673 19165 60676
rect 19199 60673 19211 60707
rect 19153 60667 19211 60673
rect 19245 60707 19303 60713
rect 19245 60673 19257 60707
rect 19291 60673 19303 60707
rect 19245 60667 19303 60673
rect 19337 60707 19395 60713
rect 19337 60673 19349 60707
rect 19383 60673 19395 60707
rect 19337 60667 19395 60673
rect 19515 60707 19573 60713
rect 19515 60673 19527 60707
rect 19561 60702 19573 60707
rect 19610 60702 19616 60716
rect 19561 60674 19616 60702
rect 19561 60673 19573 60674
rect 19515 60667 19573 60673
rect 14274 60596 14280 60648
rect 14332 60636 14338 60648
rect 14461 60639 14519 60645
rect 14461 60636 14473 60639
rect 14332 60608 14473 60636
rect 14332 60596 14338 60608
rect 14461 60605 14473 60608
rect 14507 60605 14519 60639
rect 14461 60599 14519 60605
rect 16850 60596 16856 60648
rect 16908 60636 16914 60648
rect 16945 60639 17003 60645
rect 16945 60636 16957 60639
rect 16908 60608 16957 60636
rect 16908 60596 16914 60608
rect 16945 60605 16957 60608
rect 16991 60605 17003 60639
rect 16945 60599 17003 60605
rect 18414 60596 18420 60648
rect 18472 60636 18478 60648
rect 19352 60636 19380 60667
rect 19610 60664 19616 60674
rect 19668 60664 19674 60716
rect 20806 60664 20812 60716
rect 20864 60713 20870 60716
rect 21008 60713 21036 60744
rect 22002 60732 22008 60744
rect 22060 60732 22066 60784
rect 22646 60732 22652 60784
rect 22704 60772 22710 60784
rect 25041 60775 25099 60781
rect 25041 60772 25053 60775
rect 22704 60744 25053 60772
rect 22704 60732 22710 60744
rect 25041 60741 25053 60744
rect 25087 60741 25099 60775
rect 26436 60772 26464 60812
rect 26973 60809 26985 60843
rect 27019 60840 27031 60843
rect 27522 60840 27528 60852
rect 27019 60812 27528 60840
rect 27019 60809 27031 60812
rect 26973 60803 27031 60809
rect 27522 60800 27528 60812
rect 27580 60800 27586 60852
rect 27798 60800 27804 60852
rect 27856 60840 27862 60852
rect 27856 60812 28120 60840
rect 27856 60800 27862 60812
rect 27341 60775 27399 60781
rect 27341 60772 27353 60775
rect 25041 60735 25099 60741
rect 26068 60744 26372 60772
rect 26436 60744 27353 60772
rect 20864 60707 20913 60713
rect 20864 60673 20867 60707
rect 20901 60673 20913 60707
rect 20864 60667 20913 60673
rect 20993 60707 21051 60713
rect 20993 60673 21005 60707
rect 21039 60673 21051 60707
rect 20993 60667 21051 60673
rect 21085 60707 21143 60713
rect 21085 60673 21097 60707
rect 21131 60704 21143 60707
rect 21174 60704 21180 60716
rect 21131 60676 21180 60704
rect 21131 60673 21143 60676
rect 21085 60667 21143 60673
rect 20864 60664 20870 60667
rect 21174 60664 21180 60676
rect 21232 60664 21238 60716
rect 21281 60707 21339 60713
rect 21281 60673 21293 60707
rect 21327 60704 21339 60707
rect 21542 60704 21548 60716
rect 21327 60676 21548 60704
rect 21327 60673 21339 60676
rect 21281 60667 21339 60673
rect 21542 60664 21548 60676
rect 21600 60664 21606 60716
rect 22830 60704 22836 60716
rect 22791 60676 22836 60704
rect 22830 60664 22836 60676
rect 22888 60664 22894 60716
rect 23017 60707 23075 60713
rect 23017 60673 23029 60707
rect 23063 60704 23075 60707
rect 23106 60704 23112 60716
rect 23063 60676 23112 60704
rect 23063 60673 23075 60676
rect 23017 60667 23075 60673
rect 23106 60664 23112 60676
rect 23164 60704 23170 60716
rect 23937 60707 23995 60713
rect 23937 60704 23949 60707
rect 23164 60676 23949 60704
rect 23164 60664 23170 60676
rect 23937 60673 23949 60676
rect 23983 60673 23995 60707
rect 23937 60667 23995 60673
rect 24857 60707 24915 60713
rect 24857 60673 24869 60707
rect 24903 60704 24915 60707
rect 24946 60704 24952 60716
rect 24903 60676 24952 60704
rect 24903 60673 24915 60676
rect 24857 60667 24915 60673
rect 24946 60664 24952 60676
rect 25004 60664 25010 60716
rect 25133 60707 25191 60713
rect 25133 60673 25145 60707
rect 25179 60704 25191 60707
rect 25222 60704 25228 60716
rect 25179 60676 25228 60704
rect 25179 60673 25191 60676
rect 25133 60667 25191 60673
rect 25222 60664 25228 60676
rect 25280 60664 25286 60716
rect 25314 60664 25320 60716
rect 25372 60664 25378 60716
rect 25774 60670 25780 60722
rect 25832 60704 25838 60722
rect 25961 60707 26019 60713
rect 25961 60704 25973 60707
rect 25832 60676 25973 60704
rect 25832 60670 25838 60676
rect 25961 60673 25973 60676
rect 26007 60673 26019 60707
rect 25961 60667 26019 60673
rect 19794 60636 19800 60648
rect 18472 60608 19800 60636
rect 18472 60596 18478 60608
rect 19794 60596 19800 60608
rect 19852 60596 19858 60648
rect 23753 60639 23811 60645
rect 23753 60605 23765 60639
rect 23799 60605 23811 60639
rect 25332 60636 25360 60664
rect 25498 60636 25504 60648
rect 25332 60608 25504 60636
rect 23753 60599 23811 60605
rect 15396 60540 15976 60568
rect 13403 60472 14228 60500
rect 13403 60469 13415 60472
rect 13357 60463 13415 60469
rect 14734 60460 14740 60512
rect 14792 60500 14798 60512
rect 15396 60500 15424 60540
rect 14792 60472 15424 60500
rect 14792 60460 14798 60472
rect 15746 60460 15752 60512
rect 15804 60500 15810 60512
rect 15841 60503 15899 60509
rect 15841 60500 15853 60503
rect 15804 60472 15853 60500
rect 15804 60460 15810 60472
rect 15841 60469 15853 60472
rect 15887 60469 15899 60503
rect 15948 60500 15976 60540
rect 18690 60528 18696 60580
rect 18748 60568 18754 60580
rect 23768 60568 23796 60599
rect 25498 60596 25504 60608
rect 25556 60596 25562 60648
rect 26068 60636 26096 60744
rect 26344 60713 26372 60744
rect 27341 60741 27353 60744
rect 27387 60741 27399 60775
rect 27341 60735 27399 60741
rect 26145 60707 26203 60713
rect 26145 60673 26157 60707
rect 26191 60673 26203 60707
rect 26145 60667 26203 60673
rect 26329 60707 26387 60713
rect 26329 60673 26341 60707
rect 26375 60673 26387 60707
rect 26329 60667 26387 60673
rect 26421 60707 26479 60713
rect 26421 60673 26433 60707
rect 26467 60704 26479 60707
rect 27062 60704 27068 60716
rect 26467 60676 27068 60704
rect 26467 60673 26479 60676
rect 26421 60667 26479 60673
rect 25608 60608 26096 60636
rect 26160 60636 26188 60667
rect 27062 60664 27068 60676
rect 27120 60664 27126 60716
rect 27157 60707 27215 60713
rect 27157 60673 27169 60707
rect 27203 60673 27215 60707
rect 27430 60704 27436 60716
rect 27391 60676 27436 60704
rect 27157 60667 27215 60673
rect 26786 60636 26792 60648
rect 26160 60608 26792 60636
rect 18748 60540 23796 60568
rect 18748 60528 18754 60540
rect 24394 60528 24400 60580
rect 24452 60568 24458 60580
rect 25608 60568 25636 60608
rect 26786 60596 26792 60608
rect 26844 60636 26850 60648
rect 27172 60636 27200 60667
rect 27430 60664 27436 60676
rect 27488 60664 27494 60716
rect 28092 60713 28120 60812
rect 28626 60800 28632 60852
rect 28684 60840 28690 60852
rect 28684 60812 28994 60840
rect 28684 60800 28690 60812
rect 28966 60772 28994 60812
rect 29454 60772 29460 60784
rect 28966 60744 29460 60772
rect 29454 60732 29460 60744
rect 29512 60732 29518 60784
rect 29730 60772 29736 60784
rect 29691 60744 29736 60772
rect 29730 60732 29736 60744
rect 29788 60732 29794 60784
rect 28077 60707 28135 60713
rect 28077 60673 28089 60707
rect 28123 60704 28135 60707
rect 28902 60704 28908 60716
rect 28123 60676 28396 60704
rect 28863 60676 28908 60704
rect 28123 60673 28135 60676
rect 28077 60667 28135 60673
rect 27448 60636 27476 60664
rect 26844 60608 27200 60636
rect 27264 60608 27476 60636
rect 26844 60596 26850 60608
rect 26142 60568 26148 60580
rect 24452 60540 25636 60568
rect 25884 60540 26148 60568
rect 24452 60528 24458 60540
rect 19610 60500 19616 60512
rect 15948 60472 19616 60500
rect 15841 60463 15899 60469
rect 19610 60460 19616 60472
rect 19668 60460 19674 60512
rect 20622 60500 20628 60512
rect 20583 60472 20628 60500
rect 20622 60460 20628 60472
rect 20680 60460 20686 60512
rect 22094 60460 22100 60512
rect 22152 60500 22158 60512
rect 23201 60503 23259 60509
rect 23201 60500 23213 60503
rect 22152 60472 23213 60500
rect 22152 60460 22158 60472
rect 23201 60469 23213 60472
rect 23247 60469 23259 60503
rect 23201 60463 23259 60469
rect 23566 60460 23572 60512
rect 23624 60500 23630 60512
rect 24121 60503 24179 60509
rect 24121 60500 24133 60503
rect 23624 60472 24133 60500
rect 23624 60460 23630 60472
rect 24121 60469 24133 60472
rect 24167 60469 24179 60503
rect 24121 60463 24179 60469
rect 24673 60503 24731 60509
rect 24673 60469 24685 60503
rect 24719 60500 24731 60503
rect 25884 60500 25912 60540
rect 26142 60528 26148 60540
rect 26200 60528 26206 60580
rect 26326 60528 26332 60580
rect 26384 60568 26390 60580
rect 27062 60568 27068 60580
rect 26384 60540 27068 60568
rect 26384 60528 26390 60540
rect 27062 60528 27068 60540
rect 27120 60568 27126 60580
rect 27264 60568 27292 60608
rect 27120 60540 27292 60568
rect 27120 60528 27126 60540
rect 28368 60512 28396 60676
rect 28902 60664 28908 60676
rect 28960 60664 28966 60716
rect 29086 60664 29092 60716
rect 29144 60704 29150 60716
rect 29144 60676 29408 60704
rect 29144 60664 29150 60676
rect 29380 60648 29408 60676
rect 29362 60596 29368 60648
rect 29420 60596 29426 60648
rect 29454 60596 29460 60648
rect 29512 60636 29518 60648
rect 30926 60636 30932 60648
rect 29512 60608 30932 60636
rect 29512 60596 29518 60608
rect 30926 60596 30932 60608
rect 30984 60596 30990 60648
rect 24719 60472 25912 60500
rect 24719 60469 24731 60472
rect 24673 60463 24731 60469
rect 27338 60460 27344 60512
rect 27396 60500 27402 60512
rect 28169 60503 28227 60509
rect 28169 60500 28181 60503
rect 27396 60472 28181 60500
rect 27396 60460 27402 60472
rect 28169 60469 28181 60472
rect 28215 60469 28227 60503
rect 28169 60463 28227 60469
rect 28350 60460 28356 60512
rect 28408 60460 28414 60512
rect 29089 60503 29147 60509
rect 29089 60469 29101 60503
rect 29135 60500 29147 60503
rect 29730 60500 29736 60512
rect 29135 60472 29736 60500
rect 29135 60469 29147 60472
rect 29089 60463 29147 60469
rect 29730 60460 29736 60472
rect 29788 60460 29794 60512
rect 29822 60460 29828 60512
rect 29880 60500 29886 60512
rect 29880 60472 29925 60500
rect 29880 60460 29886 60472
rect 1104 60410 30820 60432
rect 1104 60358 5915 60410
rect 5967 60358 5979 60410
rect 6031 60358 6043 60410
rect 6095 60358 6107 60410
rect 6159 60358 6171 60410
rect 6223 60358 15846 60410
rect 15898 60358 15910 60410
rect 15962 60358 15974 60410
rect 16026 60358 16038 60410
rect 16090 60358 16102 60410
rect 16154 60358 25776 60410
rect 25828 60358 25840 60410
rect 25892 60358 25904 60410
rect 25956 60358 25968 60410
rect 26020 60358 26032 60410
rect 26084 60358 30820 60410
rect 1104 60336 30820 60358
rect 13630 60256 13636 60308
rect 13688 60296 13694 60308
rect 15746 60296 15752 60308
rect 13688 60268 15752 60296
rect 13688 60256 13694 60268
rect 15746 60256 15752 60268
rect 15804 60256 15810 60308
rect 17310 60256 17316 60308
rect 17368 60296 17374 60308
rect 17865 60299 17923 60305
rect 17865 60296 17877 60299
rect 17368 60268 17877 60296
rect 17368 60256 17374 60268
rect 17865 60265 17877 60268
rect 17911 60265 17923 60299
rect 17865 60259 17923 60265
rect 21726 60256 21732 60308
rect 21784 60296 21790 60308
rect 22370 60296 22376 60308
rect 21784 60268 22094 60296
rect 22331 60268 22376 60296
rect 21784 60256 21790 60268
rect 14090 60188 14096 60240
rect 14148 60228 14154 60240
rect 14185 60231 14243 60237
rect 14185 60228 14197 60231
rect 14148 60200 14197 60228
rect 14148 60188 14154 60200
rect 14185 60197 14197 60200
rect 14231 60197 14243 60231
rect 14185 60191 14243 60197
rect 12897 60163 12955 60169
rect 12897 60129 12909 60163
rect 12943 60160 12955 60163
rect 19334 60160 19340 60172
rect 12943 60132 19340 60160
rect 12943 60129 12955 60132
rect 12897 60123 12955 60129
rect 19334 60120 19340 60132
rect 19392 60120 19398 60172
rect 20346 60120 20352 60172
rect 20404 60160 20410 60172
rect 20530 60160 20536 60172
rect 20404 60132 20536 60160
rect 20404 60120 20410 60132
rect 20530 60120 20536 60132
rect 20588 60120 20594 60172
rect 22066 60160 22094 60268
rect 22370 60256 22376 60268
rect 22428 60256 22434 60308
rect 23934 60256 23940 60308
rect 23992 60296 23998 60308
rect 25314 60296 25320 60308
rect 23992 60268 25320 60296
rect 23992 60256 23998 60268
rect 25314 60256 25320 60268
rect 25372 60256 25378 60308
rect 25593 60299 25651 60305
rect 25593 60265 25605 60299
rect 25639 60296 25651 60299
rect 26602 60296 26608 60308
rect 25639 60268 26608 60296
rect 25639 60265 25651 60268
rect 25593 60259 25651 60265
rect 26602 60256 26608 60268
rect 26660 60256 26666 60308
rect 26694 60256 26700 60308
rect 26752 60296 26758 60308
rect 28537 60299 28595 60305
rect 28537 60296 28549 60299
rect 26752 60268 28549 60296
rect 26752 60256 26758 60268
rect 28537 60265 28549 60268
rect 28583 60265 28595 60299
rect 28537 60259 28595 60265
rect 23474 60188 23480 60240
rect 23532 60228 23538 60240
rect 23532 60200 25728 60228
rect 23532 60188 23538 60200
rect 22925 60163 22983 60169
rect 22925 60160 22937 60163
rect 22066 60132 22937 60160
rect 22925 60129 22937 60132
rect 22971 60129 22983 60163
rect 25700 60160 25728 60200
rect 27154 60188 27160 60240
rect 27212 60228 27218 60240
rect 27433 60231 27491 60237
rect 27433 60228 27445 60231
rect 27212 60200 27445 60228
rect 27212 60188 27218 60200
rect 27433 60197 27445 60200
rect 27479 60197 27491 60231
rect 27433 60191 27491 60197
rect 27540 60200 28120 60228
rect 25866 60160 25872 60172
rect 25700 60132 25872 60160
rect 22925 60123 22983 60129
rect 25866 60120 25872 60132
rect 25924 60160 25930 60172
rect 27540 60160 27568 60200
rect 28092 60169 28120 60200
rect 28077 60163 28135 60169
rect 25924 60132 27568 60160
rect 27632 60132 28028 60160
rect 25924 60120 25930 60132
rect 1578 60092 1584 60104
rect 1539 60064 1584 60092
rect 1578 60052 1584 60064
rect 1636 60052 1642 60104
rect 11238 60052 11244 60104
rect 11296 60092 11302 60104
rect 11296 60064 12434 60092
rect 11296 60052 11302 60064
rect 12406 60024 12434 60064
rect 12526 60052 12532 60104
rect 12584 60092 12590 60104
rect 17678 60092 17684 60104
rect 12584 60064 12629 60092
rect 17639 60064 17684 60092
rect 12584 60052 12590 60064
rect 17678 60052 17684 60064
rect 17736 60052 17742 60104
rect 19475 60095 19533 60101
rect 19475 60061 19487 60095
rect 19521 60061 19533 60095
rect 19610 60092 19616 60104
rect 19571 60064 19616 60092
rect 19475 60055 19533 60061
rect 12713 60027 12771 60033
rect 12713 60024 12725 60027
rect 12406 59996 12725 60024
rect 12713 59993 12725 59996
rect 12759 59993 12771 60027
rect 14458 60024 14464 60036
rect 14419 59996 14464 60024
rect 12713 59987 12771 59993
rect 14458 59984 14464 59996
rect 14516 59984 14522 60036
rect 14642 60024 14648 60036
rect 14603 59996 14648 60024
rect 14642 59984 14648 59996
rect 14700 59984 14706 60036
rect 14734 59984 14740 60036
rect 14792 60024 14798 60036
rect 15470 60024 15476 60036
rect 14792 59996 14837 60024
rect 15431 59996 15476 60024
rect 14792 59984 14798 59996
rect 15470 59984 15476 59996
rect 15528 59984 15534 60036
rect 15746 59984 15752 60036
rect 15804 60024 15810 60036
rect 18966 60024 18972 60036
rect 15804 59996 18972 60024
rect 15804 59984 15810 59996
rect 18966 59984 18972 59996
rect 19024 59984 19030 60036
rect 19490 60024 19518 60055
rect 19610 60052 19616 60064
rect 19668 60052 19674 60104
rect 19705 60095 19763 60101
rect 19705 60061 19717 60095
rect 19751 60092 19763 60095
rect 19794 60092 19800 60104
rect 19751 60064 19800 60092
rect 19751 60061 19763 60064
rect 19705 60055 19763 60061
rect 19794 60052 19800 60064
rect 19852 60052 19858 60104
rect 19886 60052 19892 60104
rect 19944 60092 19950 60104
rect 20993 60095 21051 60101
rect 19944 60064 19989 60092
rect 19944 60052 19950 60064
rect 20993 60061 21005 60095
rect 21039 60092 21051 60095
rect 23109 60095 23167 60101
rect 21039 60064 21496 60092
rect 21039 60061 21051 60064
rect 20993 60055 21051 60061
rect 21468 60036 21496 60064
rect 23109 60061 23121 60095
rect 23155 60092 23167 60095
rect 23198 60092 23204 60104
rect 23155 60064 23204 60092
rect 23155 60061 23167 60064
rect 23109 60055 23167 60061
rect 23198 60052 23204 60064
rect 23256 60052 23262 60104
rect 25774 60092 25780 60104
rect 25735 60064 25780 60092
rect 25774 60052 25780 60064
rect 25832 60052 25838 60104
rect 26053 60095 26111 60101
rect 26053 60061 26065 60095
rect 26099 60092 26111 60095
rect 26326 60092 26332 60104
rect 26099 60064 26332 60092
rect 26099 60061 26111 60064
rect 26053 60055 26111 60061
rect 26326 60052 26332 60064
rect 26384 60052 26390 60104
rect 26602 60052 26608 60104
rect 26660 60092 26666 60104
rect 26881 60095 26939 60101
rect 26881 60092 26893 60095
rect 26660 60064 26893 60092
rect 26660 60052 26666 60064
rect 26881 60061 26893 60064
rect 26927 60061 26939 60095
rect 26881 60055 26939 60061
rect 27154 60052 27160 60104
rect 27212 60092 27218 60104
rect 27632 60092 27660 60132
rect 27798 60092 27804 60104
rect 27212 60064 27660 60092
rect 27759 60064 27804 60092
rect 27212 60052 27218 60064
rect 27798 60052 27804 60064
rect 27856 60052 27862 60104
rect 28000 60101 28028 60132
rect 28077 60129 28089 60163
rect 28123 60129 28135 60163
rect 28077 60123 28135 60129
rect 27985 60095 28043 60101
rect 27985 60061 27997 60095
rect 28031 60061 28043 60095
rect 27985 60055 28043 60061
rect 28169 60095 28227 60101
rect 28169 60061 28181 60095
rect 28215 60061 28227 60095
rect 28350 60092 28356 60104
rect 28311 60064 28356 60092
rect 28169 60055 28227 60061
rect 20530 60024 20536 60036
rect 19490 59996 20536 60024
rect 20530 59984 20536 59996
rect 20588 59984 20594 60036
rect 20622 59984 20628 60036
rect 20680 60024 20686 60036
rect 21238 60027 21296 60033
rect 21238 60024 21250 60027
rect 20680 59996 21250 60024
rect 20680 59984 20686 59996
rect 21238 59993 21250 59996
rect 21284 59993 21296 60027
rect 21238 59987 21296 59993
rect 21450 59984 21456 60036
rect 21508 59984 21514 60036
rect 21910 59984 21916 60036
rect 21968 60024 21974 60036
rect 25961 60027 26019 60033
rect 25961 60024 25973 60027
rect 21968 59996 25973 60024
rect 21968 59984 21974 59996
rect 25961 59993 25973 59996
rect 26007 59993 26019 60027
rect 25961 59987 26019 59993
rect 28074 59984 28080 60036
rect 28132 60024 28138 60036
rect 28184 60024 28212 60055
rect 28350 60052 28356 60064
rect 28408 60052 28414 60104
rect 29825 60095 29883 60101
rect 29825 60061 29837 60095
rect 29871 60092 29883 60095
rect 29914 60092 29920 60104
rect 29871 60064 29920 60092
rect 29871 60061 29883 60064
rect 29825 60055 29883 60061
rect 29914 60052 29920 60064
rect 29972 60052 29978 60104
rect 28132 59996 28212 60024
rect 28132 59984 28138 59996
rect 1397 59959 1455 59965
rect 1397 59925 1409 59959
rect 1443 59956 1455 59959
rect 11330 59956 11336 59968
rect 1443 59928 11336 59956
rect 1443 59925 1455 59928
rect 1397 59919 1455 59925
rect 11330 59916 11336 59928
rect 11388 59916 11394 59968
rect 16666 59916 16672 59968
rect 16724 59956 16730 59968
rect 16761 59959 16819 59965
rect 16761 59956 16773 59959
rect 16724 59928 16773 59956
rect 16724 59916 16730 59928
rect 16761 59925 16773 59928
rect 16807 59925 16819 59959
rect 16761 59919 16819 59925
rect 19150 59916 19156 59968
rect 19208 59956 19214 59968
rect 19245 59959 19303 59965
rect 19245 59956 19257 59959
rect 19208 59928 19257 59956
rect 19208 59916 19214 59928
rect 19245 59925 19257 59928
rect 19291 59925 19303 59959
rect 23290 59956 23296 59968
rect 23251 59928 23296 59956
rect 19245 59919 19303 59925
rect 23290 59916 23296 59928
rect 23348 59916 23354 59968
rect 26602 59916 26608 59968
rect 26660 59956 26666 59968
rect 26786 59956 26792 59968
rect 26660 59928 26792 59956
rect 26660 59916 26666 59928
rect 26786 59916 26792 59928
rect 26844 59956 26850 59968
rect 27065 59959 27123 59965
rect 27065 59956 27077 59959
rect 26844 59928 27077 59956
rect 26844 59916 26850 59928
rect 27065 59925 27077 59928
rect 27111 59925 27123 59959
rect 27065 59919 27123 59925
rect 28350 59916 28356 59968
rect 28408 59956 28414 59968
rect 28626 59956 28632 59968
rect 28408 59928 28632 59956
rect 28408 59916 28414 59928
rect 28626 59916 28632 59928
rect 28684 59916 28690 59968
rect 29454 59916 29460 59968
rect 29512 59956 29518 59968
rect 30009 59959 30067 59965
rect 30009 59956 30021 59959
rect 29512 59928 30021 59956
rect 29512 59916 29518 59928
rect 30009 59925 30021 59928
rect 30055 59925 30067 59959
rect 30009 59919 30067 59925
rect 1104 59866 30820 59888
rect 1104 59814 10880 59866
rect 10932 59814 10944 59866
rect 10996 59814 11008 59866
rect 11060 59814 11072 59866
rect 11124 59814 11136 59866
rect 11188 59814 20811 59866
rect 20863 59814 20875 59866
rect 20927 59814 20939 59866
rect 20991 59814 21003 59866
rect 21055 59814 21067 59866
rect 21119 59814 30820 59866
rect 1104 59792 30820 59814
rect 13538 59752 13544 59764
rect 13499 59724 13544 59752
rect 13538 59712 13544 59724
rect 13596 59712 13602 59764
rect 14274 59752 14280 59764
rect 14235 59724 14280 59752
rect 14274 59712 14280 59724
rect 14332 59712 14338 59764
rect 16850 59752 16856 59764
rect 16811 59724 16856 59752
rect 16850 59712 16856 59724
rect 16908 59712 16914 59764
rect 23845 59755 23903 59761
rect 23845 59752 23857 59755
rect 16960 59724 19656 59752
rect 12526 59684 12532 59696
rect 12487 59656 12532 59684
rect 12526 59644 12532 59656
rect 12584 59644 12590 59696
rect 12710 59684 12716 59696
rect 12671 59656 12716 59684
rect 12710 59644 12716 59656
rect 12768 59644 12774 59696
rect 16298 59644 16304 59696
rect 16356 59684 16362 59696
rect 16960 59684 16988 59724
rect 16356 59656 16988 59684
rect 16356 59644 16362 59656
rect 19150 59644 19156 59696
rect 19208 59684 19214 59696
rect 19512 59687 19570 59693
rect 19512 59684 19524 59687
rect 19208 59656 19524 59684
rect 19208 59644 19214 59656
rect 19512 59653 19524 59656
rect 19558 59653 19570 59687
rect 19628 59684 19656 59724
rect 23124 59724 23857 59752
rect 19628 59656 22094 59684
rect 19512 59647 19570 59653
rect 1578 59616 1584 59628
rect 1539 59588 1584 59616
rect 1578 59576 1584 59588
rect 1636 59576 1642 59628
rect 13446 59616 13452 59628
rect 13407 59588 13452 59616
rect 13446 59576 13452 59588
rect 13504 59576 13510 59628
rect 14090 59616 14096 59628
rect 14051 59588 14096 59616
rect 14090 59576 14096 59588
rect 14148 59576 14154 59628
rect 16669 59619 16727 59625
rect 16669 59585 16681 59619
rect 16715 59616 16727 59619
rect 16758 59616 16764 59628
rect 16715 59588 16764 59616
rect 16715 59585 16727 59588
rect 16669 59579 16727 59585
rect 16758 59576 16764 59588
rect 16816 59576 16822 59628
rect 19058 59576 19064 59628
rect 19116 59616 19122 59628
rect 19245 59619 19303 59625
rect 19245 59616 19257 59619
rect 19116 59588 19257 59616
rect 19116 59576 19122 59588
rect 19245 59585 19257 59588
rect 19291 59585 19303 59619
rect 19886 59616 19892 59628
rect 19245 59579 19303 59585
rect 19352 59588 19892 59616
rect 12894 59508 12900 59560
rect 12952 59548 12958 59560
rect 19352 59548 19380 59588
rect 19886 59576 19892 59588
rect 19944 59576 19950 59628
rect 22066 59616 22094 59656
rect 23124 59628 23152 59724
rect 23845 59721 23857 59724
rect 23891 59721 23903 59755
rect 25777 59755 25835 59761
rect 25777 59752 25789 59755
rect 23845 59715 23903 59721
rect 24136 59724 25789 59752
rect 22925 59619 22983 59625
rect 22925 59616 22937 59619
rect 22066 59588 22937 59616
rect 22925 59585 22937 59588
rect 22971 59585 22983 59619
rect 23106 59616 23112 59628
rect 23067 59588 23112 59616
rect 22925 59579 22983 59585
rect 23106 59576 23112 59588
rect 23164 59576 23170 59628
rect 23934 59576 23940 59628
rect 23992 59616 23998 59628
rect 24029 59619 24087 59625
rect 24029 59616 24041 59619
rect 23992 59588 24041 59616
rect 23992 59576 23998 59588
rect 24029 59585 24041 59588
rect 24075 59585 24087 59619
rect 24029 59579 24087 59585
rect 12952 59520 19380 59548
rect 12952 59508 12958 59520
rect 23014 59508 23020 59560
rect 23072 59548 23078 59560
rect 23474 59548 23480 59560
rect 23072 59520 23480 59548
rect 23072 59508 23078 59520
rect 23474 59508 23480 59520
rect 23532 59508 23538 59560
rect 18874 59480 18880 59492
rect 12912 59452 18880 59480
rect 1397 59415 1455 59421
rect 1397 59381 1409 59415
rect 1443 59412 1455 59415
rect 11238 59412 11244 59424
rect 1443 59384 11244 59412
rect 1443 59381 1455 59384
rect 1397 59375 1455 59381
rect 11238 59372 11244 59384
rect 11296 59372 11302 59424
rect 12912 59421 12940 59452
rect 18874 59440 18880 59452
rect 18932 59440 18938 59492
rect 20530 59440 20536 59492
rect 20588 59480 20594 59492
rect 20625 59483 20683 59489
rect 20625 59480 20637 59483
rect 20588 59452 20637 59480
rect 20588 59440 20594 59452
rect 20625 59449 20637 59452
rect 20671 59480 20683 59483
rect 24136 59480 24164 59724
rect 25777 59721 25789 59724
rect 25823 59752 25835 59755
rect 25866 59752 25872 59764
rect 25823 59724 25872 59752
rect 25823 59721 25835 59724
rect 25777 59715 25835 59721
rect 25866 59712 25872 59724
rect 25924 59712 25930 59764
rect 26878 59712 26884 59764
rect 26936 59752 26942 59764
rect 27433 59755 27491 59761
rect 27433 59752 27445 59755
rect 26936 59724 27445 59752
rect 26936 59712 26942 59724
rect 27433 59721 27445 59724
rect 27479 59721 27491 59755
rect 27433 59715 27491 59721
rect 25222 59644 25228 59696
rect 25280 59684 25286 59696
rect 31018 59684 31024 59696
rect 25280 59656 25912 59684
rect 25280 59644 25286 59656
rect 25884 59625 25912 59656
rect 27816 59656 31024 59684
rect 25593 59619 25651 59625
rect 25593 59585 25605 59619
rect 25639 59585 25651 59619
rect 25593 59579 25651 59585
rect 25869 59619 25927 59625
rect 25869 59585 25881 59619
rect 25915 59585 25927 59619
rect 26326 59616 26332 59628
rect 25869 59579 25927 59585
rect 25976 59588 26332 59616
rect 25608 59548 25636 59579
rect 25976 59548 26004 59588
rect 26326 59576 26332 59588
rect 26384 59616 26390 59628
rect 27154 59616 27160 59628
rect 26384 59588 27160 59616
rect 26384 59576 26390 59588
rect 27154 59576 27160 59588
rect 27212 59576 27218 59628
rect 27338 59576 27344 59628
rect 27396 59616 27402 59628
rect 27706 59616 27712 59628
rect 27396 59588 27712 59616
rect 27396 59576 27402 59588
rect 27706 59576 27712 59588
rect 27764 59576 27770 59628
rect 27816 59625 27844 59656
rect 31018 59644 31024 59656
rect 31076 59644 31082 59696
rect 27801 59619 27859 59625
rect 27801 59585 27813 59619
rect 27847 59585 27859 59619
rect 27801 59579 27859 59585
rect 27893 59619 27951 59625
rect 27893 59585 27905 59619
rect 27939 59585 27951 59619
rect 28074 59616 28080 59628
rect 28035 59588 28080 59616
rect 27893 59579 27951 59585
rect 25608 59520 26004 59548
rect 26878 59508 26884 59560
rect 26936 59548 26942 59560
rect 27908 59548 27936 59579
rect 28074 59576 28080 59588
rect 28132 59576 28138 59628
rect 28905 59619 28963 59625
rect 28905 59616 28917 59619
rect 28736 59588 28917 59616
rect 28736 59560 28764 59588
rect 28905 59585 28917 59588
rect 28951 59585 28963 59619
rect 28905 59579 28963 59585
rect 29733 59619 29791 59625
rect 29733 59585 29745 59619
rect 29779 59616 29791 59619
rect 29822 59616 29828 59628
rect 29779 59588 29828 59616
rect 29779 59585 29791 59588
rect 29733 59579 29791 59585
rect 29822 59576 29828 59588
rect 29880 59576 29886 59628
rect 26936 59520 27936 59548
rect 26936 59508 26942 59520
rect 28718 59508 28724 59560
rect 28776 59508 28782 59560
rect 20671 59452 24164 59480
rect 20671 59449 20683 59452
rect 20625 59443 20683 59449
rect 25222 59440 25228 59492
rect 25280 59480 25286 59492
rect 25774 59480 25780 59492
rect 25280 59452 25780 59480
rect 25280 59440 25286 59452
rect 25774 59440 25780 59452
rect 25832 59440 25838 59492
rect 26970 59440 26976 59492
rect 27028 59480 27034 59492
rect 29089 59483 29147 59489
rect 27028 59452 27476 59480
rect 27028 59440 27034 59452
rect 12897 59415 12955 59421
rect 12897 59381 12909 59415
rect 12943 59381 12955 59415
rect 12897 59375 12955 59381
rect 14826 59372 14832 59424
rect 14884 59412 14890 59424
rect 21726 59412 21732 59424
rect 14884 59384 21732 59412
rect 14884 59372 14890 59384
rect 21726 59372 21732 59384
rect 21784 59372 21790 59424
rect 23198 59372 23204 59424
rect 23256 59412 23262 59424
rect 23293 59415 23351 59421
rect 23293 59412 23305 59415
rect 23256 59384 23305 59412
rect 23256 59372 23262 59384
rect 23293 59381 23305 59384
rect 23339 59381 23351 59415
rect 23293 59375 23351 59381
rect 25409 59415 25467 59421
rect 25409 59381 25421 59415
rect 25455 59412 25467 59415
rect 27338 59412 27344 59424
rect 25455 59384 27344 59412
rect 25455 59381 25467 59384
rect 25409 59375 25467 59381
rect 27338 59372 27344 59384
rect 27396 59372 27402 59424
rect 27448 59412 27476 59452
rect 29089 59449 29101 59483
rect 29135 59480 29147 59483
rect 30742 59480 30748 59492
rect 29135 59452 30748 59480
rect 29135 59449 29147 59452
rect 29089 59443 29147 59449
rect 30742 59440 30748 59452
rect 30800 59440 30806 59492
rect 29825 59415 29883 59421
rect 29825 59412 29837 59415
rect 27448 59384 29837 59412
rect 29825 59381 29837 59384
rect 29871 59381 29883 59415
rect 29825 59375 29883 59381
rect 1104 59322 30820 59344
rect 1104 59270 5915 59322
rect 5967 59270 5979 59322
rect 6031 59270 6043 59322
rect 6095 59270 6107 59322
rect 6159 59270 6171 59322
rect 6223 59270 15846 59322
rect 15898 59270 15910 59322
rect 15962 59270 15974 59322
rect 16026 59270 16038 59322
rect 16090 59270 16102 59322
rect 16154 59270 25776 59322
rect 25828 59270 25840 59322
rect 25892 59270 25904 59322
rect 25956 59270 25968 59322
rect 26020 59270 26032 59322
rect 26084 59270 30820 59322
rect 1104 59248 30820 59270
rect 18598 59168 18604 59220
rect 18656 59208 18662 59220
rect 19797 59211 19855 59217
rect 19797 59208 19809 59211
rect 18656 59180 19809 59208
rect 18656 59168 18662 59180
rect 19797 59177 19809 59180
rect 19843 59177 19855 59211
rect 19797 59171 19855 59177
rect 20254 59168 20260 59220
rect 20312 59208 20318 59220
rect 20530 59208 20536 59220
rect 20312 59180 20536 59208
rect 20312 59168 20318 59180
rect 20530 59168 20536 59180
rect 20588 59168 20594 59220
rect 20809 59211 20867 59217
rect 20809 59177 20821 59211
rect 20855 59208 20867 59211
rect 21358 59208 21364 59220
rect 20855 59180 21364 59208
rect 20855 59177 20867 59180
rect 20809 59171 20867 59177
rect 21358 59168 21364 59180
rect 21416 59168 21422 59220
rect 23382 59168 23388 59220
rect 23440 59208 23446 59220
rect 23440 59180 27936 59208
rect 23440 59168 23446 59180
rect 13541 59143 13599 59149
rect 13541 59109 13553 59143
rect 13587 59140 13599 59143
rect 21818 59140 21824 59152
rect 13587 59112 21824 59140
rect 13587 59109 13599 59112
rect 13541 59103 13599 59109
rect 21818 59100 21824 59112
rect 21876 59100 21882 59152
rect 27908 59140 27936 59180
rect 28626 59168 28632 59220
rect 28684 59208 28690 59220
rect 28721 59211 28779 59217
rect 28721 59208 28733 59211
rect 28684 59180 28733 59208
rect 28684 59168 28690 59180
rect 28721 59177 28733 59180
rect 28767 59177 28779 59211
rect 28721 59171 28779 59177
rect 29730 59168 29736 59220
rect 29788 59208 29794 59220
rect 30374 59208 30380 59220
rect 29788 59180 30380 59208
rect 29788 59168 29794 59180
rect 30374 59168 30380 59180
rect 30432 59168 30438 59220
rect 30650 59140 30656 59152
rect 27908 59112 30656 59140
rect 30650 59100 30656 59112
rect 30708 59100 30714 59152
rect 27157 59075 27215 59081
rect 27157 59041 27169 59075
rect 27203 59072 27215 59075
rect 27430 59072 27436 59084
rect 27203 59044 27436 59072
rect 27203 59041 27215 59044
rect 27157 59035 27215 59041
rect 27430 59032 27436 59044
rect 27488 59032 27494 59084
rect 11330 58964 11336 59016
rect 11388 59004 11394 59016
rect 13357 59007 13415 59013
rect 13357 59004 13369 59007
rect 11388 58976 13369 59004
rect 11388 58964 11394 58976
rect 13357 58973 13369 58976
rect 13403 58973 13415 59007
rect 13357 58967 13415 58973
rect 13538 58964 13544 59016
rect 13596 58964 13602 59016
rect 14645 59007 14703 59013
rect 14645 58973 14657 59007
rect 14691 59004 14703 59007
rect 16390 59004 16396 59016
rect 14691 58976 16396 59004
rect 14691 58973 14703 58976
rect 14645 58967 14703 58973
rect 16390 58964 16396 58976
rect 16448 58964 16454 59016
rect 20530 58964 20536 59016
rect 20588 59004 20594 59016
rect 20625 59007 20683 59013
rect 20625 59004 20637 59007
rect 20588 58976 20637 59004
rect 20588 58964 20594 58976
rect 20625 58973 20637 58976
rect 20671 58973 20683 59007
rect 20625 58967 20683 58973
rect 26881 59007 26939 59013
rect 26881 58973 26893 59007
rect 26927 59004 26939 59007
rect 26927 58976 27476 59004
rect 26927 58973 26939 58976
rect 26881 58967 26939 58973
rect 13170 58936 13176 58948
rect 13083 58908 13176 58936
rect 13170 58896 13176 58908
rect 13228 58936 13234 58948
rect 13556 58936 13584 58964
rect 27448 58948 27476 58976
rect 29362 58964 29368 59016
rect 29420 59004 29426 59016
rect 29420 58976 30144 59004
rect 29420 58964 29426 58976
rect 30116 58948 30144 58976
rect 13228 58908 13584 58936
rect 17865 58939 17923 58945
rect 13228 58896 13234 58908
rect 17865 58905 17877 58939
rect 17911 58936 17923 58939
rect 18322 58936 18328 58948
rect 17911 58908 18328 58936
rect 17911 58905 17923 58908
rect 17865 58899 17923 58905
rect 18322 58896 18328 58908
rect 18380 58896 18386 58948
rect 19705 58939 19763 58945
rect 19705 58905 19717 58939
rect 19751 58936 19763 58939
rect 20162 58936 20168 58948
rect 19751 58908 20168 58936
rect 19751 58905 19763 58908
rect 19705 58899 19763 58905
rect 20162 58896 20168 58908
rect 20220 58896 20226 58948
rect 23842 58896 23848 58948
rect 23900 58936 23906 58948
rect 24394 58936 24400 58948
rect 23900 58908 24400 58936
rect 23900 58896 23906 58908
rect 24394 58896 24400 58908
rect 24452 58896 24458 58948
rect 27430 58896 27436 58948
rect 27488 58896 27494 58948
rect 28626 58936 28632 58948
rect 28587 58908 28632 58936
rect 28626 58896 28632 58908
rect 28684 58896 28690 58948
rect 29730 58936 29736 58948
rect 29691 58908 29736 58936
rect 29730 58896 29736 58908
rect 29788 58896 29794 58948
rect 30098 58936 30104 58948
rect 30059 58908 30104 58936
rect 30098 58896 30104 58908
rect 30156 58896 30162 58948
rect 14458 58828 14464 58880
rect 14516 58868 14522 58880
rect 14737 58871 14795 58877
rect 14737 58868 14749 58871
rect 14516 58840 14749 58868
rect 14516 58828 14522 58840
rect 14737 58837 14749 58840
rect 14783 58837 14795 58871
rect 14737 58831 14795 58837
rect 17218 58828 17224 58880
rect 17276 58868 17282 58880
rect 17957 58871 18015 58877
rect 17957 58868 17969 58871
rect 17276 58840 17969 58868
rect 17276 58828 17282 58840
rect 17957 58837 17969 58840
rect 18003 58837 18015 58871
rect 17957 58831 18015 58837
rect 1104 58778 30820 58800
rect 1104 58726 10880 58778
rect 10932 58726 10944 58778
rect 10996 58726 11008 58778
rect 11060 58726 11072 58778
rect 11124 58726 11136 58778
rect 11188 58726 20811 58778
rect 20863 58726 20875 58778
rect 20927 58726 20939 58778
rect 20991 58726 21003 58778
rect 21055 58726 21067 58778
rect 21119 58726 30820 58778
rect 1104 58704 30820 58726
rect 19150 58624 19156 58676
rect 19208 58664 19214 58676
rect 19705 58667 19763 58673
rect 19705 58664 19717 58667
rect 19208 58636 19717 58664
rect 19208 58624 19214 58636
rect 19705 58633 19717 58636
rect 19751 58633 19763 58667
rect 19705 58627 19763 58633
rect 27433 58667 27491 58673
rect 27433 58633 27445 58667
rect 27479 58664 27491 58667
rect 27614 58664 27620 58676
rect 27479 58636 27620 58664
rect 27479 58633 27491 58636
rect 27433 58627 27491 58633
rect 27614 58624 27620 58636
rect 27672 58624 27678 58676
rect 27706 58624 27712 58676
rect 27764 58624 27770 58676
rect 28626 58664 28632 58676
rect 27816 58636 28632 58664
rect 11238 58556 11244 58608
rect 11296 58596 11302 58608
rect 13357 58599 13415 58605
rect 13357 58596 13369 58599
rect 11296 58568 13369 58596
rect 11296 58556 11302 58568
rect 13357 58565 13369 58568
rect 13403 58565 13415 58599
rect 13357 58559 13415 58565
rect 15933 58599 15991 58605
rect 15933 58565 15945 58599
rect 15979 58596 15991 58599
rect 16666 58596 16672 58608
rect 15979 58568 16672 58596
rect 15979 58565 15991 58568
rect 15933 58559 15991 58565
rect 16666 58556 16672 58568
rect 16724 58556 16730 58608
rect 17221 58599 17279 58605
rect 17221 58565 17233 58599
rect 17267 58596 17279 58599
rect 17586 58596 17592 58608
rect 17267 58568 17592 58596
rect 17267 58565 17279 58568
rect 17221 58559 17279 58565
rect 17586 58556 17592 58568
rect 17644 58556 17650 58608
rect 19061 58599 19119 58605
rect 19061 58565 19073 58599
rect 19107 58596 19119 58599
rect 19242 58596 19248 58608
rect 19107 58568 19248 58596
rect 19107 58565 19119 58568
rect 19061 58559 19119 58565
rect 19242 58556 19248 58568
rect 19300 58556 19306 58608
rect 20809 58599 20867 58605
rect 20809 58565 20821 58599
rect 20855 58596 20867 58599
rect 21174 58596 21180 58608
rect 20855 58568 21180 58596
rect 20855 58565 20867 58568
rect 20809 58559 20867 58565
rect 21174 58556 21180 58568
rect 21232 58596 21238 58608
rect 21634 58596 21640 58608
rect 21232 58568 21640 58596
rect 21232 58556 21238 58568
rect 21634 58556 21640 58568
rect 21692 58556 21698 58608
rect 26237 58599 26295 58605
rect 26237 58565 26249 58599
rect 26283 58596 26295 58599
rect 26326 58596 26332 58608
rect 26283 58568 26332 58596
rect 26283 58565 26295 58568
rect 26237 58559 26295 58565
rect 26326 58556 26332 58568
rect 26384 58556 26390 58608
rect 1394 58528 1400 58540
rect 1355 58500 1400 58528
rect 1394 58488 1400 58500
rect 1452 58488 1458 58540
rect 13170 58528 13176 58540
rect 13131 58500 13176 58528
rect 13170 58488 13176 58500
rect 13228 58488 13234 58540
rect 18877 58531 18935 58537
rect 18877 58497 18889 58531
rect 18923 58497 18935 58531
rect 19518 58528 19524 58540
rect 19479 58500 19524 58528
rect 18877 58491 18935 58497
rect 17218 58460 17224 58472
rect 17179 58432 17224 58460
rect 17218 58420 17224 58432
rect 17276 58420 17282 58472
rect 17310 58420 17316 58472
rect 17368 58460 17374 58472
rect 18892 58460 18920 58491
rect 19518 58488 19524 58500
rect 19576 58488 19582 58540
rect 20070 58488 20076 58540
rect 20128 58528 20134 58540
rect 20346 58528 20352 58540
rect 20128 58500 20352 58528
rect 20128 58488 20134 58500
rect 20346 58488 20352 58500
rect 20404 58528 20410 58540
rect 20625 58531 20683 58537
rect 20625 58528 20637 58531
rect 20404 58500 20637 58528
rect 20404 58488 20410 58500
rect 20625 58497 20637 58500
rect 20671 58497 20683 58531
rect 20625 58491 20683 58497
rect 23658 58488 23664 58540
rect 23716 58528 23722 58540
rect 24394 58528 24400 58540
rect 23716 58500 24400 58528
rect 23716 58488 23722 58500
rect 24394 58488 24400 58500
rect 24452 58528 24458 58540
rect 26053 58531 26111 58537
rect 26053 58528 26065 58531
rect 24452 58500 26065 58528
rect 24452 58488 24458 58500
rect 26053 58497 26065 58500
rect 26099 58497 26111 58531
rect 26053 58491 26111 58497
rect 26970 58488 26976 58540
rect 27028 58528 27034 58540
rect 27338 58528 27344 58540
rect 27028 58500 27344 58528
rect 27028 58488 27034 58500
rect 27338 58488 27344 58500
rect 27396 58488 27402 58540
rect 27724 58537 27752 58624
rect 27816 58543 27844 58636
rect 28626 58624 28632 58636
rect 28684 58624 28690 58676
rect 30006 58624 30012 58676
rect 30064 58664 30070 58676
rect 30101 58667 30159 58673
rect 30101 58664 30113 58667
rect 30064 58636 30113 58664
rect 30064 58624 30070 58636
rect 30101 58633 30113 58636
rect 30147 58633 30159 58667
rect 30101 58627 30159 58633
rect 29086 58556 29092 58608
rect 29144 58596 29150 58608
rect 30650 58596 30656 58608
rect 29144 58568 29592 58596
rect 29144 58556 29150 58568
rect 27801 58537 27859 58543
rect 27709 58531 27767 58537
rect 27709 58497 27721 58531
rect 27755 58497 27767 58531
rect 27801 58503 27813 58537
rect 27847 58503 27859 58537
rect 27801 58497 27859 58503
rect 27893 58531 27951 58537
rect 27893 58497 27905 58531
rect 27939 58528 27951 58531
rect 28077 58531 28135 58537
rect 27939 58500 28028 58528
rect 27939 58497 27951 58500
rect 27709 58491 27767 58497
rect 27893 58491 27951 58497
rect 21174 58460 21180 58472
rect 17368 58432 17413 58460
rect 18892 58432 21180 58460
rect 17368 58420 17374 58432
rect 21174 58420 21180 58432
rect 21232 58420 21238 58472
rect 1578 58392 1584 58404
rect 1539 58364 1584 58392
rect 1578 58352 1584 58364
rect 1636 58352 1642 58404
rect 16117 58395 16175 58401
rect 16117 58361 16129 58395
rect 16163 58392 16175 58395
rect 16482 58392 16488 58404
rect 16163 58364 16488 58392
rect 16163 58361 16175 58364
rect 16117 58355 16175 58361
rect 16482 58352 16488 58364
rect 16540 58352 16546 58404
rect 16758 58392 16764 58404
rect 16719 58364 16764 58392
rect 16758 58352 16764 58364
rect 16816 58352 16822 58404
rect 26326 58352 26332 58404
rect 26384 58392 26390 58404
rect 28000 58392 28028 58500
rect 28077 58497 28089 58531
rect 28123 58497 28135 58531
rect 28626 58528 28632 58540
rect 28587 58500 28632 58528
rect 28077 58491 28135 58497
rect 26384 58364 28028 58392
rect 26384 58352 26390 58364
rect 13538 58324 13544 58336
rect 13499 58296 13544 58324
rect 13538 58284 13544 58296
rect 13596 58284 13602 58336
rect 26970 58284 26976 58336
rect 27028 58324 27034 58336
rect 28092 58324 28120 58491
rect 28626 58488 28632 58500
rect 28684 58488 28690 58540
rect 29362 58528 29368 58540
rect 29323 58500 29368 58528
rect 29362 58488 29368 58500
rect 29420 58488 29426 58540
rect 29564 58537 29592 58568
rect 29656 58568 30656 58596
rect 29656 58537 29684 58568
rect 30650 58556 30656 58568
rect 30708 58596 30714 58608
rect 31202 58596 31208 58608
rect 30708 58568 31208 58596
rect 30708 58556 30714 58568
rect 31202 58556 31208 58568
rect 31260 58556 31266 58608
rect 29549 58531 29607 58537
rect 29549 58497 29561 58531
rect 29595 58497 29607 58531
rect 29549 58491 29607 58497
rect 29641 58531 29699 58537
rect 29641 58497 29653 58531
rect 29687 58497 29699 58531
rect 29641 58491 29699 58497
rect 29917 58531 29975 58537
rect 29917 58497 29929 58531
rect 29963 58528 29975 58531
rect 30006 58528 30012 58540
rect 29963 58500 30012 58528
rect 29963 58497 29975 58500
rect 29917 58491 29975 58497
rect 30006 58488 30012 58500
rect 30064 58488 30070 58540
rect 30374 58488 30380 58540
rect 30432 58488 30438 58540
rect 29733 58463 29791 58469
rect 28966 58432 29684 58460
rect 28813 58395 28871 58401
rect 28813 58361 28825 58395
rect 28859 58392 28871 58395
rect 28966 58392 28994 58432
rect 28859 58364 28994 58392
rect 29656 58392 29684 58432
rect 29733 58429 29745 58463
rect 29779 58460 29791 58463
rect 30392 58460 30420 58488
rect 31478 58460 31484 58472
rect 29779 58432 31484 58460
rect 29779 58429 29791 58432
rect 29733 58423 29791 58429
rect 31478 58420 31484 58432
rect 31536 58420 31542 58472
rect 30374 58392 30380 58404
rect 29656 58364 30380 58392
rect 28859 58361 28871 58364
rect 28813 58355 28871 58361
rect 30374 58352 30380 58364
rect 30432 58352 30438 58404
rect 27028 58296 28120 58324
rect 27028 58284 27034 58296
rect 29822 58284 29828 58336
rect 29880 58324 29886 58336
rect 30098 58324 30104 58336
rect 29880 58296 30104 58324
rect 29880 58284 29886 58296
rect 30098 58284 30104 58296
rect 30156 58284 30162 58336
rect 1104 58234 30820 58256
rect 1104 58182 5915 58234
rect 5967 58182 5979 58234
rect 6031 58182 6043 58234
rect 6095 58182 6107 58234
rect 6159 58182 6171 58234
rect 6223 58182 15846 58234
rect 15898 58182 15910 58234
rect 15962 58182 15974 58234
rect 16026 58182 16038 58234
rect 16090 58182 16102 58234
rect 16154 58182 25776 58234
rect 25828 58182 25840 58234
rect 25892 58182 25904 58234
rect 25956 58182 25968 58234
rect 26020 58182 26032 58234
rect 26084 58182 30820 58234
rect 1104 58160 30820 58182
rect 17221 58123 17279 58129
rect 17221 58089 17233 58123
rect 17267 58120 17279 58123
rect 18506 58120 18512 58132
rect 17267 58092 18512 58120
rect 17267 58089 17279 58092
rect 17221 58083 17279 58089
rect 18506 58080 18512 58092
rect 18564 58080 18570 58132
rect 25884 58092 28948 58120
rect 25884 58064 25912 58092
rect 13538 58012 13544 58064
rect 13596 58052 13602 58064
rect 21542 58052 21548 58064
rect 13596 58024 21548 58052
rect 13596 58012 13602 58024
rect 21542 58012 21548 58024
rect 21600 58012 21606 58064
rect 25866 58012 25872 58064
rect 25924 58012 25930 58064
rect 26513 58055 26571 58061
rect 26513 58021 26525 58055
rect 26559 58052 26571 58055
rect 27154 58052 27160 58064
rect 26559 58024 27160 58052
rect 26559 58021 26571 58024
rect 26513 58015 26571 58021
rect 27154 58012 27160 58024
rect 27212 58012 27218 58064
rect 15102 57944 15108 57996
rect 15160 57984 15166 57996
rect 17862 57984 17868 57996
rect 15160 57956 17868 57984
rect 15160 57944 15166 57956
rect 17862 57944 17868 57956
rect 17920 57944 17926 57996
rect 23014 57944 23020 57996
rect 23072 57984 23078 57996
rect 23658 57984 23664 57996
rect 23072 57956 23664 57984
rect 23072 57944 23078 57956
rect 23658 57944 23664 57956
rect 23716 57944 23722 57996
rect 28000 57956 28856 57984
rect 1397 57919 1455 57925
rect 1397 57885 1409 57919
rect 1443 57916 1455 57919
rect 2130 57916 2136 57928
rect 1443 57888 2136 57916
rect 1443 57885 1455 57888
rect 1397 57879 1455 57885
rect 2130 57876 2136 57888
rect 2188 57876 2194 57928
rect 13814 57876 13820 57928
rect 13872 57916 13878 57928
rect 15473 57919 15531 57925
rect 15473 57916 15485 57919
rect 13872 57888 15485 57916
rect 13872 57876 13878 57888
rect 15473 57885 15485 57888
rect 15519 57885 15531 57919
rect 15473 57879 15531 57885
rect 17218 57876 17224 57928
rect 17276 57916 17282 57928
rect 17497 57919 17555 57925
rect 17497 57916 17509 57919
rect 17276 57888 17509 57916
rect 17276 57876 17282 57888
rect 17497 57885 17509 57888
rect 17543 57885 17555 57919
rect 20717 57919 20775 57925
rect 20717 57916 20729 57919
rect 17497 57879 17555 57885
rect 17880 57888 20729 57916
rect 17880 57860 17908 57888
rect 20717 57885 20729 57888
rect 20763 57885 20775 57919
rect 20717 57879 20775 57885
rect 27065 57919 27123 57925
rect 27065 57885 27077 57919
rect 27111 57916 27123 57919
rect 27154 57916 27160 57928
rect 27111 57888 27160 57916
rect 27111 57885 27123 57888
rect 27065 57879 27123 57885
rect 27154 57876 27160 57888
rect 27212 57876 27218 57928
rect 15286 57848 15292 57860
rect 15247 57820 15292 57848
rect 15286 57808 15292 57820
rect 15344 57808 15350 57860
rect 16298 57848 16304 57860
rect 16259 57820 16304 57848
rect 16298 57808 16304 57820
rect 16356 57808 16362 57860
rect 16577 57851 16635 57857
rect 16577 57817 16589 57851
rect 16623 57848 16635 57851
rect 17310 57848 17316 57860
rect 16623 57820 17316 57848
rect 16623 57817 16635 57820
rect 16577 57811 16635 57817
rect 17310 57808 17316 57820
rect 17368 57848 17374 57860
rect 17773 57851 17831 57857
rect 17773 57848 17785 57851
rect 17368 57820 17785 57848
rect 17368 57808 17374 57820
rect 17773 57817 17785 57820
rect 17819 57817 17831 57851
rect 17773 57811 17831 57817
rect 17862 57808 17868 57860
rect 17920 57808 17926 57860
rect 18230 57808 18236 57860
rect 18288 57848 18294 57860
rect 18417 57851 18475 57857
rect 18417 57848 18429 57851
rect 18288 57820 18429 57848
rect 18288 57808 18294 57820
rect 18417 57817 18429 57820
rect 18463 57817 18475 57851
rect 18417 57811 18475 57817
rect 26329 57851 26387 57857
rect 26329 57817 26341 57851
rect 26375 57848 26387 57851
rect 26970 57848 26976 57860
rect 26375 57820 26976 57848
rect 26375 57817 26387 57820
rect 26329 57811 26387 57817
rect 26970 57808 26976 57820
rect 27028 57808 27034 57860
rect 27338 57808 27344 57860
rect 27396 57848 27402 57860
rect 27893 57851 27951 57857
rect 27893 57848 27905 57851
rect 27396 57820 27905 57848
rect 27396 57808 27402 57820
rect 27893 57817 27905 57820
rect 27939 57817 27951 57851
rect 27893 57811 27951 57817
rect 1578 57780 1584 57792
rect 1539 57752 1584 57780
rect 1578 57740 1584 57752
rect 1636 57740 1642 57792
rect 12986 57740 12992 57792
rect 13044 57780 13050 57792
rect 14182 57780 14188 57792
rect 13044 57752 14188 57780
rect 13044 57740 13050 57752
rect 14182 57740 14188 57752
rect 14240 57740 14246 57792
rect 15562 57740 15568 57792
rect 15620 57780 15626 57792
rect 16007 57783 16065 57789
rect 16007 57780 16019 57783
rect 15620 57752 16019 57780
rect 15620 57740 15626 57752
rect 16007 57749 16019 57752
rect 16053 57749 16065 57783
rect 16482 57780 16488 57792
rect 16443 57752 16488 57780
rect 16007 57743 16065 57749
rect 16482 57740 16488 57752
rect 16540 57740 16546 57792
rect 17586 57740 17592 57792
rect 17644 57780 17650 57792
rect 17681 57783 17739 57789
rect 17681 57780 17693 57783
rect 17644 57752 17693 57780
rect 17644 57740 17650 57752
rect 17681 57749 17693 57752
rect 17727 57780 17739 57783
rect 18509 57783 18567 57789
rect 18509 57780 18521 57783
rect 17727 57752 18521 57780
rect 17727 57749 17739 57752
rect 17681 57743 17739 57749
rect 18509 57749 18521 57752
rect 18555 57749 18567 57783
rect 18509 57743 18567 57749
rect 20438 57740 20444 57792
rect 20496 57780 20502 57792
rect 20901 57783 20959 57789
rect 20901 57780 20913 57783
rect 20496 57752 20913 57780
rect 20496 57740 20502 57752
rect 20901 57749 20913 57752
rect 20947 57749 20959 57783
rect 20901 57743 20959 57749
rect 26694 57740 26700 57792
rect 26752 57780 26758 57792
rect 27157 57783 27215 57789
rect 27157 57780 27169 57783
rect 26752 57752 27169 57780
rect 26752 57740 26758 57752
rect 27157 57749 27169 57752
rect 27203 57749 27215 57783
rect 27157 57743 27215 57749
rect 27430 57740 27436 57792
rect 27488 57780 27494 57792
rect 28000 57789 28028 57956
rect 28350 57876 28356 57928
rect 28408 57916 28414 57928
rect 28721 57919 28779 57925
rect 28721 57916 28733 57919
rect 28408 57888 28733 57916
rect 28408 57876 28414 57888
rect 27985 57783 28043 57789
rect 27985 57780 27997 57783
rect 27488 57752 27997 57780
rect 27488 57740 27494 57752
rect 27985 57749 27997 57752
rect 28031 57749 28043 57783
rect 27985 57743 28043 57749
rect 28166 57740 28172 57792
rect 28224 57780 28230 57792
rect 28537 57783 28595 57789
rect 28537 57780 28549 57783
rect 28224 57752 28549 57780
rect 28224 57740 28230 57752
rect 28537 57749 28549 57752
rect 28583 57749 28595 57783
rect 28644 57780 28672 57888
rect 28721 57885 28733 57888
rect 28767 57885 28779 57919
rect 28721 57879 28779 57885
rect 28828 57848 28856 57956
rect 28920 57925 28948 58092
rect 29362 58080 29368 58132
rect 29420 58120 29426 58132
rect 29549 58123 29607 58129
rect 29549 58120 29561 58123
rect 29420 58092 29561 58120
rect 29420 58080 29426 58092
rect 29549 58089 29561 58092
rect 29595 58089 29607 58123
rect 29549 58083 29607 58089
rect 28905 57919 28963 57925
rect 28905 57885 28917 57919
rect 28951 57885 28963 57919
rect 28905 57879 28963 57885
rect 28997 57919 29055 57925
rect 28997 57885 29009 57919
rect 29043 57885 29055 57919
rect 28997 57879 29055 57885
rect 29012 57848 29040 57879
rect 29086 57876 29092 57928
rect 29144 57916 29150 57928
rect 29362 57916 29368 57928
rect 29144 57888 29368 57916
rect 29144 57876 29150 57888
rect 29362 57876 29368 57888
rect 29420 57876 29426 57928
rect 29733 57919 29791 57925
rect 29733 57885 29745 57919
rect 29779 57885 29791 57919
rect 30009 57919 30067 57925
rect 30009 57916 30021 57919
rect 29733 57879 29791 57885
rect 29840 57888 30021 57916
rect 29748 57848 29776 57879
rect 28828 57820 29040 57848
rect 29104 57820 29776 57848
rect 29104 57792 29132 57820
rect 29086 57780 29092 57792
rect 28644 57752 29092 57780
rect 28537 57743 28595 57749
rect 29086 57740 29092 57752
rect 29144 57740 29150 57792
rect 29178 57740 29184 57792
rect 29236 57780 29242 57792
rect 29840 57780 29868 57888
rect 30009 57885 30021 57888
rect 30055 57885 30067 57919
rect 30009 57879 30067 57885
rect 29236 57752 29868 57780
rect 29917 57783 29975 57789
rect 29236 57740 29242 57752
rect 29917 57749 29929 57783
rect 29963 57780 29975 57783
rect 30098 57780 30104 57792
rect 29963 57752 30104 57780
rect 29963 57749 29975 57752
rect 29917 57743 29975 57749
rect 30098 57740 30104 57752
rect 30156 57740 30162 57792
rect 1104 57690 30820 57712
rect 1104 57638 10880 57690
rect 10932 57638 10944 57690
rect 10996 57638 11008 57690
rect 11060 57638 11072 57690
rect 11124 57638 11136 57690
rect 11188 57638 20811 57690
rect 20863 57638 20875 57690
rect 20927 57638 20939 57690
rect 20991 57638 21003 57690
rect 21055 57638 21067 57690
rect 21119 57638 30820 57690
rect 1104 57616 30820 57638
rect 1394 57536 1400 57588
rect 1452 57576 1458 57588
rect 2133 57579 2191 57585
rect 2133 57576 2145 57579
rect 1452 57548 2145 57576
rect 1452 57536 1458 57548
rect 2133 57545 2145 57548
rect 2179 57545 2191 57579
rect 2133 57539 2191 57545
rect 15286 57536 15292 57588
rect 15344 57576 15350 57588
rect 20530 57576 20536 57588
rect 15344 57548 20536 57576
rect 15344 57536 15350 57548
rect 20530 57536 20536 57548
rect 20588 57536 20594 57588
rect 25406 57536 25412 57588
rect 25464 57576 25470 57588
rect 25869 57579 25927 57585
rect 25869 57576 25881 57579
rect 25464 57548 25881 57576
rect 25464 57536 25470 57548
rect 25869 57545 25881 57548
rect 25915 57545 25927 57579
rect 25869 57539 25927 57545
rect 29730 57536 29736 57588
rect 29788 57576 29794 57588
rect 29825 57579 29883 57585
rect 29825 57576 29837 57579
rect 29788 57548 29837 57576
rect 29788 57536 29794 57548
rect 29825 57545 29837 57548
rect 29871 57545 29883 57579
rect 29825 57539 29883 57545
rect 14918 57517 14924 57520
rect 14912 57508 14924 57517
rect 14879 57480 14924 57508
rect 14912 57471 14924 57480
rect 14918 57468 14924 57471
rect 14976 57468 14982 57520
rect 20254 57468 20260 57520
rect 20312 57508 20318 57520
rect 20312 57480 21036 57508
rect 20312 57468 20318 57480
rect 1397 57443 1455 57449
rect 1397 57409 1409 57443
rect 1443 57440 1455 57443
rect 1854 57440 1860 57452
rect 1443 57412 1860 57440
rect 1443 57409 1455 57412
rect 1397 57403 1455 57409
rect 1854 57400 1860 57412
rect 1912 57400 1918 57452
rect 2317 57443 2375 57449
rect 2317 57409 2329 57443
rect 2363 57440 2375 57443
rect 2682 57440 2688 57452
rect 2363 57412 2688 57440
rect 2363 57409 2375 57412
rect 2317 57403 2375 57409
rect 2682 57400 2688 57412
rect 2740 57400 2746 57452
rect 13630 57400 13636 57452
rect 13688 57440 13694 57452
rect 13771 57443 13829 57449
rect 13771 57440 13783 57443
rect 13688 57412 13783 57440
rect 13688 57400 13694 57412
rect 13771 57409 13783 57412
rect 13817 57409 13829 57443
rect 13771 57403 13829 57409
rect 13906 57446 13964 57452
rect 13906 57412 13918 57446
rect 13952 57412 13964 57446
rect 13906 57406 13964 57412
rect 14001 57443 14059 57449
rect 14001 57409 14013 57443
rect 14047 57440 14059 57443
rect 14090 57440 14096 57452
rect 14047 57412 14096 57440
rect 14047 57409 14059 57412
rect 13924 57372 13952 57406
rect 14001 57403 14059 57409
rect 14090 57400 14096 57412
rect 14148 57400 14154 57452
rect 14182 57400 14188 57452
rect 14240 57440 14246 57452
rect 17037 57443 17095 57449
rect 14240 57412 14285 57440
rect 14240 57400 14246 57412
rect 17037 57409 17049 57443
rect 17083 57440 17095 57443
rect 17954 57440 17960 57452
rect 17083 57412 17960 57440
rect 17083 57409 17095 57412
rect 17037 57403 17095 57409
rect 17954 57400 17960 57412
rect 18012 57400 18018 57452
rect 19334 57400 19340 57452
rect 19392 57440 19398 57452
rect 19475 57443 19533 57449
rect 19475 57440 19487 57443
rect 19392 57412 19487 57440
rect 19392 57400 19398 57412
rect 19475 57409 19487 57412
rect 19521 57409 19533 57443
rect 19610 57440 19616 57452
rect 19571 57412 19616 57440
rect 19475 57403 19533 57409
rect 19610 57400 19616 57412
rect 19668 57400 19674 57452
rect 19705 57443 19763 57449
rect 19705 57409 19717 57443
rect 19751 57440 19763 57443
rect 19794 57440 19800 57452
rect 19751 57412 19800 57440
rect 19751 57409 19763 57412
rect 19705 57403 19763 57409
rect 19794 57400 19800 57412
rect 19852 57400 19858 57452
rect 19886 57400 19892 57452
rect 19944 57440 19950 57452
rect 20622 57440 20628 57452
rect 19944 57412 19989 57440
rect 20583 57412 20628 57440
rect 19944 57400 19950 57412
rect 20622 57400 20628 57412
rect 20680 57400 20686 57452
rect 20717 57443 20775 57449
rect 20717 57409 20729 57443
rect 20763 57409 20775 57443
rect 20717 57403 20775 57409
rect 14645 57375 14703 57381
rect 13924 57344 13965 57372
rect 13814 57264 13820 57316
rect 13872 57304 13878 57316
rect 13937 57304 13965 57344
rect 14645 57341 14657 57375
rect 14691 57341 14703 57375
rect 19628 57372 19656 57400
rect 20732 57372 20760 57403
rect 20806 57400 20812 57452
rect 20864 57440 20870 57452
rect 21008 57449 21036 57480
rect 21082 57468 21088 57520
rect 21140 57508 21146 57520
rect 26237 57511 26295 57517
rect 21140 57480 22094 57508
rect 21140 57468 21146 57480
rect 20993 57443 21051 57449
rect 20864 57412 20909 57440
rect 20864 57400 20870 57412
rect 20993 57409 21005 57443
rect 21039 57409 21051 57443
rect 22066 57440 22094 57480
rect 26237 57477 26249 57511
rect 26283 57508 26295 57511
rect 26602 57508 26608 57520
rect 26283 57480 26608 57508
rect 26283 57477 26295 57480
rect 26237 57471 26295 57477
rect 26602 57468 26608 57480
rect 26660 57468 26666 57520
rect 26712 57480 29316 57508
rect 22833 57443 22891 57449
rect 22833 57440 22845 57443
rect 22066 57412 22845 57440
rect 20993 57403 21051 57409
rect 22833 57409 22845 57412
rect 22879 57409 22891 57443
rect 22833 57403 22891 57409
rect 23017 57443 23075 57449
rect 23017 57409 23029 57443
rect 23063 57440 23075 57443
rect 23106 57440 23112 57452
rect 23063 57412 23112 57440
rect 23063 57409 23075 57412
rect 23017 57403 23075 57409
rect 23106 57400 23112 57412
rect 23164 57400 23170 57452
rect 23934 57440 23940 57452
rect 23895 57412 23940 57440
rect 23934 57400 23940 57412
rect 23992 57400 23998 57452
rect 26050 57440 26056 57452
rect 26011 57412 26056 57440
rect 26050 57400 26056 57412
rect 26108 57400 26114 57452
rect 26326 57440 26332 57452
rect 26287 57412 26332 57440
rect 26326 57400 26332 57412
rect 26384 57400 26390 57452
rect 19628 57344 20760 57372
rect 14645 57335 14703 57341
rect 13872 57276 13965 57304
rect 13872 57264 13878 57276
rect 1578 57236 1584 57248
rect 1539 57208 1584 57236
rect 1578 57196 1584 57208
rect 1636 57196 1642 57248
rect 13541 57239 13599 57245
rect 13541 57205 13553 57239
rect 13587 57236 13599 57239
rect 14182 57236 14188 57248
rect 13587 57208 14188 57236
rect 13587 57205 13599 57208
rect 13541 57199 13599 57205
rect 14182 57196 14188 57208
rect 14240 57196 14246 57248
rect 14660 57236 14688 57335
rect 21726 57332 21732 57384
rect 21784 57372 21790 57384
rect 25866 57372 25872 57384
rect 21784 57344 25872 57372
rect 21784 57332 21790 57344
rect 25866 57332 25872 57344
rect 25924 57332 25930 57384
rect 20714 57264 20720 57316
rect 20772 57304 20778 57316
rect 21266 57304 21272 57316
rect 20772 57276 21272 57304
rect 20772 57264 20778 57276
rect 21266 57264 21272 57276
rect 21324 57264 21330 57316
rect 23201 57307 23259 57313
rect 23201 57273 23213 57307
rect 23247 57304 23259 57307
rect 26712 57304 26740 57480
rect 26970 57440 26976 57452
rect 26931 57412 26976 57440
rect 26970 57400 26976 57412
rect 27028 57400 27034 57452
rect 27338 57332 27344 57384
rect 27396 57372 27402 57384
rect 28353 57375 28411 57381
rect 28353 57372 28365 57375
rect 27396 57344 28365 57372
rect 27396 57332 27402 57344
rect 28353 57341 28365 57344
rect 28399 57341 28411 57375
rect 28353 57335 28411 57341
rect 28629 57375 28687 57381
rect 28629 57341 28641 57375
rect 28675 57372 28687 57375
rect 29178 57372 29184 57384
rect 28675 57344 29184 57372
rect 28675 57341 28687 57344
rect 28629 57335 28687 57341
rect 29178 57332 29184 57344
rect 29236 57332 29242 57384
rect 29288 57372 29316 57480
rect 29730 57440 29736 57452
rect 29691 57412 29736 57440
rect 29730 57400 29736 57412
rect 29788 57400 29794 57452
rect 29288 57344 29776 57372
rect 29748 57316 29776 57344
rect 23247 57276 26740 57304
rect 23247 57273 23259 57276
rect 23201 57267 23259 57273
rect 29730 57264 29736 57316
rect 29788 57264 29794 57316
rect 15378 57236 15384 57248
rect 14660 57208 15384 57236
rect 15378 57196 15384 57208
rect 15436 57196 15442 57248
rect 15654 57196 15660 57248
rect 15712 57236 15718 57248
rect 16025 57239 16083 57245
rect 16025 57236 16037 57239
rect 15712 57208 16037 57236
rect 15712 57196 15718 57208
rect 16025 57205 16037 57208
rect 16071 57205 16083 57239
rect 18322 57236 18328 57248
rect 18283 57208 18328 57236
rect 16025 57199 16083 57205
rect 18322 57196 18328 57208
rect 18380 57196 18386 57248
rect 18414 57196 18420 57248
rect 18472 57236 18478 57248
rect 19245 57239 19303 57245
rect 19245 57236 19257 57239
rect 18472 57208 19257 57236
rect 18472 57196 18478 57208
rect 19245 57205 19257 57208
rect 19291 57205 19303 57239
rect 20346 57236 20352 57248
rect 20307 57208 20352 57236
rect 19245 57199 19303 57205
rect 20346 57196 20352 57208
rect 20404 57196 20410 57248
rect 21542 57196 21548 57248
rect 21600 57236 21606 57248
rect 23014 57236 23020 57248
rect 21600 57208 23020 57236
rect 21600 57196 21606 57208
rect 23014 57196 23020 57208
rect 23072 57196 23078 57248
rect 23753 57239 23811 57245
rect 23753 57205 23765 57239
rect 23799 57236 23811 57239
rect 24118 57236 24124 57248
rect 23799 57208 24124 57236
rect 23799 57205 23811 57208
rect 23753 57199 23811 57205
rect 24118 57196 24124 57208
rect 24176 57196 24182 57248
rect 24394 57196 24400 57248
rect 24452 57236 24458 57248
rect 27157 57239 27215 57245
rect 27157 57236 27169 57239
rect 24452 57208 27169 57236
rect 24452 57196 24458 57208
rect 27157 57205 27169 57208
rect 27203 57205 27215 57239
rect 27157 57199 27215 57205
rect 28166 57196 28172 57248
rect 28224 57236 28230 57248
rect 30650 57236 30656 57248
rect 28224 57208 30656 57236
rect 28224 57196 28230 57208
rect 30650 57196 30656 57208
rect 30708 57196 30714 57248
rect 1104 57146 30820 57168
rect 1104 57094 5915 57146
rect 5967 57094 5979 57146
rect 6031 57094 6043 57146
rect 6095 57094 6107 57146
rect 6159 57094 6171 57146
rect 6223 57094 15846 57146
rect 15898 57094 15910 57146
rect 15962 57094 15974 57146
rect 16026 57094 16038 57146
rect 16090 57094 16102 57146
rect 16154 57094 25776 57146
rect 25828 57094 25840 57146
rect 25892 57094 25904 57146
rect 25956 57094 25968 57146
rect 26020 57094 26032 57146
rect 26084 57094 30820 57146
rect 1104 57072 30820 57094
rect 2130 57032 2136 57044
rect 2091 57004 2136 57032
rect 2130 56992 2136 57004
rect 2188 56992 2194 57044
rect 13630 56992 13636 57044
rect 13688 57032 13694 57044
rect 16206 57032 16212 57044
rect 13688 57004 15516 57032
rect 16167 57004 16212 57032
rect 13688 56992 13694 57004
rect 15488 56973 15516 57004
rect 16206 56992 16212 57004
rect 16264 56992 16270 57044
rect 16761 57035 16819 57041
rect 16761 57001 16773 57035
rect 16807 57032 16819 57035
rect 17678 57032 17684 57044
rect 16807 57004 17684 57032
rect 16807 57001 16819 57004
rect 16761 56995 16819 57001
rect 17678 56992 17684 57004
rect 17736 56992 17742 57044
rect 21082 57032 21088 57044
rect 17788 57004 21088 57032
rect 13541 56967 13599 56973
rect 13541 56933 13553 56967
rect 13587 56964 13599 56967
rect 15473 56967 15531 56973
rect 13587 56936 14136 56964
rect 13587 56933 13599 56936
rect 13541 56927 13599 56933
rect 14108 56905 14136 56936
rect 15473 56933 15485 56967
rect 15519 56964 15531 56967
rect 17788 56964 17816 57004
rect 21082 56992 21088 57004
rect 21140 56992 21146 57044
rect 21542 56992 21548 57044
rect 21600 57032 21606 57044
rect 21600 57004 22784 57032
rect 21600 56992 21606 57004
rect 15519 56936 17816 56964
rect 15519 56933 15531 56936
rect 15473 56927 15531 56933
rect 21358 56924 21364 56976
rect 21416 56964 21422 56976
rect 22554 56964 22560 56976
rect 21416 56936 22560 56964
rect 21416 56924 21422 56936
rect 22554 56924 22560 56936
rect 22612 56924 22618 56976
rect 14093 56899 14151 56905
rect 14093 56865 14105 56899
rect 14139 56865 14151 56899
rect 17218 56896 17224 56908
rect 17179 56868 17224 56896
rect 14093 56859 14151 56865
rect 17218 56856 17224 56868
rect 17276 56856 17282 56908
rect 17494 56856 17500 56908
rect 17552 56896 17558 56908
rect 17862 56896 17868 56908
rect 17552 56868 17868 56896
rect 17552 56856 17558 56868
rect 17862 56856 17868 56868
rect 17920 56856 17926 56908
rect 21376 56896 21404 56924
rect 21376 56868 21496 56896
rect 1394 56828 1400 56840
rect 1355 56800 1400 56828
rect 1394 56788 1400 56800
rect 1452 56788 1458 56840
rect 2317 56831 2375 56837
rect 2317 56797 2329 56831
rect 2363 56828 2375 56831
rect 2590 56828 2596 56840
rect 2363 56800 2596 56828
rect 2363 56797 2375 56800
rect 2317 56791 2375 56797
rect 2590 56788 2596 56800
rect 2648 56788 2654 56840
rect 13357 56831 13415 56837
rect 13357 56797 13369 56831
rect 13403 56828 13415 56831
rect 13998 56828 14004 56840
rect 13403 56800 14004 56828
rect 13403 56797 13415 56800
rect 13357 56791 13415 56797
rect 13998 56788 14004 56800
rect 14056 56788 14062 56840
rect 14182 56788 14188 56840
rect 14240 56828 14246 56840
rect 14349 56831 14407 56837
rect 14349 56828 14361 56831
rect 14240 56800 14361 56828
rect 14240 56788 14246 56800
rect 14349 56797 14361 56800
rect 14395 56797 14407 56831
rect 14349 56791 14407 56797
rect 16025 56831 16083 56837
rect 16025 56797 16037 56831
rect 16071 56828 16083 56831
rect 17678 56828 17684 56840
rect 16071 56800 17684 56828
rect 16071 56797 16083 56800
rect 16025 56791 16083 56797
rect 17678 56788 17684 56800
rect 17736 56788 17742 56840
rect 18141 56831 18199 56837
rect 18141 56797 18153 56831
rect 18187 56797 18199 56831
rect 19242 56828 19248 56840
rect 19203 56800 19248 56828
rect 18141 56791 18199 56797
rect 17310 56760 17316 56772
rect 17271 56732 17316 56760
rect 17310 56720 17316 56732
rect 17368 56720 17374 56772
rect 18156 56760 18184 56791
rect 19242 56788 19248 56800
rect 19300 56788 19306 56840
rect 19512 56831 19570 56837
rect 19512 56797 19524 56831
rect 19558 56828 19570 56831
rect 20346 56828 20352 56840
rect 19558 56800 20352 56828
rect 19558 56797 19570 56800
rect 19512 56791 19570 56797
rect 20346 56788 20352 56800
rect 20404 56788 20410 56840
rect 21266 56788 21272 56840
rect 21324 56837 21330 56840
rect 21468 56837 21496 56868
rect 21324 56831 21373 56837
rect 21324 56797 21327 56831
rect 21361 56797 21373 56831
rect 21324 56791 21373 56797
rect 21453 56831 21511 56837
rect 21453 56797 21465 56831
rect 21499 56797 21511 56831
rect 21453 56791 21511 56797
rect 21324 56788 21330 56791
rect 21542 56788 21548 56840
rect 21600 56828 21606 56840
rect 21729 56831 21787 56837
rect 21600 56800 21693 56828
rect 21600 56788 21606 56800
rect 21729 56797 21741 56831
rect 21775 56828 21787 56831
rect 21818 56828 21824 56840
rect 21775 56800 21824 56828
rect 21775 56797 21787 56800
rect 21729 56791 21787 56797
rect 21818 56788 21824 56800
rect 21876 56788 21882 56840
rect 22569 56837 22597 56924
rect 22465 56831 22523 56837
rect 22296 56825 22416 56828
rect 22465 56825 22477 56831
rect 22296 56800 22477 56825
rect 19794 56760 19800 56772
rect 18156 56732 19800 56760
rect 19794 56720 19800 56732
rect 19852 56720 19858 56772
rect 20254 56720 20260 56772
rect 20312 56760 20318 56772
rect 20438 56760 20444 56772
rect 20312 56732 20444 56760
rect 20312 56720 20318 56732
rect 20438 56720 20444 56732
rect 20496 56760 20502 56772
rect 21560 56760 21588 56788
rect 20496 56732 21588 56760
rect 20496 56720 20502 56732
rect 1578 56692 1584 56704
rect 1539 56664 1584 56692
rect 1578 56652 1584 56664
rect 1636 56652 1642 56704
rect 17221 56695 17279 56701
rect 17221 56661 17233 56695
rect 17267 56692 17279 56695
rect 17586 56692 17592 56704
rect 17267 56664 17592 56692
rect 17267 56661 17279 56664
rect 17221 56655 17279 56661
rect 17586 56652 17592 56664
rect 17644 56652 17650 56704
rect 20622 56692 20628 56704
rect 20583 56664 20628 56692
rect 20622 56652 20628 56664
rect 20680 56652 20686 56704
rect 21085 56695 21143 56701
rect 21085 56661 21097 56695
rect 21131 56692 21143 56695
rect 21818 56692 21824 56704
rect 21131 56664 21824 56692
rect 21131 56661 21143 56664
rect 21085 56655 21143 56661
rect 21818 56652 21824 56664
rect 21876 56652 21882 56704
rect 22094 56652 22100 56704
rect 22152 56692 22158 56704
rect 22189 56695 22247 56701
rect 22189 56692 22201 56695
rect 22152 56664 22201 56692
rect 22152 56652 22158 56664
rect 22189 56661 22201 56664
rect 22235 56661 22247 56695
rect 22296 56692 22324 56800
rect 22388 56797 22477 56800
rect 22511 56797 22523 56831
rect 22465 56791 22523 56797
rect 22554 56831 22612 56837
rect 22554 56797 22566 56831
rect 22600 56797 22612 56831
rect 22554 56791 22612 56797
rect 22649 56831 22707 56837
rect 22649 56797 22661 56831
rect 22695 56806 22707 56831
rect 22756 56806 22784 57004
rect 23658 56992 23664 57044
rect 23716 57032 23722 57044
rect 23716 57004 25544 57032
rect 23716 56992 23722 57004
rect 23474 56924 23480 56976
rect 23532 56964 23538 56976
rect 24486 56964 24492 56976
rect 23532 56936 24492 56964
rect 23532 56924 23538 56936
rect 24486 56924 24492 56936
rect 24544 56924 24550 56976
rect 25516 56964 25544 57004
rect 25590 56992 25596 57044
rect 25648 57032 25654 57044
rect 25685 57035 25743 57041
rect 25685 57032 25697 57035
rect 25648 57004 25697 57032
rect 25648 56992 25654 57004
rect 25685 57001 25697 57004
rect 25731 57001 25743 57035
rect 26326 57032 26332 57044
rect 25685 56995 25743 57001
rect 26252 57004 26332 57032
rect 25516 56936 26004 56964
rect 24946 56856 24952 56908
rect 25004 56896 25010 56908
rect 25590 56896 25596 56908
rect 25004 56868 25596 56896
rect 25004 56856 25010 56868
rect 25590 56856 25596 56868
rect 25648 56856 25654 56908
rect 25976 56896 26004 56936
rect 25976 56868 26096 56896
rect 22695 56797 22784 56806
rect 22649 56791 22784 56797
rect 22845 56831 22903 56837
rect 22845 56797 22857 56831
rect 22891 56828 22903 56831
rect 23014 56828 23020 56840
rect 22891 56800 23020 56828
rect 22891 56797 22903 56800
rect 22845 56791 22903 56797
rect 22664 56778 22784 56791
rect 23014 56788 23020 56800
rect 23072 56788 23078 56840
rect 24118 56788 24124 56840
rect 24176 56828 24182 56840
rect 24578 56828 24584 56840
rect 24176 56800 24584 56828
rect 24176 56788 24182 56800
rect 24578 56788 24584 56800
rect 24636 56788 24642 56840
rect 25222 56788 25228 56840
rect 25280 56828 25286 56840
rect 25869 56831 25927 56837
rect 25869 56828 25881 56831
rect 25280 56800 25881 56828
rect 25280 56788 25286 56800
rect 25869 56797 25881 56800
rect 25915 56828 25927 56831
rect 25958 56828 25964 56840
rect 25915 56800 25964 56828
rect 25915 56797 25927 56800
rect 25869 56791 25927 56797
rect 25958 56788 25964 56800
rect 26016 56788 26022 56840
rect 26068 56837 26096 56868
rect 26252 56840 26280 57004
rect 26326 56992 26332 57004
rect 26384 56992 26390 57044
rect 27709 57035 27767 57041
rect 27709 57001 27721 57035
rect 27755 57032 27767 57035
rect 28399 57035 28457 57041
rect 27755 57004 28304 57032
rect 27755 57001 27767 57004
rect 27709 56995 27767 57001
rect 27338 56964 27344 56976
rect 27264 56936 27344 56964
rect 27264 56896 27292 56936
rect 27338 56924 27344 56936
rect 27396 56924 27402 56976
rect 27920 56936 28028 56964
rect 27080 56868 27292 56896
rect 26053 56831 26111 56837
rect 26053 56797 26065 56831
rect 26099 56797 26111 56831
rect 26053 56791 26111 56797
rect 26145 56831 26203 56837
rect 26145 56797 26157 56831
rect 26191 56828 26203 56831
rect 26234 56828 26240 56840
rect 26191 56800 26240 56828
rect 26191 56797 26203 56800
rect 26145 56791 26203 56797
rect 26234 56788 26240 56800
rect 26292 56788 26298 56840
rect 26973 56831 27031 56837
rect 26973 56797 26985 56831
rect 27019 56797 27031 56831
rect 26973 56791 27031 56797
rect 23382 56760 23388 56772
rect 23343 56732 23388 56760
rect 23382 56720 23388 56732
rect 23440 56720 23446 56772
rect 24394 56760 24400 56772
rect 24355 56732 24400 56760
rect 24394 56720 24400 56732
rect 24452 56720 24458 56772
rect 24946 56760 24952 56772
rect 24907 56732 24952 56760
rect 24946 56720 24952 56732
rect 25004 56720 25010 56772
rect 26988 56760 27016 56791
rect 25884 56732 27016 56760
rect 25884 56704 25912 56732
rect 22462 56692 22468 56704
rect 22296 56664 22468 56692
rect 22189 56655 22247 56661
rect 22462 56652 22468 56664
rect 22520 56652 22526 56704
rect 22738 56652 22744 56704
rect 22796 56692 22802 56704
rect 23477 56695 23535 56701
rect 23477 56692 23489 56695
rect 22796 56664 23489 56692
rect 22796 56652 22802 56664
rect 23477 56661 23489 56664
rect 23523 56661 23535 56695
rect 23477 56655 23535 56661
rect 24486 56652 24492 56704
rect 24544 56692 24550 56704
rect 24673 56695 24731 56701
rect 24673 56692 24685 56695
rect 24544 56664 24685 56692
rect 24544 56652 24550 56664
rect 24673 56661 24685 56664
rect 24719 56661 24731 56695
rect 24673 56655 24731 56661
rect 24765 56695 24823 56701
rect 24765 56661 24777 56695
rect 24811 56692 24823 56695
rect 25222 56692 25228 56704
rect 24811 56664 25228 56692
rect 24811 56661 24823 56664
rect 24765 56655 24823 56661
rect 25222 56652 25228 56664
rect 25280 56652 25286 56704
rect 25866 56652 25872 56704
rect 25924 56652 25930 56704
rect 26050 56652 26056 56704
rect 26108 56692 26114 56704
rect 27080 56692 27108 56868
rect 27264 56837 27292 56868
rect 27430 56856 27436 56908
rect 27488 56896 27494 56908
rect 27920 56896 27948 56936
rect 27488 56868 27948 56896
rect 28000 56896 28028 56936
rect 28169 56899 28227 56905
rect 28169 56896 28181 56899
rect 28000 56868 28181 56896
rect 27488 56856 27494 56868
rect 28169 56865 28181 56868
rect 28215 56865 28227 56899
rect 28276 56896 28304 57004
rect 28399 57001 28411 57035
rect 28445 57032 28457 57035
rect 29086 57032 29092 57044
rect 28445 57004 29092 57032
rect 28445 57001 28457 57004
rect 28399 56995 28457 57001
rect 29086 56992 29092 57004
rect 29144 56992 29150 57044
rect 29733 57035 29791 57041
rect 29733 57001 29745 57035
rect 29779 57032 29791 57035
rect 30558 57032 30564 57044
rect 29779 57004 30564 57032
rect 29779 57001 29791 57004
rect 29733 56995 29791 57001
rect 28276 56868 28574 56896
rect 28169 56859 28227 56865
rect 27157 56831 27215 56837
rect 27157 56797 27169 56831
rect 27203 56797 27215 56831
rect 27157 56791 27215 56797
rect 27249 56831 27307 56837
rect 27249 56797 27261 56831
rect 27295 56797 27307 56831
rect 27249 56791 27307 56797
rect 27172 56760 27200 56791
rect 27338 56788 27344 56840
rect 27396 56828 27402 56840
rect 27525 56831 27583 56837
rect 27396 56800 27441 56828
rect 27396 56788 27402 56800
rect 27525 56797 27537 56831
rect 27571 56828 27583 56831
rect 28546 56830 28574 56868
rect 29086 56856 29092 56908
rect 29144 56896 29150 56908
rect 30116 56896 30144 57004
rect 30558 56992 30564 57004
rect 30616 56992 30622 57044
rect 29144 56868 30144 56896
rect 29144 56856 29150 56868
rect 28718 56830 28724 56840
rect 27571 56822 27844 56828
rect 28546 56826 28580 56830
rect 28644 56826 28724 56830
rect 27571 56800 28233 56822
rect 28546 56802 28724 56826
rect 27571 56797 27583 56800
rect 27525 56791 27583 56797
rect 27816 56794 28233 56800
rect 28552 56798 28672 56802
rect 28205 56760 28233 56794
rect 28718 56788 28724 56802
rect 28776 56788 28782 56840
rect 29730 56828 29736 56840
rect 29691 56800 29736 56828
rect 29730 56788 29736 56800
rect 29788 56788 29794 56840
rect 30006 56760 30012 56772
rect 27172 56732 28101 56760
rect 28205 56732 30012 56760
rect 26108 56664 27108 56692
rect 28073 56692 28101 56732
rect 30006 56720 30012 56732
rect 30064 56720 30070 56772
rect 28166 56692 28172 56704
rect 28073 56664 28172 56692
rect 26108 56652 26114 56664
rect 28166 56652 28172 56664
rect 28224 56652 28230 56704
rect 1104 56602 30820 56624
rect 1104 56550 10880 56602
rect 10932 56550 10944 56602
rect 10996 56550 11008 56602
rect 11060 56550 11072 56602
rect 11124 56550 11136 56602
rect 11188 56550 20811 56602
rect 20863 56550 20875 56602
rect 20927 56550 20939 56602
rect 20991 56550 21003 56602
rect 21055 56550 21067 56602
rect 21119 56550 30820 56602
rect 1104 56528 30820 56550
rect 1854 56448 1860 56500
rect 1912 56488 1918 56500
rect 2133 56491 2191 56497
rect 2133 56488 2145 56491
rect 1912 56460 2145 56488
rect 1912 56448 1918 56460
rect 2133 56457 2145 56460
rect 2179 56457 2191 56491
rect 15378 56488 15384 56500
rect 15339 56460 15384 56488
rect 2133 56451 2191 56457
rect 15378 56448 15384 56460
rect 15436 56448 15442 56500
rect 22462 56448 22468 56500
rect 22520 56488 22526 56500
rect 23014 56488 23020 56500
rect 22520 56460 23020 56488
rect 22520 56448 22526 56460
rect 23014 56448 23020 56460
rect 23072 56488 23078 56500
rect 23201 56491 23259 56497
rect 23201 56488 23213 56491
rect 23072 56460 23213 56488
rect 23072 56448 23078 56460
rect 23201 56457 23213 56460
rect 23247 56457 23259 56491
rect 23201 56451 23259 56457
rect 23566 56448 23572 56500
rect 23624 56488 23630 56500
rect 24394 56488 24400 56500
rect 23624 56460 24400 56488
rect 23624 56448 23630 56460
rect 24394 56448 24400 56460
rect 24452 56448 24458 56500
rect 24489 56491 24547 56497
rect 24489 56457 24501 56491
rect 24535 56457 24547 56491
rect 24489 56451 24547 56457
rect 14461 56423 14519 56429
rect 14461 56389 14473 56423
rect 14507 56420 14519 56423
rect 16482 56420 16488 56432
rect 14507 56392 16488 56420
rect 14507 56389 14519 56392
rect 14461 56383 14519 56389
rect 16482 56380 16488 56392
rect 16540 56380 16546 56432
rect 17304 56423 17362 56429
rect 17304 56389 17316 56423
rect 17350 56420 17362 56423
rect 18414 56420 18420 56432
rect 17350 56392 18420 56420
rect 17350 56389 17362 56392
rect 17304 56383 17362 56389
rect 18414 56380 18420 56392
rect 18472 56380 18478 56432
rect 22738 56420 22744 56432
rect 21836 56392 22744 56420
rect 1397 56355 1455 56361
rect 1397 56321 1409 56355
rect 1443 56352 1455 56355
rect 2130 56352 2136 56364
rect 1443 56324 2136 56352
rect 1443 56321 1455 56324
rect 1397 56315 1455 56321
rect 2130 56312 2136 56324
rect 2188 56312 2194 56364
rect 2314 56352 2320 56364
rect 2275 56324 2320 56352
rect 2314 56312 2320 56324
rect 2372 56312 2378 56364
rect 14553 56355 14611 56361
rect 14553 56321 14565 56355
rect 14599 56352 14611 56355
rect 14734 56352 14740 56364
rect 14599 56324 14740 56352
rect 14599 56321 14611 56324
rect 14553 56315 14611 56321
rect 14734 56312 14740 56324
rect 14792 56312 14798 56364
rect 15197 56355 15255 56361
rect 15197 56321 15209 56355
rect 15243 56352 15255 56355
rect 15562 56352 15568 56364
rect 15243 56324 15568 56352
rect 15243 56321 15255 56324
rect 15197 56315 15255 56321
rect 15562 56312 15568 56324
rect 15620 56312 15626 56364
rect 15933 56355 15991 56361
rect 15933 56321 15945 56355
rect 15979 56352 15991 56355
rect 17586 56352 17592 56364
rect 15979 56324 17592 56352
rect 15979 56321 15991 56324
rect 15933 56315 15991 56321
rect 17586 56312 17592 56324
rect 17644 56312 17650 56364
rect 18877 56355 18935 56361
rect 18877 56321 18889 56355
rect 18923 56352 18935 56355
rect 19058 56352 19064 56364
rect 18923 56324 19064 56352
rect 18923 56321 18935 56324
rect 18877 56315 18935 56321
rect 19058 56312 19064 56324
rect 19116 56312 19122 56364
rect 21836 56361 21864 56392
rect 22738 56380 22744 56392
rect 22796 56380 22802 56432
rect 24210 56380 24216 56432
rect 24268 56420 24274 56432
rect 24504 56420 24532 56451
rect 25038 56448 25044 56500
rect 25096 56488 25102 56500
rect 25406 56488 25412 56500
rect 25096 56460 25412 56488
rect 25096 56448 25102 56460
rect 25406 56448 25412 56460
rect 25464 56448 25470 56500
rect 25682 56448 25688 56500
rect 25740 56488 25746 56500
rect 25777 56491 25835 56497
rect 25777 56488 25789 56491
rect 25740 56460 25789 56488
rect 25740 56448 25746 56460
rect 25777 56457 25789 56460
rect 25823 56457 25835 56491
rect 25777 56451 25835 56457
rect 25866 56448 25872 56500
rect 25924 56488 25930 56500
rect 28353 56491 28411 56497
rect 28353 56488 28365 56491
rect 25924 56460 28365 56488
rect 25924 56448 25930 56460
rect 28353 56457 28365 56460
rect 28399 56457 28411 56491
rect 29178 56488 29184 56500
rect 28353 56451 28411 56457
rect 28828 56460 29184 56488
rect 24268 56392 24532 56420
rect 25976 56392 27292 56420
rect 24268 56380 24274 56392
rect 25976 56364 26004 56392
rect 22094 56361 22100 56364
rect 21821 56355 21879 56361
rect 21821 56321 21833 56355
rect 21867 56321 21879 56355
rect 21821 56315 21879 56321
rect 22088 56315 22100 56361
rect 22152 56352 22158 56364
rect 22152 56324 22188 56352
rect 22094 56312 22100 56315
rect 22152 56312 22158 56324
rect 23290 56312 23296 56364
rect 23348 56352 23354 56364
rect 24118 56352 24124 56364
rect 23348 56324 24124 56352
rect 23348 56312 23354 56324
rect 24118 56312 24124 56324
rect 24176 56352 24182 56364
rect 24305 56355 24363 56361
rect 24305 56352 24317 56355
rect 24176 56324 24317 56352
rect 24176 56312 24182 56324
rect 24305 56321 24317 56324
rect 24351 56321 24363 56355
rect 24305 56315 24363 56321
rect 24394 56312 24400 56364
rect 24452 56352 24458 56364
rect 24673 56355 24731 56361
rect 24673 56352 24685 56355
rect 24452 56324 24685 56352
rect 24452 56312 24458 56324
rect 24673 56321 24685 56324
rect 24719 56321 24731 56355
rect 25958 56352 25964 56364
rect 25919 56324 25964 56352
rect 24673 56315 24731 56321
rect 25958 56312 25964 56324
rect 26016 56312 26022 56364
rect 26145 56355 26203 56361
rect 26145 56321 26157 56355
rect 26191 56321 26203 56355
rect 26145 56315 26203 56321
rect 14458 56284 14464 56296
rect 14419 56256 14464 56284
rect 14458 56244 14464 56256
rect 14516 56244 14522 56296
rect 17037 56287 17095 56293
rect 17037 56253 17049 56287
rect 17083 56253 17095 56287
rect 26160 56284 26188 56315
rect 26234 56312 26240 56364
rect 26292 56352 26298 56364
rect 27264 56361 27292 56392
rect 27249 56355 27307 56361
rect 26292 56324 26337 56352
rect 26292 56312 26298 56324
rect 27249 56321 27261 56355
rect 27295 56321 27307 56355
rect 27249 56315 27307 56321
rect 28537 56355 28595 56361
rect 28537 56321 28549 56355
rect 28583 56321 28595 56355
rect 28718 56352 28724 56364
rect 28679 56324 28724 56352
rect 28537 56315 28595 56321
rect 17037 56247 17095 56253
rect 23124 56256 26188 56284
rect 26973 56287 27031 56293
rect 13998 56216 14004 56228
rect 13959 56188 14004 56216
rect 13998 56176 14004 56188
rect 14056 56176 14062 56228
rect 1578 56148 1584 56160
rect 1539 56120 1584 56148
rect 1578 56108 1584 56120
rect 1636 56108 1642 56160
rect 14090 56108 14096 56160
rect 14148 56148 14154 56160
rect 16025 56151 16083 56157
rect 16025 56148 16037 56151
rect 14148 56120 16037 56148
rect 14148 56108 14154 56120
rect 16025 56117 16037 56120
rect 16071 56117 16083 56151
rect 17052 56148 17080 56247
rect 18046 56148 18052 56160
rect 17052 56120 18052 56148
rect 16025 56111 16083 56117
rect 18046 56108 18052 56120
rect 18104 56108 18110 56160
rect 18417 56151 18475 56157
rect 18417 56117 18429 56151
rect 18463 56148 18475 56151
rect 19334 56148 19340 56160
rect 18463 56120 19340 56148
rect 18463 56117 18475 56120
rect 18417 56111 18475 56117
rect 19334 56108 19340 56120
rect 19392 56108 19398 56160
rect 20162 56148 20168 56160
rect 20123 56120 20168 56148
rect 20162 56108 20168 56120
rect 20220 56108 20226 56160
rect 21542 56108 21548 56160
rect 21600 56148 21606 56160
rect 23124 56148 23152 56256
rect 26973 56253 26985 56287
rect 27019 56284 27031 56287
rect 27154 56284 27160 56296
rect 27019 56256 27160 56284
rect 27019 56253 27031 56256
rect 26973 56247 27031 56253
rect 27154 56244 27160 56256
rect 27212 56244 27218 56296
rect 28552 56284 28580 56315
rect 28718 56312 28724 56324
rect 28776 56312 28782 56364
rect 28828 56361 28856 56460
rect 29178 56448 29184 56460
rect 29236 56448 29242 56500
rect 29730 56448 29736 56500
rect 29788 56488 29794 56500
rect 29914 56488 29920 56500
rect 29788 56460 29920 56488
rect 29788 56448 29794 56460
rect 29914 56448 29920 56460
rect 29972 56448 29978 56500
rect 29086 56380 29092 56432
rect 29144 56420 29150 56432
rect 29144 56392 29316 56420
rect 29144 56380 29150 56392
rect 29288 56361 29316 56392
rect 28813 56355 28871 56361
rect 28813 56321 28825 56355
rect 28859 56321 28871 56355
rect 28813 56315 28871 56321
rect 29273 56355 29331 56361
rect 29273 56321 29285 56355
rect 29319 56321 29331 56355
rect 29273 56315 29331 56321
rect 29549 56355 29607 56361
rect 29549 56321 29561 56355
rect 29595 56352 29607 56355
rect 30006 56352 30012 56364
rect 29595 56324 30012 56352
rect 29595 56321 29607 56324
rect 29549 56315 29607 56321
rect 30006 56312 30012 56324
rect 30064 56312 30070 56364
rect 29086 56284 29092 56296
rect 28552 56256 29092 56284
rect 29086 56244 29092 56256
rect 29144 56244 29150 56296
rect 24118 56216 24124 56228
rect 24079 56188 24124 56216
rect 24118 56176 24124 56188
rect 24176 56176 24182 56228
rect 27338 56176 27344 56228
rect 27396 56216 27402 56228
rect 30742 56216 30748 56228
rect 27396 56188 30748 56216
rect 27396 56176 27402 56188
rect 30742 56176 30748 56188
rect 30800 56216 30806 56228
rect 31570 56216 31576 56228
rect 30800 56188 31576 56216
rect 30800 56176 30806 56188
rect 31570 56176 31576 56188
rect 31628 56176 31634 56228
rect 21600 56120 23152 56148
rect 21600 56108 21606 56120
rect 24210 56108 24216 56160
rect 24268 56148 24274 56160
rect 26602 56148 26608 56160
rect 24268 56120 26608 56148
rect 24268 56108 24274 56120
rect 26602 56108 26608 56120
rect 26660 56108 26666 56160
rect 1104 56058 30820 56080
rect 1104 56006 5915 56058
rect 5967 56006 5979 56058
rect 6031 56006 6043 56058
rect 6095 56006 6107 56058
rect 6159 56006 6171 56058
rect 6223 56006 15846 56058
rect 15898 56006 15910 56058
rect 15962 56006 15974 56058
rect 16026 56006 16038 56058
rect 16090 56006 16102 56058
rect 16154 56006 25776 56058
rect 25828 56006 25840 56058
rect 25892 56006 25904 56058
rect 25956 56006 25968 56058
rect 26020 56006 26032 56058
rect 26084 56006 30820 56058
rect 1104 55984 30820 56006
rect 1394 55904 1400 55956
rect 1452 55944 1458 55956
rect 1673 55947 1731 55953
rect 1673 55944 1685 55947
rect 1452 55916 1685 55944
rect 1452 55904 1458 55916
rect 1673 55913 1685 55916
rect 1719 55913 1731 55947
rect 1673 55907 1731 55913
rect 2682 55904 2688 55956
rect 2740 55944 2746 55956
rect 15378 55944 15384 55956
rect 2740 55916 15384 55944
rect 2740 55904 2746 55916
rect 15378 55904 15384 55916
rect 15436 55904 15442 55956
rect 21085 55947 21143 55953
rect 21085 55913 21097 55947
rect 21131 55944 21143 55947
rect 21174 55944 21180 55956
rect 21131 55916 21180 55944
rect 21131 55913 21143 55916
rect 21085 55907 21143 55913
rect 21174 55904 21180 55916
rect 21232 55904 21238 55956
rect 21266 55904 21272 55956
rect 21324 55944 21330 55956
rect 23201 55947 23259 55953
rect 23201 55944 23213 55947
rect 21324 55916 23213 55944
rect 21324 55904 21330 55916
rect 23201 55913 23213 55916
rect 23247 55913 23259 55947
rect 24394 55944 24400 55956
rect 24355 55916 24400 55944
rect 23201 55907 23259 55913
rect 2314 55836 2320 55888
rect 2372 55876 2378 55888
rect 15194 55876 15200 55888
rect 2372 55848 15200 55876
rect 2372 55836 2378 55848
rect 15194 55836 15200 55848
rect 15252 55836 15258 55888
rect 15841 55879 15899 55885
rect 15841 55845 15853 55879
rect 15887 55876 15899 55879
rect 16298 55876 16304 55888
rect 15887 55848 16304 55876
rect 15887 55845 15899 55848
rect 15841 55839 15899 55845
rect 16298 55836 16304 55848
rect 16356 55836 16362 55888
rect 21818 55836 21824 55888
rect 21876 55836 21882 55888
rect 16206 55808 16212 55820
rect 16167 55780 16212 55808
rect 16206 55768 16212 55780
rect 16264 55768 16270 55820
rect 21836 55808 21864 55836
rect 23216 55808 23244 55907
rect 24394 55904 24400 55916
rect 24452 55904 24458 55956
rect 24486 55904 24492 55956
rect 24544 55904 24550 55956
rect 24578 55904 24584 55956
rect 24636 55944 24642 55956
rect 25682 55944 25688 55956
rect 24636 55916 25688 55944
rect 24636 55904 24642 55916
rect 25682 55904 25688 55916
rect 25740 55904 25746 55956
rect 30742 55904 30748 55956
rect 30800 55944 30806 55956
rect 31386 55944 31392 55956
rect 30800 55916 31392 55944
rect 30800 55904 30806 55916
rect 31386 55904 31392 55916
rect 31444 55904 31450 55956
rect 24504 55876 24532 55904
rect 24504 55848 25176 55876
rect 24394 55808 24400 55820
rect 21836 55780 21938 55808
rect 23216 55780 24400 55808
rect 1854 55740 1860 55752
rect 1815 55712 1860 55740
rect 1854 55700 1860 55712
rect 1912 55700 1918 55752
rect 18690 55700 18696 55752
rect 18748 55740 18754 55752
rect 21821 55743 21879 55749
rect 21821 55740 21833 55743
rect 18748 55712 21833 55740
rect 18748 55700 18754 55712
rect 21821 55709 21833 55712
rect 21867 55709 21879 55743
rect 21910 55740 21938 55780
rect 24394 55768 24400 55780
rect 24452 55768 24458 55820
rect 25041 55811 25099 55817
rect 25041 55777 25053 55811
rect 25087 55777 25099 55811
rect 25041 55771 25099 55777
rect 22077 55743 22135 55749
rect 22077 55740 22089 55743
rect 21910 55712 22089 55740
rect 21821 55703 21879 55709
rect 22077 55709 22089 55712
rect 22123 55709 22135 55743
rect 22077 55703 22135 55709
rect 22462 55700 22468 55752
rect 22520 55740 22526 55752
rect 23106 55740 23112 55752
rect 22520 55712 23112 55740
rect 22520 55700 22526 55712
rect 23106 55700 23112 55712
rect 23164 55700 23170 55752
rect 24578 55740 24584 55752
rect 24539 55712 24584 55740
rect 24578 55700 24584 55712
rect 24636 55700 24642 55752
rect 24673 55743 24731 55749
rect 24673 55709 24685 55743
rect 24719 55709 24731 55743
rect 24673 55703 24731 55709
rect 16393 55675 16451 55681
rect 16393 55641 16405 55675
rect 16439 55672 16451 55675
rect 16574 55672 16580 55684
rect 16439 55644 16580 55672
rect 16439 55641 16451 55644
rect 16393 55635 16451 55641
rect 16574 55632 16580 55644
rect 16632 55632 16638 55684
rect 16942 55672 16948 55684
rect 16903 55644 16948 55672
rect 16942 55632 16948 55644
rect 17000 55632 17006 55684
rect 19610 55672 19616 55684
rect 19571 55644 19616 55672
rect 19610 55632 19616 55644
rect 19668 55632 19674 55684
rect 22296 55644 24256 55672
rect 16301 55607 16359 55613
rect 16301 55573 16313 55607
rect 16347 55604 16359 55607
rect 17770 55604 17776 55616
rect 16347 55576 17776 55604
rect 16347 55573 16359 55576
rect 16301 55567 16359 55573
rect 17770 55564 17776 55576
rect 17828 55564 17834 55616
rect 18230 55604 18236 55616
rect 18191 55576 18236 55604
rect 18230 55564 18236 55576
rect 18288 55564 18294 55616
rect 21910 55564 21916 55616
rect 21968 55604 21974 55616
rect 22296 55604 22324 55644
rect 24228 55616 24256 55644
rect 24486 55632 24492 55684
rect 24544 55672 24550 55684
rect 24688 55672 24716 55703
rect 24544 55644 24716 55672
rect 25056 55672 25084 55771
rect 25148 55740 25176 55848
rect 30558 55836 30564 55888
rect 30616 55876 30622 55888
rect 31294 55876 31300 55888
rect 30616 55848 31300 55876
rect 30616 55836 30622 55848
rect 31294 55836 31300 55848
rect 31352 55836 31358 55888
rect 25958 55768 25964 55820
rect 26016 55768 26022 55820
rect 27157 55811 27215 55817
rect 27157 55777 27169 55811
rect 27203 55808 27215 55811
rect 27430 55808 27436 55820
rect 27203 55780 27436 55808
rect 27203 55777 27215 55780
rect 27157 55771 27215 55777
rect 27430 55768 27436 55780
rect 27488 55768 27494 55820
rect 28169 55811 28227 55817
rect 28169 55777 28181 55811
rect 28215 55808 28227 55811
rect 28902 55808 28908 55820
rect 28215 55780 28908 55808
rect 28215 55777 28227 55780
rect 28169 55771 28227 55777
rect 28902 55768 28908 55780
rect 28960 55768 28966 55820
rect 30650 55768 30656 55820
rect 30708 55808 30714 55820
rect 31662 55808 31668 55820
rect 30708 55780 31668 55808
rect 30708 55768 30714 55780
rect 31662 55768 31668 55780
rect 31720 55768 31726 55820
rect 25976 55740 26004 55768
rect 25148 55712 25820 55740
rect 25498 55672 25504 55684
rect 25056 55644 25360 55672
rect 25459 55644 25504 55672
rect 24544 55632 24550 55644
rect 25332 55616 25360 55644
rect 25498 55632 25504 55644
rect 25556 55632 25562 55684
rect 25682 55672 25688 55684
rect 25643 55644 25688 55672
rect 25682 55632 25688 55644
rect 25740 55632 25746 55684
rect 21968 55576 22324 55604
rect 21968 55564 21974 55576
rect 22554 55564 22560 55616
rect 22612 55604 22618 55616
rect 22738 55604 22744 55616
rect 22612 55576 22744 55604
rect 22612 55564 22618 55576
rect 22738 55564 22744 55576
rect 22796 55564 22802 55616
rect 24210 55564 24216 55616
rect 24268 55604 24274 55616
rect 24765 55607 24823 55613
rect 24765 55604 24777 55607
rect 24268 55576 24777 55604
rect 24268 55564 24274 55576
rect 24765 55573 24777 55576
rect 24811 55573 24823 55607
rect 24765 55567 24823 55573
rect 24949 55607 25007 55613
rect 24949 55573 24961 55607
rect 24995 55604 25007 55607
rect 25038 55604 25044 55616
rect 24995 55576 25044 55604
rect 24995 55573 25007 55576
rect 24949 55567 25007 55573
rect 25038 55564 25044 55576
rect 25096 55564 25102 55616
rect 25314 55564 25320 55616
rect 25372 55564 25378 55616
rect 25792 55613 25820 55712
rect 25884 55712 26004 55740
rect 26881 55743 26939 55749
rect 25884 55613 25912 55712
rect 26881 55709 26893 55743
rect 26927 55740 26939 55743
rect 28442 55740 28448 55752
rect 26927 55712 27200 55740
rect 28403 55712 28448 55740
rect 26927 55709 26939 55712
rect 26881 55703 26939 55709
rect 27172 55684 27200 55712
rect 28442 55700 28448 55712
rect 28500 55700 28506 55752
rect 25958 55632 25964 55684
rect 26016 55672 26022 55684
rect 26053 55675 26111 55681
rect 26053 55672 26065 55675
rect 26016 55644 26065 55672
rect 26016 55632 26022 55644
rect 26053 55641 26065 55644
rect 26099 55641 26111 55675
rect 26053 55635 26111 55641
rect 27154 55632 27160 55684
rect 27212 55632 27218 55684
rect 29730 55672 29736 55684
rect 29691 55644 29736 55672
rect 29730 55632 29736 55644
rect 29788 55632 29794 55684
rect 30101 55675 30159 55681
rect 30101 55641 30113 55675
rect 30147 55672 30159 55675
rect 30926 55672 30932 55684
rect 30147 55644 30932 55672
rect 30147 55641 30159 55644
rect 30101 55635 30159 55641
rect 30926 55632 30932 55644
rect 30984 55672 30990 55684
rect 31754 55672 31760 55684
rect 30984 55644 31760 55672
rect 30984 55632 30990 55644
rect 31754 55632 31760 55644
rect 31812 55632 31818 55684
rect 25777 55607 25835 55613
rect 25777 55573 25789 55607
rect 25823 55573 25835 55607
rect 25777 55567 25835 55573
rect 25869 55607 25927 55613
rect 25869 55573 25881 55607
rect 25915 55573 25927 55607
rect 25869 55567 25927 55573
rect 26510 55564 26516 55616
rect 26568 55604 26574 55616
rect 26786 55604 26792 55616
rect 26568 55576 26792 55604
rect 26568 55564 26574 55576
rect 26786 55564 26792 55576
rect 26844 55564 26850 55616
rect 28626 55564 28632 55616
rect 28684 55604 28690 55616
rect 29362 55604 29368 55616
rect 28684 55576 29368 55604
rect 28684 55564 28690 55576
rect 29362 55564 29368 55576
rect 29420 55564 29426 55616
rect 1104 55514 30820 55536
rect 1104 55462 10880 55514
rect 10932 55462 10944 55514
rect 10996 55462 11008 55514
rect 11060 55462 11072 55514
rect 11124 55462 11136 55514
rect 11188 55462 20811 55514
rect 20863 55462 20875 55514
rect 20927 55462 20939 55514
rect 20991 55462 21003 55514
rect 21055 55462 21067 55514
rect 21119 55462 30820 55514
rect 1104 55440 30820 55462
rect 2130 55400 2136 55412
rect 2091 55372 2136 55400
rect 2130 55360 2136 55372
rect 2188 55360 2194 55412
rect 16574 55360 16580 55412
rect 16632 55400 16638 55412
rect 17310 55400 17316 55412
rect 16632 55372 17316 55400
rect 16632 55360 16638 55372
rect 17310 55360 17316 55372
rect 17368 55360 17374 55412
rect 17954 55360 17960 55412
rect 18012 55400 18018 55412
rect 18049 55403 18107 55409
rect 18049 55400 18061 55403
rect 18012 55372 18061 55400
rect 18012 55360 18018 55372
rect 18049 55369 18061 55372
rect 18095 55369 18107 55403
rect 18049 55363 18107 55369
rect 18874 55360 18880 55412
rect 18932 55400 18938 55412
rect 18932 55372 20208 55400
rect 18932 55360 18938 55372
rect 16117 55335 16175 55341
rect 16117 55301 16129 55335
rect 16163 55332 16175 55335
rect 16206 55332 16212 55344
rect 16163 55304 16212 55332
rect 16163 55301 16175 55304
rect 16117 55295 16175 55301
rect 16206 55292 16212 55304
rect 16264 55292 16270 55344
rect 18322 55332 18328 55344
rect 17144 55304 18328 55332
rect 1394 55264 1400 55276
rect 1355 55236 1400 55264
rect 1394 55224 1400 55236
rect 1452 55224 1458 55276
rect 2317 55267 2375 55273
rect 2317 55233 2329 55267
rect 2363 55264 2375 55267
rect 4798 55264 4804 55276
rect 2363 55236 4804 55264
rect 2363 55233 2375 55236
rect 2317 55227 2375 55233
rect 4798 55224 4804 55236
rect 4856 55224 4862 55276
rect 15933 55267 15991 55273
rect 15933 55233 15945 55267
rect 15979 55264 15991 55267
rect 17144 55264 17172 55304
rect 18322 55292 18328 55304
rect 18380 55292 18386 55344
rect 15979 55236 17172 55264
rect 15979 55233 15991 55236
rect 15933 55227 15991 55233
rect 17218 55224 17224 55276
rect 17276 55264 17282 55276
rect 17276 55236 17321 55264
rect 17276 55224 17282 55236
rect 17678 55224 17684 55276
rect 17736 55264 17742 55276
rect 17865 55267 17923 55273
rect 17865 55264 17877 55267
rect 17736 55236 17877 55264
rect 17736 55224 17742 55236
rect 17865 55233 17877 55236
rect 17911 55233 17923 55267
rect 19794 55264 19800 55276
rect 19755 55236 19800 55264
rect 17865 55227 17923 55233
rect 19794 55224 19800 55236
rect 19852 55224 19858 55276
rect 20180 55273 20208 55372
rect 20714 55360 20720 55412
rect 20772 55400 20778 55412
rect 20809 55403 20867 55409
rect 20809 55400 20821 55403
rect 20772 55372 20821 55400
rect 20772 55360 20778 55372
rect 20809 55369 20821 55372
rect 20855 55369 20867 55403
rect 20809 55363 20867 55369
rect 23106 55360 23112 55412
rect 23164 55400 23170 55412
rect 23658 55400 23664 55412
rect 23164 55372 23664 55400
rect 23164 55360 23170 55372
rect 23658 55360 23664 55372
rect 23716 55400 23722 55412
rect 24581 55403 24639 55409
rect 24581 55400 24593 55403
rect 23716 55372 24593 55400
rect 23716 55360 23722 55372
rect 24581 55369 24593 55372
rect 24627 55369 24639 55403
rect 24581 55363 24639 55369
rect 24946 55360 24952 55412
rect 25004 55400 25010 55412
rect 25317 55403 25375 55409
rect 25317 55400 25329 55403
rect 25004 55372 25329 55400
rect 25004 55360 25010 55372
rect 25317 55369 25329 55372
rect 25363 55369 25375 55403
rect 25774 55400 25780 55412
rect 25735 55372 25780 55400
rect 25317 55363 25375 55369
rect 25774 55360 25780 55372
rect 25832 55360 25838 55412
rect 26973 55403 27031 55409
rect 26973 55369 26985 55403
rect 27019 55400 27031 55403
rect 27522 55400 27528 55412
rect 27019 55372 27528 55400
rect 27019 55369 27031 55372
rect 26973 55363 27031 55369
rect 27522 55360 27528 55372
rect 27580 55360 27586 55412
rect 29178 55400 29184 55412
rect 28184 55372 29184 55400
rect 25406 55332 25412 55344
rect 23584 55304 25412 55332
rect 19889 55267 19947 55273
rect 19889 55233 19901 55267
rect 19935 55233 19947 55267
rect 19889 55227 19947 55233
rect 19981 55267 20039 55273
rect 19981 55233 19993 55267
rect 20027 55233 20039 55267
rect 19981 55227 20039 55233
rect 20165 55267 20223 55273
rect 20165 55233 20177 55267
rect 20211 55233 20223 55267
rect 20165 55227 20223 55233
rect 20717 55267 20775 55273
rect 20717 55233 20729 55267
rect 20763 55264 20775 55267
rect 21266 55264 21272 55276
rect 20763 55236 21272 55264
rect 20763 55233 20775 55236
rect 20717 55227 20775 55233
rect 19702 55156 19708 55208
rect 19760 55196 19766 55208
rect 19901 55196 19929 55227
rect 19760 55168 19929 55196
rect 19996 55196 20024 55227
rect 21266 55224 21272 55236
rect 21324 55224 21330 55276
rect 22465 55267 22523 55273
rect 22465 55233 22477 55267
rect 22511 55264 22523 55267
rect 23290 55264 23296 55276
rect 22511 55236 23296 55264
rect 22511 55233 22523 55236
rect 22465 55227 22523 55233
rect 23290 55224 23296 55236
rect 23348 55224 23354 55276
rect 23584 55273 23612 55304
rect 25406 55292 25412 55304
rect 25464 55292 25470 55344
rect 25866 55332 25872 55344
rect 25827 55304 25872 55332
rect 25866 55292 25872 55304
rect 25924 55292 25930 55344
rect 26418 55292 26424 55344
rect 26476 55332 26482 55344
rect 27341 55335 27399 55341
rect 27341 55332 27353 55335
rect 26476 55304 27353 55332
rect 26476 55292 26482 55304
rect 27341 55301 27353 55304
rect 27387 55301 27399 55335
rect 27341 55295 27399 55301
rect 23569 55267 23627 55273
rect 23569 55233 23581 55267
rect 23615 55233 23627 55267
rect 23569 55227 23627 55233
rect 23661 55267 23719 55273
rect 23661 55233 23673 55267
rect 23707 55264 23719 55267
rect 24213 55267 24271 55273
rect 24213 55264 24225 55267
rect 23707 55236 24225 55264
rect 23707 55233 23719 55236
rect 23661 55227 23719 55233
rect 24213 55233 24225 55236
rect 24259 55233 24271 55267
rect 24213 55227 24271 55233
rect 24397 55267 24455 55273
rect 24397 55233 24409 55267
rect 24443 55264 24455 55267
rect 24578 55264 24584 55276
rect 24443 55236 24584 55264
rect 24443 55233 24455 55236
rect 24397 55227 24455 55233
rect 24578 55224 24584 55236
rect 24636 55264 24642 55276
rect 28184 55273 28212 55372
rect 29178 55360 29184 55372
rect 29236 55360 29242 55412
rect 30101 55403 30159 55409
rect 30101 55369 30113 55403
rect 30147 55400 30159 55403
rect 30282 55400 30288 55412
rect 30147 55372 30288 55400
rect 30147 55369 30159 55372
rect 30101 55363 30159 55369
rect 30282 55360 30288 55372
rect 30340 55360 30346 55412
rect 28442 55292 28448 55344
rect 28500 55332 28506 55344
rect 30926 55332 30932 55344
rect 28500 55304 29592 55332
rect 28500 55292 28506 55304
rect 25501 55267 25559 55273
rect 25501 55264 25513 55267
rect 24636 55236 25513 55264
rect 24636 55224 24642 55236
rect 25501 55233 25513 55236
rect 25547 55233 25559 55267
rect 25501 55227 25559 55233
rect 27157 55267 27215 55273
rect 27157 55233 27169 55267
rect 27203 55233 27215 55267
rect 27157 55227 27215 55233
rect 27433 55267 27491 55273
rect 27433 55233 27445 55267
rect 27479 55233 27491 55267
rect 27433 55227 27491 55233
rect 28169 55267 28227 55273
rect 28169 55233 28181 55267
rect 28215 55233 28227 55267
rect 28169 55227 28227 55233
rect 28353 55267 28411 55273
rect 28353 55233 28365 55267
rect 28399 55264 28411 55267
rect 28626 55264 28632 55276
rect 28399 55236 28632 55264
rect 28399 55233 28411 55236
rect 28353 55227 28411 55233
rect 20254 55196 20260 55208
rect 19996 55168 20260 55196
rect 19760 55156 19766 55168
rect 20254 55156 20260 55168
rect 20312 55156 20318 55208
rect 20622 55156 20628 55208
rect 20680 55196 20686 55208
rect 22281 55199 22339 55205
rect 22281 55196 22293 55199
rect 20680 55168 22293 55196
rect 20680 55156 20686 55168
rect 22281 55165 22293 55168
rect 22327 55165 22339 55199
rect 22281 55159 22339 55165
rect 22649 55199 22707 55205
rect 22649 55165 22661 55199
rect 22695 55196 22707 55199
rect 23198 55196 23204 55208
rect 22695 55168 23204 55196
rect 22695 55165 22707 55168
rect 22649 55159 22707 55165
rect 23198 55156 23204 55168
rect 23256 55156 23262 55208
rect 23385 55199 23443 55205
rect 23385 55165 23397 55199
rect 23431 55165 23443 55199
rect 23385 55159 23443 55165
rect 23477 55199 23535 55205
rect 23477 55165 23489 55199
rect 23523 55196 23535 55199
rect 24486 55196 24492 55208
rect 23523 55168 23796 55196
rect 24447 55168 24492 55196
rect 23523 55165 23535 55168
rect 23477 55159 23535 55165
rect 1578 55128 1584 55140
rect 1539 55100 1584 55128
rect 1578 55088 1584 55100
rect 1636 55088 1642 55140
rect 23400 55128 23428 55159
rect 23658 55128 23664 55140
rect 23400 55100 23664 55128
rect 23658 55088 23664 55100
rect 23716 55088 23722 55140
rect 14642 55020 14648 55072
rect 14700 55060 14706 55072
rect 18782 55060 18788 55072
rect 14700 55032 18788 55060
rect 14700 55020 14706 55032
rect 18782 55020 18788 55032
rect 18840 55020 18846 55072
rect 19521 55063 19579 55069
rect 19521 55029 19533 55063
rect 19567 55060 19579 55063
rect 19794 55060 19800 55072
rect 19567 55032 19800 55060
rect 19567 55029 19579 55032
rect 19521 55023 19579 55029
rect 19794 55020 19800 55032
rect 19852 55020 19858 55072
rect 23198 55060 23204 55072
rect 23159 55032 23204 55060
rect 23198 55020 23204 55032
rect 23256 55020 23262 55072
rect 23566 55020 23572 55072
rect 23624 55060 23630 55072
rect 23768 55060 23796 55168
rect 24486 55156 24492 55168
rect 24544 55156 24550 55208
rect 24765 55199 24823 55205
rect 24765 55196 24777 55199
rect 24688 55168 24777 55196
rect 24210 55088 24216 55140
rect 24268 55128 24274 55140
rect 24688 55128 24716 55168
rect 24765 55165 24777 55168
rect 24811 55165 24823 55199
rect 24765 55159 24823 55165
rect 24857 55199 24915 55205
rect 24857 55165 24869 55199
rect 24903 55196 24915 55199
rect 25038 55196 25044 55208
rect 24903 55168 25044 55196
rect 24903 55165 24915 55168
rect 24857 55159 24915 55165
rect 25038 55156 25044 55168
rect 25096 55196 25102 55208
rect 25314 55196 25320 55208
rect 25096 55168 25320 55196
rect 25096 55156 25102 55168
rect 25314 55156 25320 55168
rect 25372 55156 25378 55208
rect 25593 55199 25651 55205
rect 25593 55165 25605 55199
rect 25639 55196 25651 55199
rect 25961 55199 26019 55205
rect 25961 55196 25973 55199
rect 25639 55168 25728 55196
rect 25639 55165 25651 55168
rect 25593 55159 25651 55165
rect 24268 55100 24716 55128
rect 24268 55088 24274 55100
rect 25222 55088 25228 55140
rect 25280 55128 25286 55140
rect 25700 55128 25728 55168
rect 25280 55100 25728 55128
rect 25792 55168 25973 55196
rect 25280 55088 25286 55100
rect 23624 55032 23796 55060
rect 23624 55020 23630 55032
rect 25314 55020 25320 55072
rect 25372 55060 25378 55072
rect 25792 55060 25820 55168
rect 25961 55165 25973 55168
rect 26007 55165 26019 55199
rect 25961 55159 26019 55165
rect 27172 55128 27200 55227
rect 27338 55128 27344 55140
rect 27172 55100 27344 55128
rect 27338 55088 27344 55100
rect 27396 55088 27402 55140
rect 25372 55032 25820 55060
rect 25372 55020 25378 55032
rect 26234 55020 26240 55072
rect 26292 55060 26298 55072
rect 27448 55060 27476 55227
rect 28626 55224 28632 55236
rect 28684 55224 28690 55276
rect 28721 55267 28779 55273
rect 28721 55233 28733 55267
rect 28767 55233 28779 55267
rect 28721 55227 28779 55233
rect 28445 55199 28503 55205
rect 28445 55165 28457 55199
rect 28491 55165 28503 55199
rect 28445 55159 28503 55165
rect 28537 55199 28595 55205
rect 28537 55165 28549 55199
rect 28583 55165 28595 55199
rect 28537 55159 28595 55165
rect 28166 55088 28172 55140
rect 28224 55128 28230 55140
rect 28460 55128 28488 55159
rect 28224 55100 28488 55128
rect 28224 55088 28230 55100
rect 26292 55032 27476 55060
rect 28552 55060 28580 55159
rect 28626 55060 28632 55072
rect 28552 55032 28632 55060
rect 26292 55020 26298 55032
rect 28626 55020 28632 55032
rect 28684 55020 28690 55072
rect 28736 55060 28764 55227
rect 28810 55224 28816 55276
rect 28868 55264 28874 55276
rect 29564 55273 29592 55304
rect 29656 55304 30932 55332
rect 29656 55273 29684 55304
rect 30926 55292 30932 55304
rect 30984 55292 30990 55344
rect 29365 55267 29423 55273
rect 29365 55266 29377 55267
rect 29288 55264 29377 55266
rect 28868 55238 29377 55264
rect 28868 55236 29316 55238
rect 28868 55224 28874 55236
rect 29365 55233 29377 55238
rect 29411 55233 29423 55267
rect 29365 55227 29423 55233
rect 29549 55267 29607 55273
rect 29549 55233 29561 55267
rect 29595 55233 29607 55267
rect 29549 55227 29607 55233
rect 29641 55267 29699 55273
rect 29641 55233 29653 55267
rect 29687 55233 29699 55267
rect 29641 55227 29699 55233
rect 29917 55267 29975 55273
rect 29917 55233 29929 55267
rect 29963 55264 29975 55267
rect 30006 55264 30012 55276
rect 29963 55236 30012 55264
rect 29963 55233 29975 55236
rect 29917 55227 29975 55233
rect 30006 55224 30012 55236
rect 30064 55224 30070 55276
rect 29733 55199 29791 55205
rect 29733 55165 29745 55199
rect 29779 55196 29791 55199
rect 31662 55196 31668 55208
rect 29779 55168 31668 55196
rect 29779 55165 29791 55168
rect 29733 55159 29791 55165
rect 31662 55156 31668 55168
rect 31720 55156 31726 55208
rect 28905 55131 28963 55137
rect 28905 55097 28917 55131
rect 28951 55128 28963 55131
rect 30834 55128 30840 55140
rect 28951 55100 30840 55128
rect 28951 55097 28963 55100
rect 28905 55091 28963 55097
rect 30834 55088 30840 55100
rect 30892 55088 30898 55140
rect 30006 55060 30012 55072
rect 28736 55032 30012 55060
rect 30006 55020 30012 55032
rect 30064 55020 30070 55072
rect 1104 54970 30820 54992
rect 1104 54918 5915 54970
rect 5967 54918 5979 54970
rect 6031 54918 6043 54970
rect 6095 54918 6107 54970
rect 6159 54918 6171 54970
rect 6223 54918 15846 54970
rect 15898 54918 15910 54970
rect 15962 54918 15974 54970
rect 16026 54918 16038 54970
rect 16090 54918 16102 54970
rect 16154 54918 25776 54970
rect 25828 54918 25840 54970
rect 25892 54918 25904 54970
rect 25956 54918 25968 54970
rect 26020 54918 26032 54970
rect 26084 54918 30820 54970
rect 1104 54896 30820 54918
rect 15470 54816 15476 54868
rect 15528 54856 15534 54868
rect 15841 54859 15899 54865
rect 15841 54856 15853 54859
rect 15528 54828 15853 54856
rect 15528 54816 15534 54828
rect 15841 54825 15853 54828
rect 15887 54825 15899 54859
rect 21818 54856 21824 54868
rect 15841 54819 15899 54825
rect 15948 54828 21824 54856
rect 13354 54748 13360 54800
rect 13412 54788 13418 54800
rect 15948 54788 15976 54828
rect 21818 54816 21824 54828
rect 21876 54816 21882 54868
rect 23658 54816 23664 54868
rect 23716 54856 23722 54868
rect 24578 54856 24584 54868
rect 23716 54828 24584 54856
rect 23716 54816 23722 54828
rect 24578 54816 24584 54828
rect 24636 54865 24642 54868
rect 24636 54859 24685 54865
rect 24636 54825 24639 54859
rect 24673 54825 24685 54859
rect 24636 54819 24685 54825
rect 25961 54859 26019 54865
rect 25961 54825 25973 54859
rect 26007 54856 26019 54859
rect 26142 54856 26148 54868
rect 26007 54828 26148 54856
rect 26007 54825 26019 54828
rect 25961 54819 26019 54825
rect 24636 54816 24642 54819
rect 26142 54816 26148 54828
rect 26200 54816 26206 54868
rect 26970 54816 26976 54868
rect 27028 54856 27034 54868
rect 27893 54859 27951 54865
rect 27893 54856 27905 54859
rect 27028 54828 27905 54856
rect 27028 54816 27034 54828
rect 27893 54825 27905 54828
rect 27939 54825 27951 54859
rect 27893 54819 27951 54825
rect 28626 54816 28632 54868
rect 28684 54856 28690 54868
rect 30374 54856 30380 54868
rect 28684 54828 30380 54856
rect 28684 54816 28690 54828
rect 30374 54816 30380 54828
rect 30432 54856 30438 54868
rect 31202 54856 31208 54868
rect 30432 54828 31208 54856
rect 30432 54816 30438 54828
rect 31202 54816 31208 54828
rect 31260 54816 31266 54868
rect 13412 54760 15976 54788
rect 13412 54748 13418 54760
rect 17402 54748 17408 54800
rect 17460 54788 17466 54800
rect 22646 54788 22652 54800
rect 17460 54760 22652 54788
rect 17460 54748 17466 54760
rect 22646 54748 22652 54760
rect 22704 54788 22710 54800
rect 26050 54788 26056 54800
rect 22704 54760 26056 54788
rect 22704 54748 22710 54760
rect 26050 54748 26056 54760
rect 26108 54748 26114 54800
rect 27430 54748 27436 54800
rect 27488 54788 27494 54800
rect 28813 54791 28871 54797
rect 28813 54788 28825 54791
rect 27488 54760 28825 54788
rect 27488 54748 27494 54760
rect 28813 54757 28825 54760
rect 28859 54757 28871 54791
rect 28813 54751 28871 54757
rect 20438 54720 20444 54732
rect 6886 54692 20444 54720
rect 1397 54655 1455 54661
rect 1397 54621 1409 54655
rect 1443 54652 1455 54655
rect 2130 54652 2136 54664
rect 1443 54624 2136 54652
rect 1443 54621 1455 54624
rect 1397 54615 1455 54621
rect 2130 54612 2136 54624
rect 2188 54612 2194 54664
rect 2590 54544 2596 54596
rect 2648 54584 2654 54596
rect 6886 54584 6914 54692
rect 20438 54680 20444 54692
rect 20496 54680 20502 54732
rect 23658 54680 23664 54732
rect 23716 54720 23722 54732
rect 24026 54720 24032 54732
rect 23716 54692 24032 54720
rect 23716 54680 23722 54692
rect 24026 54680 24032 54692
rect 24084 54720 24090 54732
rect 24397 54723 24455 54729
rect 24397 54720 24409 54723
rect 24084 54692 24409 54720
rect 24084 54680 24090 54692
rect 24397 54689 24409 54692
rect 24443 54689 24455 54723
rect 24397 54683 24455 54689
rect 26970 54680 26976 54732
rect 27028 54720 27034 54732
rect 30009 54723 30067 54729
rect 30009 54720 30021 54723
rect 27028 54692 30021 54720
rect 27028 54680 27034 54692
rect 30009 54689 30021 54692
rect 30055 54720 30067 54723
rect 30926 54720 30932 54732
rect 30055 54692 30932 54720
rect 30055 54689 30067 54692
rect 30009 54683 30067 54689
rect 30926 54680 30932 54692
rect 30984 54680 30990 54732
rect 15657 54655 15715 54661
rect 15657 54621 15669 54655
rect 15703 54621 15715 54655
rect 16298 54652 16304 54664
rect 16259 54624 16304 54652
rect 15657 54615 15715 54621
rect 2648 54556 6914 54584
rect 15672 54584 15700 54615
rect 16298 54612 16304 54624
rect 16356 54612 16362 54664
rect 26145 54655 26203 54661
rect 26145 54621 26157 54655
rect 26191 54621 26203 54655
rect 26145 54615 26203 54621
rect 17034 54584 17040 54596
rect 15672 54556 17040 54584
rect 2648 54544 2654 54556
rect 17034 54544 17040 54556
rect 17092 54544 17098 54596
rect 22094 54544 22100 54596
rect 22152 54584 22158 54596
rect 26160 54584 26188 54615
rect 26234 54612 26240 54664
rect 26292 54652 26298 54664
rect 26421 54655 26479 54661
rect 26421 54652 26433 54655
rect 26292 54624 26433 54652
rect 26292 54612 26298 54624
rect 26421 54621 26433 54624
rect 26467 54621 26479 54655
rect 26421 54615 26479 54621
rect 27525 54655 27583 54661
rect 27525 54621 27537 54655
rect 27571 54652 27583 54655
rect 29730 54652 29736 54664
rect 27571 54624 28994 54652
rect 29691 54624 29736 54652
rect 27571 54621 27583 54624
rect 27525 54615 27583 54621
rect 27338 54584 27344 54596
rect 22152 54556 22197 54584
rect 26160 54556 27344 54584
rect 22152 54544 22158 54556
rect 27338 54544 27344 54556
rect 27396 54544 27402 54596
rect 27614 54544 27620 54596
rect 27672 54584 27678 54596
rect 27709 54587 27767 54593
rect 27709 54584 27721 54587
rect 27672 54556 27721 54584
rect 27672 54544 27678 54556
rect 27709 54553 27721 54556
rect 27755 54553 27767 54587
rect 28626 54584 28632 54596
rect 28587 54556 28632 54584
rect 27709 54547 27767 54553
rect 28626 54544 28632 54556
rect 28684 54544 28690 54596
rect 28966 54584 28994 54624
rect 29730 54612 29736 54624
rect 29788 54612 29794 54664
rect 30374 54612 30380 54664
rect 30432 54652 30438 54664
rect 31294 54652 31300 54664
rect 30432 54624 31300 54652
rect 30432 54612 30438 54624
rect 31294 54612 31300 54624
rect 31352 54612 31358 54664
rect 30282 54584 30288 54596
rect 28966 54556 30288 54584
rect 30282 54544 30288 54556
rect 30340 54544 30346 54596
rect 1578 54516 1584 54528
rect 1539 54488 1584 54516
rect 1578 54476 1584 54488
rect 1636 54476 1642 54528
rect 16485 54519 16543 54525
rect 16485 54485 16497 54519
rect 16531 54516 16543 54519
rect 16666 54516 16672 54528
rect 16531 54488 16672 54516
rect 16531 54485 16543 54488
rect 16485 54479 16543 54485
rect 16666 54476 16672 54488
rect 16724 54476 16730 54528
rect 22278 54476 22284 54528
rect 22336 54516 22342 54528
rect 23382 54516 23388 54528
rect 22336 54488 23388 54516
rect 22336 54476 22342 54488
rect 23382 54476 23388 54488
rect 23440 54476 23446 54528
rect 24210 54476 24216 54528
rect 24268 54516 24274 54528
rect 26142 54516 26148 54528
rect 24268 54488 26148 54516
rect 24268 54476 24274 54488
rect 26142 54476 26148 54488
rect 26200 54516 26206 54528
rect 26329 54519 26387 54525
rect 26329 54516 26341 54519
rect 26200 54488 26341 54516
rect 26200 54476 26206 54488
rect 26329 54485 26341 54488
rect 26375 54485 26387 54519
rect 26329 54479 26387 54485
rect 28166 54476 28172 54528
rect 28224 54516 28230 54528
rect 31294 54516 31300 54528
rect 28224 54488 31300 54516
rect 28224 54476 28230 54488
rect 31294 54476 31300 54488
rect 31352 54476 31358 54528
rect 1104 54426 30820 54448
rect 1104 54374 10880 54426
rect 10932 54374 10944 54426
rect 10996 54374 11008 54426
rect 11060 54374 11072 54426
rect 11124 54374 11136 54426
rect 11188 54374 20811 54426
rect 20863 54374 20875 54426
rect 20927 54374 20939 54426
rect 20991 54374 21003 54426
rect 21055 54374 21067 54426
rect 21119 54374 30820 54426
rect 1104 54352 30820 54374
rect 1394 54272 1400 54324
rect 1452 54312 1458 54324
rect 2133 54315 2191 54321
rect 2133 54312 2145 54315
rect 1452 54284 2145 54312
rect 1452 54272 1458 54284
rect 2133 54281 2145 54284
rect 2179 54281 2191 54315
rect 2133 54275 2191 54281
rect 17402 54272 17408 54324
rect 17460 54312 17466 54324
rect 18049 54315 18107 54321
rect 18049 54312 18061 54315
rect 17460 54284 18061 54312
rect 17460 54272 17466 54284
rect 18049 54281 18061 54284
rect 18095 54281 18107 54315
rect 18049 54275 18107 54281
rect 19886 54272 19892 54324
rect 19944 54312 19950 54324
rect 21085 54315 21143 54321
rect 21085 54312 21097 54315
rect 19944 54284 21097 54312
rect 19944 54272 19950 54284
rect 21085 54281 21097 54284
rect 21131 54312 21143 54315
rect 25314 54312 25320 54324
rect 21131 54284 25320 54312
rect 21131 54281 21143 54284
rect 21085 54275 21143 54281
rect 25314 54272 25320 54284
rect 25372 54272 25378 54324
rect 27338 54272 27344 54324
rect 27396 54312 27402 54324
rect 27396 54284 28488 54312
rect 27396 54272 27402 54284
rect 16850 54204 16856 54256
rect 16908 54253 16914 54256
rect 16908 54247 16972 54253
rect 16908 54213 16926 54247
rect 16960 54213 16972 54247
rect 16908 54207 16972 54213
rect 16908 54204 16914 54207
rect 19334 54204 19340 54256
rect 19392 54244 19398 54256
rect 19392 54216 22094 54244
rect 19392 54204 19398 54216
rect 1394 54176 1400 54188
rect 1355 54148 1400 54176
rect 1394 54136 1400 54148
rect 1452 54136 1458 54188
rect 2317 54179 2375 54185
rect 2317 54145 2329 54179
rect 2363 54176 2375 54179
rect 7558 54176 7564 54188
rect 2363 54148 7564 54176
rect 2363 54145 2375 54148
rect 2317 54139 2375 54145
rect 7558 54136 7564 54148
rect 7616 54136 7622 54188
rect 16666 54176 16672 54188
rect 16627 54148 16672 54176
rect 16666 54136 16672 54148
rect 16724 54136 16730 54188
rect 19794 54136 19800 54188
rect 19852 54176 19858 54188
rect 19961 54179 20019 54185
rect 19961 54176 19973 54179
rect 19852 54148 19973 54176
rect 19852 54136 19858 54148
rect 19961 54145 19973 54148
rect 20007 54145 20019 54179
rect 22066 54176 22094 54216
rect 22830 54204 22836 54256
rect 22888 54244 22894 54256
rect 28460 54253 28488 54284
rect 29362 54272 29368 54324
rect 29420 54272 29426 54324
rect 29454 54272 29460 54324
rect 29512 54312 29518 54324
rect 30101 54315 30159 54321
rect 29512 54284 29684 54312
rect 29512 54272 29518 54284
rect 28445 54247 28503 54253
rect 22888 54216 27844 54244
rect 22888 54204 22894 54216
rect 23109 54179 23167 54185
rect 23109 54176 23121 54179
rect 22066 54148 23121 54176
rect 19961 54139 20019 54145
rect 23109 54145 23121 54148
rect 23155 54145 23167 54179
rect 23290 54176 23296 54188
rect 23251 54148 23296 54176
rect 23109 54139 23167 54145
rect 23290 54136 23296 54148
rect 23348 54136 23354 54188
rect 25222 54176 25228 54188
rect 25183 54148 25228 54176
rect 25222 54136 25228 54148
rect 25280 54136 25286 54188
rect 27430 54136 27436 54188
rect 27488 54176 27494 54188
rect 27525 54179 27583 54185
rect 27525 54176 27537 54179
rect 27488 54148 27537 54176
rect 27488 54136 27494 54148
rect 27525 54145 27537 54148
rect 27571 54145 27583 54179
rect 27525 54139 27583 54145
rect 27709 54179 27767 54185
rect 27709 54145 27721 54179
rect 27755 54145 27767 54179
rect 27709 54139 27767 54145
rect 19702 54108 19708 54120
rect 19663 54080 19708 54108
rect 19702 54068 19708 54080
rect 19760 54068 19766 54120
rect 25038 54068 25044 54120
rect 25096 54108 25102 54120
rect 27614 54108 27620 54120
rect 25096 54080 27620 54108
rect 25096 54068 25102 54080
rect 27614 54068 27620 54080
rect 27672 54108 27678 54120
rect 27724 54108 27752 54139
rect 27672 54080 27752 54108
rect 27816 54108 27844 54216
rect 28445 54213 28457 54247
rect 28491 54213 28503 54247
rect 29380 54244 29408 54272
rect 29380 54216 29592 54244
rect 28445 54207 28503 54213
rect 29362 54176 29368 54188
rect 29323 54148 29368 54176
rect 29362 54136 29368 54148
rect 29420 54136 29426 54188
rect 29564 54185 29592 54216
rect 29549 54179 29607 54185
rect 29549 54145 29561 54179
rect 29595 54145 29607 54179
rect 29656 54176 29684 54284
rect 30101 54281 30113 54315
rect 30147 54312 30159 54315
rect 30190 54312 30196 54324
rect 30147 54284 30196 54312
rect 30147 54281 30159 54284
rect 30101 54275 30159 54281
rect 30190 54272 30196 54284
rect 30248 54272 30254 54324
rect 29733 54179 29791 54185
rect 29733 54176 29745 54179
rect 29656 54148 29745 54176
rect 29549 54139 29607 54145
rect 29733 54145 29745 54148
rect 29779 54145 29791 54179
rect 29733 54139 29791 54145
rect 29917 54179 29975 54185
rect 29917 54145 29929 54179
rect 29963 54176 29975 54179
rect 30006 54176 30012 54188
rect 29963 54148 30012 54176
rect 29963 54145 29975 54148
rect 29917 54139 29975 54145
rect 29641 54111 29699 54117
rect 29641 54108 29653 54111
rect 27816 54080 29653 54108
rect 27672 54068 27678 54080
rect 29641 54077 29653 54080
rect 29687 54077 29699 54111
rect 29748 54108 29776 54139
rect 30006 54136 30012 54148
rect 30064 54136 30070 54188
rect 31386 54108 31392 54120
rect 29748 54080 31392 54108
rect 29641 54071 29699 54077
rect 31386 54068 31392 54080
rect 31444 54068 31450 54120
rect 28629 54043 28687 54049
rect 28629 54009 28641 54043
rect 28675 54040 28687 54043
rect 29086 54040 29092 54052
rect 28675 54012 29092 54040
rect 28675 54009 28687 54012
rect 28629 54003 28687 54009
rect 29086 54000 29092 54012
rect 29144 54040 29150 54052
rect 30282 54040 30288 54052
rect 29144 54012 30288 54040
rect 29144 54000 29150 54012
rect 30282 54000 30288 54012
rect 30340 54000 30346 54052
rect 1578 53972 1584 53984
rect 1539 53944 1584 53972
rect 1578 53932 1584 53944
rect 1636 53932 1642 53984
rect 23477 53975 23535 53981
rect 23477 53941 23489 53975
rect 23523 53972 23535 53975
rect 24026 53972 24032 53984
rect 23523 53944 24032 53972
rect 23523 53941 23535 53944
rect 23477 53935 23535 53941
rect 24026 53932 24032 53944
rect 24084 53932 24090 53984
rect 24486 53932 24492 53984
rect 24544 53972 24550 53984
rect 25317 53975 25375 53981
rect 25317 53972 25329 53975
rect 24544 53944 25329 53972
rect 24544 53932 24550 53944
rect 25317 53941 25329 53944
rect 25363 53941 25375 53975
rect 25317 53935 25375 53941
rect 27154 53932 27160 53984
rect 27212 53972 27218 53984
rect 27617 53975 27675 53981
rect 27617 53972 27629 53975
rect 27212 53944 27629 53972
rect 27212 53932 27218 53944
rect 27617 53941 27629 53944
rect 27663 53941 27675 53975
rect 27617 53935 27675 53941
rect 29638 53932 29644 53984
rect 29696 53972 29702 53984
rect 30190 53972 30196 53984
rect 29696 53944 30196 53972
rect 29696 53932 29702 53944
rect 30190 53932 30196 53944
rect 30248 53932 30254 53984
rect 1104 53882 30820 53904
rect 1104 53830 5915 53882
rect 5967 53830 5979 53882
rect 6031 53830 6043 53882
rect 6095 53830 6107 53882
rect 6159 53830 6171 53882
rect 6223 53830 15846 53882
rect 15898 53830 15910 53882
rect 15962 53830 15974 53882
rect 16026 53830 16038 53882
rect 16090 53830 16102 53882
rect 16154 53830 25776 53882
rect 25828 53830 25840 53882
rect 25892 53830 25904 53882
rect 25956 53830 25968 53882
rect 26020 53830 26032 53882
rect 26084 53830 30820 53882
rect 1104 53808 30820 53830
rect 2130 53768 2136 53780
rect 2091 53740 2136 53768
rect 2130 53728 2136 53740
rect 2188 53728 2194 53780
rect 18046 53768 18052 53780
rect 18007 53740 18052 53768
rect 18046 53728 18052 53740
rect 18104 53728 18110 53780
rect 18690 53768 18696 53780
rect 18651 53740 18696 53768
rect 18690 53728 18696 53740
rect 18748 53728 18754 53780
rect 19426 53768 19432 53780
rect 19387 53740 19432 53768
rect 19426 53728 19432 53740
rect 19484 53728 19490 53780
rect 29638 53728 29644 53780
rect 29696 53768 29702 53780
rect 30009 53771 30067 53777
rect 30009 53768 30021 53771
rect 29696 53740 30021 53768
rect 29696 53728 29702 53740
rect 30009 53737 30021 53740
rect 30055 53768 30067 53771
rect 31018 53768 31024 53780
rect 30055 53740 31024 53768
rect 30055 53737 30067 53740
rect 30009 53731 30067 53737
rect 31018 53728 31024 53740
rect 31076 53728 31082 53780
rect 22186 53660 22192 53712
rect 22244 53700 22250 53712
rect 22244 53672 29868 53700
rect 22244 53660 22250 53672
rect 19334 53592 19340 53644
rect 19392 53592 19398 53644
rect 19794 53592 19800 53644
rect 19852 53632 19858 53644
rect 23106 53632 23112 53644
rect 19852 53604 23112 53632
rect 19852 53592 19858 53604
rect 23106 53592 23112 53604
rect 23164 53592 23170 53644
rect 24394 53592 24400 53644
rect 24452 53632 24458 53644
rect 25866 53632 25872 53644
rect 24452 53604 25872 53632
rect 24452 53592 24458 53604
rect 25866 53592 25872 53604
rect 25924 53632 25930 53644
rect 25924 53604 26924 53632
rect 25924 53592 25930 53604
rect 1397 53567 1455 53573
rect 1397 53533 1409 53567
rect 1443 53564 1455 53567
rect 2222 53564 2228 53576
rect 1443 53536 2228 53564
rect 1443 53533 1455 53536
rect 1397 53527 1455 53533
rect 2222 53524 2228 53536
rect 2280 53524 2286 53576
rect 2317 53567 2375 53573
rect 2317 53533 2329 53567
rect 2363 53564 2375 53567
rect 6270 53564 6276 53576
rect 2363 53536 6276 53564
rect 2363 53533 2375 53536
rect 2317 53527 2375 53533
rect 6270 53524 6276 53536
rect 6328 53524 6334 53576
rect 17862 53564 17868 53576
rect 17823 53536 17868 53564
rect 17862 53524 17868 53536
rect 17920 53524 17926 53576
rect 18509 53567 18567 53573
rect 18509 53533 18521 53567
rect 18555 53564 18567 53567
rect 19352 53564 19380 53592
rect 19978 53564 19984 53576
rect 18555 53536 19380 53564
rect 19939 53536 19984 53564
rect 18555 53533 18567 53536
rect 18509 53527 18567 53533
rect 19978 53524 19984 53536
rect 20036 53524 20042 53576
rect 22370 53564 22376 53576
rect 22331 53536 22376 53564
rect 22370 53524 22376 53536
rect 22428 53524 22434 53576
rect 25777 53567 25835 53573
rect 25777 53533 25789 53567
rect 25823 53533 25835 53567
rect 25777 53527 25835 53533
rect 19337 53499 19395 53505
rect 19337 53465 19349 53499
rect 19383 53496 19395 53499
rect 21174 53496 21180 53508
rect 19383 53468 21180 53496
rect 19383 53465 19395 53468
rect 19337 53459 19395 53465
rect 21174 53456 21180 53468
rect 21232 53456 21238 53508
rect 22554 53456 22560 53508
rect 22612 53496 22618 53508
rect 23106 53496 23112 53508
rect 22612 53468 23112 53496
rect 22612 53456 22618 53468
rect 23106 53456 23112 53468
rect 23164 53456 23170 53508
rect 25792 53496 25820 53527
rect 26142 53524 26148 53576
rect 26200 53564 26206 53576
rect 26896 53573 26924 53604
rect 26697 53567 26755 53573
rect 26697 53564 26709 53567
rect 26200 53536 26709 53564
rect 26200 53524 26206 53536
rect 26697 53533 26709 53536
rect 26743 53533 26755 53567
rect 26697 53527 26755 53533
rect 26881 53567 26939 53573
rect 26881 53533 26893 53567
rect 26927 53533 26939 53567
rect 26881 53527 26939 53533
rect 26970 53524 26976 53576
rect 27028 53564 27034 53576
rect 27982 53564 27988 53576
rect 27028 53536 27073 53564
rect 27943 53536 27988 53564
rect 27028 53524 27034 53536
rect 27982 53524 27988 53536
rect 28040 53524 28046 53576
rect 28718 53564 28724 53576
rect 28679 53536 28724 53564
rect 28718 53524 28724 53536
rect 28776 53524 28782 53576
rect 29730 53564 29736 53576
rect 29691 53536 29736 53564
rect 29730 53524 29736 53536
rect 29788 53524 29794 53576
rect 25792 53468 26648 53496
rect 1578 53428 1584 53440
rect 1539 53400 1584 53428
rect 1578 53388 1584 53400
rect 1636 53388 1642 53440
rect 21266 53428 21272 53440
rect 21227 53400 21272 53428
rect 21266 53388 21272 53400
rect 21324 53388 21330 53440
rect 22462 53428 22468 53440
rect 22423 53400 22468 53428
rect 22462 53388 22468 53400
rect 22520 53388 22526 53440
rect 25958 53428 25964 53440
rect 25919 53400 25964 53428
rect 25958 53388 25964 53400
rect 26016 53388 26022 53440
rect 26510 53428 26516 53440
rect 26471 53400 26516 53428
rect 26510 53388 26516 53400
rect 26568 53388 26574 53440
rect 26620 53428 26648 53468
rect 27706 53428 27712 53440
rect 26620 53400 27712 53428
rect 27706 53388 27712 53400
rect 27764 53388 27770 53440
rect 28166 53428 28172 53440
rect 28127 53400 28172 53428
rect 28166 53388 28172 53400
rect 28224 53388 28230 53440
rect 28905 53431 28963 53437
rect 28905 53397 28917 53431
rect 28951 53428 28963 53431
rect 29086 53428 29092 53440
rect 28951 53400 29092 53428
rect 28951 53397 28963 53400
rect 28905 53391 28963 53397
rect 29086 53388 29092 53400
rect 29144 53388 29150 53440
rect 29730 53388 29736 53440
rect 29788 53428 29794 53440
rect 29840 53428 29868 53672
rect 29788 53400 29868 53428
rect 29788 53388 29794 53400
rect 1104 53338 30820 53360
rect 1104 53286 10880 53338
rect 10932 53286 10944 53338
rect 10996 53286 11008 53338
rect 11060 53286 11072 53338
rect 11124 53286 11136 53338
rect 11188 53286 20811 53338
rect 20863 53286 20875 53338
rect 20927 53286 20939 53338
rect 20991 53286 21003 53338
rect 21055 53286 21067 53338
rect 21119 53286 30820 53338
rect 1104 53264 30820 53286
rect 1394 53184 1400 53236
rect 1452 53224 1458 53236
rect 1673 53227 1731 53233
rect 1673 53224 1685 53227
rect 1452 53196 1685 53224
rect 1452 53184 1458 53196
rect 1673 53193 1685 53196
rect 1719 53193 1731 53227
rect 1673 53187 1731 53193
rect 2222 53184 2228 53236
rect 2280 53224 2286 53236
rect 17770 53224 17776 53236
rect 2280 53196 17264 53224
rect 17731 53196 17776 53224
rect 2280 53184 2286 53196
rect 1857 53091 1915 53097
rect 1857 53057 1869 53091
rect 1903 53088 1915 53091
rect 1946 53088 1952 53100
rect 1903 53060 1952 53088
rect 1903 53057 1915 53060
rect 1857 53051 1915 53057
rect 1946 53048 1952 53060
rect 2004 53048 2010 53100
rect 14182 53097 14188 53100
rect 14176 53051 14188 53097
rect 14240 53088 14246 53100
rect 14240 53060 14276 53088
rect 14182 53048 14188 53051
rect 14240 53048 14246 53060
rect 13906 53020 13912 53032
rect 13867 52992 13912 53020
rect 13906 52980 13912 52992
rect 13964 52980 13970 53032
rect 17236 53020 17264 53196
rect 17770 53184 17776 53196
rect 17828 53184 17834 53236
rect 18509 53227 18567 53233
rect 18509 53193 18521 53227
rect 18555 53224 18567 53227
rect 19242 53224 19248 53236
rect 18555 53196 19248 53224
rect 18555 53193 18567 53196
rect 18509 53187 18567 53193
rect 19242 53184 19248 53196
rect 19300 53184 19306 53236
rect 19702 53184 19708 53236
rect 19760 53224 19766 53236
rect 19889 53227 19947 53233
rect 19889 53224 19901 53227
rect 19760 53196 19901 53224
rect 19760 53184 19766 53196
rect 19889 53193 19901 53196
rect 19935 53193 19947 53227
rect 19889 53187 19947 53193
rect 21269 53227 21327 53233
rect 21269 53193 21281 53227
rect 21315 53224 21327 53227
rect 22094 53224 22100 53236
rect 21315 53196 22100 53224
rect 21315 53193 21327 53196
rect 21269 53187 21327 53193
rect 22094 53184 22100 53196
rect 22152 53184 22158 53236
rect 27433 53227 27491 53233
rect 27433 53193 27445 53227
rect 27479 53224 27491 53227
rect 27890 53224 27896 53236
rect 27479 53196 27896 53224
rect 27479 53193 27491 53196
rect 27433 53187 27491 53193
rect 27890 53184 27896 53196
rect 27948 53184 27954 53236
rect 28166 53184 28172 53236
rect 28224 53224 28230 53236
rect 29270 53224 29276 53236
rect 28224 53196 28856 53224
rect 29231 53196 29276 53224
rect 28224 53184 28230 53196
rect 17681 53159 17739 53165
rect 17681 53125 17693 53159
rect 17727 53156 17739 53159
rect 18230 53156 18236 53168
rect 17727 53128 18236 53156
rect 17727 53125 17739 53128
rect 17681 53119 17739 53125
rect 18230 53116 18236 53128
rect 18288 53116 18294 53168
rect 19061 53159 19119 53165
rect 19061 53125 19073 53159
rect 19107 53156 19119 53159
rect 20162 53156 20168 53168
rect 19107 53128 20168 53156
rect 19107 53125 19119 53128
rect 19061 53119 19119 53125
rect 20162 53116 20168 53128
rect 20220 53116 20226 53168
rect 20714 53116 20720 53168
rect 20772 53156 20778 53168
rect 21913 53159 21971 53165
rect 21913 53156 21925 53159
rect 20772 53128 21925 53156
rect 20772 53116 20778 53128
rect 21913 53125 21925 53128
rect 21959 53125 21971 53159
rect 21913 53119 21971 53125
rect 25314 53116 25320 53168
rect 25372 53156 25378 53168
rect 26329 53159 26387 53165
rect 26329 53156 26341 53159
rect 25372 53128 26341 53156
rect 25372 53116 25378 53128
rect 26329 53125 26341 53128
rect 26375 53125 26387 53159
rect 26329 53119 26387 53125
rect 26510 53116 26516 53168
rect 26568 53156 26574 53168
rect 26568 53128 28120 53156
rect 26568 53116 26574 53128
rect 18322 53088 18328 53100
rect 18283 53060 18328 53088
rect 18322 53048 18328 53060
rect 18380 53048 18386 53100
rect 19150 53048 19156 53100
rect 19208 53088 19214 53100
rect 19705 53091 19763 53097
rect 19705 53088 19717 53091
rect 19208 53060 19717 53088
rect 19208 53048 19214 53060
rect 19705 53057 19717 53060
rect 19751 53057 19763 53091
rect 19705 53051 19763 53057
rect 21085 53091 21143 53097
rect 21085 53057 21097 53091
rect 21131 53088 21143 53091
rect 21818 53088 21824 53100
rect 21131 53060 21824 53088
rect 21131 53057 21143 53060
rect 21085 53051 21143 53057
rect 21818 53048 21824 53060
rect 21876 53048 21882 53100
rect 22094 53048 22100 53100
rect 22152 53088 22158 53100
rect 22370 53088 22376 53100
rect 22152 53060 22376 53088
rect 22152 53048 22158 53060
rect 22370 53048 22376 53060
rect 22428 53088 22434 53100
rect 22557 53091 22615 53097
rect 22557 53088 22569 53091
rect 22428 53060 22569 53088
rect 22428 53048 22434 53060
rect 22557 53057 22569 53060
rect 22603 53057 22615 53091
rect 22557 53051 22615 53057
rect 23569 53091 23627 53097
rect 23569 53057 23581 53091
rect 23615 53088 23627 53091
rect 23658 53088 23664 53100
rect 23615 53060 23664 53088
rect 23615 53057 23627 53060
rect 23569 53051 23627 53057
rect 23658 53048 23664 53060
rect 23716 53048 23722 53100
rect 26142 53088 26148 53100
rect 26103 53060 26148 53088
rect 26142 53048 26148 53060
rect 26200 53048 26206 53100
rect 26421 53091 26479 53097
rect 26421 53057 26433 53091
rect 26467 53057 26479 53091
rect 26421 53051 26479 53057
rect 23290 53020 23296 53032
rect 17236 52992 23296 53020
rect 23290 52980 23296 52992
rect 23348 52980 23354 53032
rect 26436 53020 26464 53051
rect 27338 53048 27344 53100
rect 27396 53088 27402 53100
rect 27614 53088 27620 53100
rect 27396 53060 27620 53088
rect 27396 53048 27402 53060
rect 27614 53048 27620 53060
rect 27672 53088 27678 53100
rect 27709 53091 27767 53097
rect 27709 53088 27721 53091
rect 27672 53060 27721 53088
rect 27672 53048 27678 53060
rect 27709 53057 27721 53060
rect 27755 53057 27767 53091
rect 27709 53051 27767 53057
rect 27801 53091 27859 53097
rect 27801 53057 27813 53091
rect 27847 53057 27859 53091
rect 27801 53051 27859 53057
rect 26970 53020 26976 53032
rect 23676 52992 26976 53020
rect 19242 52952 19248 52964
rect 19203 52924 19248 52952
rect 19242 52912 19248 52924
rect 19300 52912 19306 52964
rect 21910 52912 21916 52964
rect 21968 52952 21974 52964
rect 22649 52955 22707 52961
rect 22649 52952 22661 52955
rect 21968 52924 22661 52952
rect 21968 52912 21974 52924
rect 22649 52921 22661 52924
rect 22695 52921 22707 52955
rect 22649 52915 22707 52921
rect 23676 52896 23704 52992
rect 26970 52980 26976 52992
rect 27028 52980 27034 53032
rect 25866 52912 25872 52964
rect 25924 52912 25930 52964
rect 25961 52955 26019 52961
rect 25961 52921 25973 52955
rect 26007 52952 26019 52955
rect 27706 52952 27712 52964
rect 26007 52924 27712 52952
rect 26007 52921 26019 52924
rect 25961 52915 26019 52921
rect 27706 52912 27712 52924
rect 27764 52912 27770 52964
rect 27816 52952 27844 53051
rect 27890 53048 27896 53100
rect 27948 53088 27954 53100
rect 28092 53097 28120 53128
rect 28442 53116 28448 53168
rect 28500 53156 28506 53168
rect 28500 53128 28764 53156
rect 28500 53116 28506 53128
rect 28077 53091 28135 53097
rect 27948 53060 27993 53088
rect 27948 53048 27954 53060
rect 28077 53057 28089 53091
rect 28123 53057 28135 53091
rect 28077 53051 28135 53057
rect 28537 53091 28595 53097
rect 28537 53057 28549 53091
rect 28583 53088 28595 53091
rect 28626 53088 28632 53100
rect 28583 53060 28632 53088
rect 28583 53057 28595 53060
rect 28537 53051 28595 53057
rect 28626 53048 28632 53060
rect 28684 53048 28690 53100
rect 28736 53097 28764 53128
rect 28721 53091 28779 53097
rect 28721 53057 28733 53091
rect 28767 53057 28779 53091
rect 28828 53088 28856 53196
rect 29270 53184 29276 53196
rect 29328 53184 29334 53236
rect 28905 53091 28963 53097
rect 28905 53088 28917 53091
rect 28828 53060 28917 53088
rect 28721 53051 28779 53057
rect 28905 53057 28917 53060
rect 28951 53057 28963 53091
rect 28905 53051 28963 53057
rect 29089 53091 29147 53097
rect 29089 53057 29101 53091
rect 29135 53088 29147 53091
rect 29638 53088 29644 53100
rect 29135 53060 29644 53088
rect 29135 53057 29147 53060
rect 29089 53051 29147 53057
rect 29638 53048 29644 53060
rect 29696 53048 29702 53100
rect 29825 53091 29883 53097
rect 29825 53057 29837 53091
rect 29871 53088 29883 53091
rect 30006 53088 30012 53100
rect 29871 53060 30012 53088
rect 29871 53057 29883 53060
rect 29825 53051 29883 53057
rect 30006 53048 30012 53060
rect 30064 53048 30070 53100
rect 28813 53023 28871 53029
rect 28813 52989 28825 53023
rect 28859 53020 28871 53023
rect 29730 53020 29736 53032
rect 28859 52992 29736 53020
rect 28859 52989 28871 52992
rect 28813 52983 28871 52989
rect 29730 52980 29736 52992
rect 29788 53020 29794 53032
rect 30926 53020 30932 53032
rect 29788 52992 30932 53020
rect 29788 52980 29794 52992
rect 30926 52980 30932 52992
rect 30984 52980 30990 53032
rect 29270 52952 29276 52964
rect 27816 52924 29276 52952
rect 29270 52912 29276 52924
rect 29328 52912 29334 52964
rect 14274 52844 14280 52896
rect 14332 52884 14338 52896
rect 15289 52887 15347 52893
rect 15289 52884 15301 52887
rect 14332 52856 15301 52884
rect 14332 52844 14338 52856
rect 15289 52853 15301 52856
rect 15335 52884 15347 52887
rect 19794 52884 19800 52896
rect 15335 52856 19800 52884
rect 15335 52853 15347 52856
rect 15289 52847 15347 52853
rect 19794 52844 19800 52856
rect 19852 52844 19858 52896
rect 20622 52844 20628 52896
rect 20680 52884 20686 52896
rect 22005 52887 22063 52893
rect 22005 52884 22017 52887
rect 20680 52856 22017 52884
rect 20680 52844 20686 52856
rect 22005 52853 22017 52856
rect 22051 52853 22063 52887
rect 23658 52884 23664 52896
rect 23619 52856 23664 52884
rect 22005 52847 22063 52853
rect 23658 52844 23664 52856
rect 23716 52844 23722 52896
rect 25884 52884 25912 52912
rect 26326 52884 26332 52896
rect 25884 52856 26332 52884
rect 26326 52844 26332 52856
rect 26384 52844 26390 52896
rect 28626 52844 28632 52896
rect 28684 52884 28690 52896
rect 29822 52884 29828 52896
rect 28684 52856 29828 52884
rect 28684 52844 28690 52856
rect 29822 52844 29828 52856
rect 29880 52844 29886 52896
rect 30009 52887 30067 52893
rect 30009 52853 30021 52887
rect 30055 52884 30067 52887
rect 31662 52884 31668 52896
rect 30055 52856 31668 52884
rect 30055 52853 30067 52856
rect 30009 52847 30067 52853
rect 31662 52844 31668 52856
rect 31720 52844 31726 52896
rect 1104 52794 30820 52816
rect 1104 52742 5915 52794
rect 5967 52742 5979 52794
rect 6031 52742 6043 52794
rect 6095 52742 6107 52794
rect 6159 52742 6171 52794
rect 6223 52742 15846 52794
rect 15898 52742 15910 52794
rect 15962 52742 15974 52794
rect 16026 52742 16038 52794
rect 16090 52742 16102 52794
rect 16154 52742 25776 52794
rect 25828 52742 25840 52794
rect 25892 52742 25904 52794
rect 25956 52742 25968 52794
rect 26020 52742 26032 52794
rect 26084 52742 30820 52794
rect 1104 52720 30820 52742
rect 13354 52680 13360 52692
rect 13315 52652 13360 52680
rect 13354 52640 13360 52652
rect 13412 52680 13418 52692
rect 13538 52680 13544 52692
rect 13412 52652 13544 52680
rect 13412 52640 13418 52652
rect 13538 52640 13544 52652
rect 13596 52640 13602 52692
rect 13906 52640 13912 52692
rect 13964 52680 13970 52692
rect 15381 52683 15439 52689
rect 15381 52680 15393 52683
rect 13964 52652 15393 52680
rect 13964 52640 13970 52652
rect 15381 52649 15393 52652
rect 15427 52649 15439 52683
rect 15381 52643 15439 52649
rect 17681 52683 17739 52689
rect 17681 52649 17693 52683
rect 17727 52680 17739 52683
rect 17862 52680 17868 52692
rect 17727 52652 17868 52680
rect 17727 52649 17739 52652
rect 17681 52643 17739 52649
rect 17862 52640 17868 52652
rect 17920 52640 17926 52692
rect 18322 52640 18328 52692
rect 18380 52680 18386 52692
rect 19337 52683 19395 52689
rect 19337 52680 19349 52683
rect 18380 52652 19349 52680
rect 18380 52640 18386 52652
rect 19337 52649 19349 52652
rect 19383 52649 19395 52683
rect 19337 52643 19395 52649
rect 20530 52640 20536 52692
rect 20588 52680 20594 52692
rect 20717 52683 20775 52689
rect 20717 52680 20729 52683
rect 20588 52652 20729 52680
rect 20588 52640 20594 52652
rect 20717 52649 20729 52652
rect 20763 52649 20775 52683
rect 23290 52680 23296 52692
rect 23251 52652 23296 52680
rect 20717 52643 20775 52649
rect 23290 52640 23296 52652
rect 23348 52640 23354 52692
rect 26602 52640 26608 52692
rect 26660 52680 26666 52692
rect 27157 52683 27215 52689
rect 27157 52680 27169 52683
rect 26660 52652 27169 52680
rect 26660 52640 26666 52652
rect 27157 52649 27169 52652
rect 27203 52649 27215 52683
rect 29178 52680 29184 52692
rect 27157 52643 27215 52649
rect 27448 52652 27752 52680
rect 1397 52615 1455 52621
rect 1397 52581 1409 52615
rect 1443 52612 1455 52615
rect 1486 52612 1492 52624
rect 1443 52584 1492 52612
rect 1443 52581 1455 52584
rect 1397 52575 1455 52581
rect 1486 52572 1492 52584
rect 1544 52572 1550 52624
rect 2038 52612 2044 52624
rect 1999 52584 2044 52612
rect 2038 52572 2044 52584
rect 2096 52572 2102 52624
rect 14093 52615 14151 52621
rect 14093 52581 14105 52615
rect 14139 52612 14151 52615
rect 14182 52612 14188 52624
rect 14139 52584 14188 52612
rect 14139 52581 14151 52584
rect 14093 52575 14151 52581
rect 14182 52572 14188 52584
rect 14240 52572 14246 52624
rect 18506 52572 18512 52624
rect 18564 52612 18570 52624
rect 21726 52612 21732 52624
rect 18564 52584 21732 52612
rect 18564 52572 18570 52584
rect 21726 52572 21732 52584
rect 21784 52572 21790 52624
rect 27448 52612 27476 52652
rect 26252 52584 27476 52612
rect 2866 52504 2872 52556
rect 2924 52544 2930 52556
rect 19797 52547 19855 52553
rect 2924 52516 14780 52544
rect 2924 52504 2930 52516
rect 1578 52476 1584 52488
rect 1539 52448 1584 52476
rect 1578 52436 1584 52448
rect 1636 52436 1642 52488
rect 2222 52476 2228 52488
rect 2183 52448 2228 52476
rect 2222 52436 2228 52448
rect 2280 52436 2286 52488
rect 11790 52476 11796 52488
rect 11751 52448 11796 52476
rect 11790 52436 11796 52448
rect 11848 52436 11854 52488
rect 11882 52436 11888 52488
rect 11940 52476 11946 52488
rect 12069 52479 12127 52485
rect 12069 52476 12081 52479
rect 11940 52448 12081 52476
rect 11940 52436 11946 52448
rect 12069 52445 12081 52448
rect 12115 52445 12127 52479
rect 12069 52439 12127 52445
rect 14274 52436 14280 52488
rect 14332 52476 14338 52488
rect 14752 52485 14780 52516
rect 19797 52513 19809 52547
rect 19843 52544 19855 52547
rect 20622 52544 20628 52556
rect 19843 52516 20628 52544
rect 19843 52513 19855 52516
rect 19797 52507 19855 52513
rect 20622 52504 20628 52516
rect 20680 52504 20686 52556
rect 21910 52544 21916 52556
rect 21871 52516 21916 52544
rect 21910 52504 21916 52516
rect 21968 52504 21974 52556
rect 23750 52504 23756 52556
rect 23808 52544 23814 52556
rect 24302 52544 24308 52556
rect 23808 52516 24308 52544
rect 23808 52504 23814 52516
rect 24302 52504 24308 52516
rect 24360 52504 24366 52556
rect 26252 52553 26280 52584
rect 27522 52572 27528 52624
rect 27580 52612 27586 52624
rect 27580 52584 27665 52612
rect 27580 52572 27586 52584
rect 26237 52547 26295 52553
rect 26237 52513 26249 52547
rect 26283 52513 26295 52547
rect 26237 52507 26295 52513
rect 14369 52479 14427 52485
rect 14369 52476 14381 52479
rect 14332 52448 14381 52476
rect 14332 52436 14338 52448
rect 14369 52445 14381 52448
rect 14415 52445 14427 52479
rect 14369 52439 14427 52445
rect 14461 52479 14519 52485
rect 14461 52445 14473 52479
rect 14507 52445 14519 52479
rect 14461 52439 14519 52445
rect 14553 52479 14611 52485
rect 14553 52445 14565 52479
rect 14599 52445 14611 52479
rect 14553 52439 14611 52445
rect 14737 52479 14795 52485
rect 14737 52445 14749 52479
rect 14783 52445 14795 52479
rect 14737 52439 14795 52445
rect 14476 52408 14504 52439
rect 14384 52380 14504 52408
rect 14568 52408 14596 52439
rect 14826 52436 14832 52488
rect 14884 52476 14890 52488
rect 15197 52479 15255 52485
rect 15197 52476 15209 52479
rect 14884 52448 15209 52476
rect 14884 52436 14890 52448
rect 15197 52445 15209 52448
rect 15243 52445 15255 52479
rect 15197 52439 15255 52445
rect 17129 52479 17187 52485
rect 17129 52445 17141 52479
rect 17175 52476 17187 52479
rect 17957 52479 18015 52485
rect 17957 52476 17969 52479
rect 17175 52448 17969 52476
rect 17175 52445 17187 52448
rect 17129 52439 17187 52445
rect 17957 52445 17969 52448
rect 18003 52476 18015 52479
rect 18046 52476 18052 52488
rect 18003 52448 18052 52476
rect 18003 52445 18015 52448
rect 17957 52439 18015 52445
rect 18046 52436 18052 52448
rect 18104 52436 18110 52488
rect 18233 52479 18291 52485
rect 18233 52445 18245 52479
rect 18279 52476 18291 52479
rect 18322 52476 18328 52488
rect 18279 52448 18328 52476
rect 18279 52445 18291 52448
rect 18233 52439 18291 52445
rect 18322 52436 18328 52448
rect 18380 52436 18386 52488
rect 20714 52476 20720 52488
rect 19720 52448 20024 52476
rect 14918 52408 14924 52420
rect 14568 52380 14924 52408
rect 14384 52352 14412 52380
rect 14918 52368 14924 52380
rect 14976 52368 14982 52420
rect 16945 52411 17003 52417
rect 16945 52377 16957 52411
rect 16991 52377 17003 52411
rect 16945 52371 17003 52377
rect 14366 52300 14372 52352
rect 14424 52300 14430 52352
rect 16960 52340 16988 52371
rect 17770 52368 17776 52420
rect 17828 52408 17834 52420
rect 18141 52411 18199 52417
rect 18141 52408 18153 52411
rect 17828 52380 18153 52408
rect 17828 52368 17834 52380
rect 18141 52377 18153 52380
rect 18187 52377 18199 52411
rect 19720 52408 19748 52448
rect 19886 52408 19892 52420
rect 18141 52371 18199 52377
rect 18248 52380 19748 52408
rect 19847 52380 19892 52408
rect 18248 52340 18276 52380
rect 19886 52368 19892 52380
rect 19944 52368 19950 52420
rect 19996 52408 20024 52448
rect 20548 52448 20720 52476
rect 20548 52408 20576 52448
rect 20714 52436 20720 52448
rect 20772 52436 20778 52488
rect 26142 52436 26148 52488
rect 26200 52476 26206 52488
rect 26421 52479 26479 52485
rect 26421 52476 26433 52479
rect 26200 52448 26433 52476
rect 26200 52436 26206 52448
rect 26421 52445 26433 52448
rect 26467 52445 26479 52479
rect 26421 52439 26479 52445
rect 26697 52479 26755 52485
rect 26697 52445 26709 52479
rect 26743 52476 26755 52479
rect 26970 52476 26976 52488
rect 26743 52448 26976 52476
rect 26743 52445 26755 52448
rect 26697 52439 26755 52445
rect 26970 52436 26976 52448
rect 27028 52436 27034 52488
rect 27338 52436 27344 52488
rect 27396 52476 27402 52488
rect 27637 52485 27665 52584
rect 27433 52479 27491 52485
rect 27433 52476 27445 52479
rect 27396 52448 27445 52476
rect 27396 52436 27402 52448
rect 27433 52445 27445 52448
rect 27479 52445 27491 52479
rect 27433 52439 27491 52445
rect 27525 52476 27583 52482
rect 27525 52442 27537 52476
rect 27571 52442 27583 52476
rect 27525 52436 27583 52442
rect 27617 52479 27675 52485
rect 27617 52445 27629 52479
rect 27663 52445 27675 52479
rect 27724 52476 27752 52652
rect 27908 52652 29184 52680
rect 27801 52479 27859 52485
rect 27801 52476 27813 52479
rect 27724 52448 27813 52476
rect 27617 52439 27675 52445
rect 27801 52445 27813 52448
rect 27847 52445 27859 52479
rect 27908 52476 27936 52652
rect 29178 52640 29184 52652
rect 29236 52640 29242 52692
rect 29454 52640 29460 52692
rect 29512 52680 29518 52692
rect 29825 52683 29883 52689
rect 29825 52680 29837 52683
rect 29512 52652 29837 52680
rect 29512 52640 29518 52652
rect 29825 52649 29837 52652
rect 29871 52680 29883 52683
rect 30006 52680 30012 52692
rect 29871 52652 30012 52680
rect 29871 52649 29883 52652
rect 29825 52643 29883 52649
rect 30006 52640 30012 52652
rect 30064 52640 30070 52692
rect 28626 52612 28632 52624
rect 28552 52584 28632 52612
rect 27982 52504 27988 52556
rect 28040 52544 28046 52556
rect 28552 52553 28580 52584
rect 28626 52572 28632 52584
rect 28684 52612 28690 52624
rect 30834 52612 30840 52624
rect 28684 52584 30840 52612
rect 28684 52572 28690 52584
rect 30834 52572 30840 52584
rect 30892 52572 30898 52624
rect 28537 52547 28595 52553
rect 28040 52516 28304 52544
rect 28040 52504 28046 52516
rect 28276 52485 28304 52516
rect 28537 52513 28549 52547
rect 28583 52513 28595 52547
rect 28902 52544 28908 52556
rect 28537 52507 28595 52513
rect 28828 52516 28908 52544
rect 28261 52479 28319 52485
rect 27908 52448 28120 52476
rect 27801 52439 27859 52445
rect 22186 52417 22192 52420
rect 19996 52380 20576 52408
rect 20625 52411 20683 52417
rect 20625 52377 20637 52411
rect 20671 52377 20683 52411
rect 20625 52371 20683 52377
rect 22180 52371 22192 52417
rect 22244 52408 22250 52420
rect 22244 52380 22280 52408
rect 19794 52340 19800 52352
rect 16960 52312 18276 52340
rect 19755 52312 19800 52340
rect 19794 52300 19800 52312
rect 19852 52300 19858 52352
rect 20438 52300 20444 52352
rect 20496 52340 20502 52352
rect 20640 52340 20668 52371
rect 22186 52368 22192 52371
rect 22244 52368 22250 52380
rect 23934 52368 23940 52420
rect 23992 52408 23998 52420
rect 24302 52408 24308 52420
rect 23992 52380 24308 52408
rect 23992 52368 23998 52380
rect 24302 52368 24308 52380
rect 24360 52368 24366 52420
rect 26605 52411 26663 52417
rect 26605 52408 26617 52411
rect 25976 52380 26617 52408
rect 25976 52352 26004 52380
rect 26605 52377 26617 52380
rect 26651 52377 26663 52411
rect 27540 52408 27568 52436
rect 27982 52408 27988 52420
rect 27540 52380 27988 52408
rect 26605 52371 26663 52377
rect 27982 52368 27988 52380
rect 28040 52368 28046 52420
rect 20496 52312 20668 52340
rect 20496 52300 20502 52312
rect 23014 52300 23020 52352
rect 23072 52340 23078 52352
rect 25958 52340 25964 52352
rect 23072 52312 25964 52340
rect 23072 52300 23078 52312
rect 25958 52300 25964 52312
rect 26016 52300 26022 52352
rect 26694 52300 26700 52352
rect 26752 52340 26758 52352
rect 26878 52340 26884 52352
rect 26752 52312 26884 52340
rect 26752 52300 26758 52312
rect 26878 52300 26884 52312
rect 26936 52300 26942 52352
rect 27430 52300 27436 52352
rect 27488 52340 27494 52352
rect 28092 52340 28120 52448
rect 28261 52445 28273 52479
rect 28307 52445 28319 52479
rect 28442 52476 28448 52488
rect 28403 52448 28448 52476
rect 28261 52439 28319 52445
rect 28442 52436 28448 52448
rect 28500 52436 28506 52488
rect 28626 52476 28632 52488
rect 28587 52448 28632 52476
rect 28626 52436 28632 52448
rect 28684 52436 28690 52488
rect 28828 52485 28856 52516
rect 28902 52504 28908 52516
rect 28960 52504 28966 52556
rect 28994 52504 29000 52556
rect 29052 52544 29058 52556
rect 29270 52544 29276 52556
rect 29052 52516 29276 52544
rect 29052 52504 29058 52516
rect 29270 52504 29276 52516
rect 29328 52504 29334 52556
rect 28813 52479 28871 52485
rect 28813 52445 28825 52479
rect 28859 52445 28871 52479
rect 28813 52439 28871 52445
rect 29730 52408 29736 52420
rect 29691 52380 29736 52408
rect 29730 52368 29736 52380
rect 29788 52368 29794 52420
rect 28994 52340 29000 52352
rect 27488 52312 28120 52340
rect 28955 52312 29000 52340
rect 27488 52300 27494 52312
rect 28994 52300 29000 52312
rect 29052 52300 29058 52352
rect 29546 52300 29552 52352
rect 29604 52340 29610 52352
rect 29604 52312 30880 52340
rect 29604 52300 29610 52312
rect 1104 52250 30820 52272
rect 1104 52198 10880 52250
rect 10932 52198 10944 52250
rect 10996 52198 11008 52250
rect 11060 52198 11072 52250
rect 11124 52198 11136 52250
rect 11188 52198 20811 52250
rect 20863 52198 20875 52250
rect 20927 52198 20939 52250
rect 20991 52198 21003 52250
rect 21055 52198 21067 52250
rect 21119 52198 30820 52250
rect 1104 52176 30820 52198
rect 1857 52139 1915 52145
rect 1857 52105 1869 52139
rect 1903 52136 1915 52139
rect 2222 52136 2228 52148
rect 1903 52108 2228 52136
rect 1903 52105 1915 52108
rect 1857 52099 1915 52105
rect 2222 52096 2228 52108
rect 2280 52096 2286 52148
rect 11701 52139 11759 52145
rect 11701 52105 11713 52139
rect 11747 52136 11759 52139
rect 11790 52136 11796 52148
rect 11747 52108 11796 52136
rect 11747 52105 11759 52108
rect 11701 52099 11759 52105
rect 11790 52096 11796 52108
rect 11848 52096 11854 52148
rect 11900 52108 16896 52136
rect 11900 52068 11928 52108
rect 6886 52040 11928 52068
rect 1673 52003 1731 52009
rect 1673 51969 1685 52003
rect 1719 52000 1731 52003
rect 6886 52000 6914 52040
rect 13998 52028 14004 52080
rect 14056 52068 14062 52080
rect 14277 52071 14335 52077
rect 14277 52068 14289 52071
rect 14056 52040 14289 52068
rect 14056 52028 14062 52040
rect 14277 52037 14289 52040
rect 14323 52068 14335 52071
rect 14642 52068 14648 52080
rect 14323 52040 14648 52068
rect 14323 52037 14335 52040
rect 14277 52031 14335 52037
rect 14642 52028 14648 52040
rect 14700 52028 14706 52080
rect 16868 52068 16896 52108
rect 16942 52096 16948 52148
rect 17000 52136 17006 52148
rect 17221 52139 17279 52145
rect 17221 52136 17233 52139
rect 17000 52108 17233 52136
rect 17000 52096 17006 52108
rect 17221 52105 17233 52108
rect 17267 52105 17279 52139
rect 18233 52139 18291 52145
rect 17221 52099 17279 52105
rect 17328 52108 18184 52136
rect 17328 52068 17356 52108
rect 18046 52068 18052 52080
rect 16868 52040 17356 52068
rect 18007 52040 18052 52068
rect 18046 52028 18052 52040
rect 18104 52028 18110 52080
rect 18156 52068 18184 52108
rect 18233 52105 18245 52139
rect 18279 52136 18291 52139
rect 19794 52136 19800 52148
rect 18279 52108 19800 52136
rect 18279 52105 18291 52108
rect 18233 52099 18291 52105
rect 19794 52096 19800 52108
rect 19852 52096 19858 52148
rect 22373 52139 22431 52145
rect 22373 52105 22385 52139
rect 22419 52136 22431 52139
rect 22462 52136 22468 52148
rect 22419 52108 22468 52136
rect 22419 52105 22431 52108
rect 22373 52099 22431 52105
rect 22462 52096 22468 52108
rect 22520 52096 22526 52148
rect 23014 52096 23020 52148
rect 23072 52136 23078 52148
rect 23566 52136 23572 52148
rect 23072 52108 23572 52136
rect 23072 52096 23078 52108
rect 23566 52096 23572 52108
rect 23624 52096 23630 52148
rect 24394 52096 24400 52148
rect 24452 52136 24458 52148
rect 25869 52139 25927 52145
rect 25869 52136 25881 52139
rect 24452 52108 25881 52136
rect 24452 52096 24458 52108
rect 25869 52105 25881 52108
rect 25915 52105 25927 52139
rect 25869 52099 25927 52105
rect 25958 52096 25964 52148
rect 26016 52136 26022 52148
rect 27065 52139 27123 52145
rect 26016 52108 26061 52136
rect 26016 52096 26022 52108
rect 27065 52105 27077 52139
rect 27111 52136 27123 52139
rect 27430 52136 27436 52148
rect 27111 52108 27436 52136
rect 27111 52105 27123 52108
rect 27065 52099 27123 52105
rect 27430 52096 27436 52108
rect 27488 52096 27494 52148
rect 28718 52096 28724 52148
rect 28776 52136 28782 52148
rect 29362 52136 29368 52148
rect 28776 52108 29368 52136
rect 28776 52096 28782 52108
rect 29362 52096 29368 52108
rect 29420 52096 29426 52148
rect 30101 52139 30159 52145
rect 30101 52105 30113 52139
rect 30147 52136 30159 52139
rect 30852 52136 30880 52312
rect 30147 52108 30880 52136
rect 30147 52105 30159 52108
rect 30101 52099 30159 52105
rect 21895 52071 21953 52077
rect 21895 52068 21907 52071
rect 18156 52040 21907 52068
rect 21895 52037 21907 52040
rect 21941 52037 21953 52071
rect 21895 52031 21953 52037
rect 25682 52028 25688 52080
rect 25740 52068 25746 52080
rect 26145 52071 26203 52077
rect 26145 52068 26157 52071
rect 25740 52040 26157 52068
rect 25740 52028 25746 52040
rect 26145 52037 26157 52040
rect 26191 52037 26203 52071
rect 26145 52031 26203 52037
rect 26602 52028 26608 52080
rect 26660 52068 26666 52080
rect 26660 52040 27476 52068
rect 26660 52028 26666 52040
rect 1719 51972 6914 52000
rect 11517 52003 11575 52009
rect 1719 51969 1731 51972
rect 1673 51963 1731 51969
rect 11517 51969 11529 52003
rect 11563 52000 11575 52003
rect 11606 52000 11612 52012
rect 11563 51972 11612 52000
rect 11563 51969 11575 51972
rect 11517 51963 11575 51969
rect 11606 51960 11612 51972
rect 11664 51960 11670 52012
rect 14458 51960 14464 52012
rect 14516 52000 14522 52012
rect 14993 52003 15051 52009
rect 14993 52000 15005 52003
rect 14516 51972 15005 52000
rect 14516 51960 14522 51972
rect 14993 51969 15005 51972
rect 15039 51969 15051 52003
rect 17034 52000 17040 52012
rect 16995 51972 17040 52000
rect 14993 51963 15051 51969
rect 17034 51960 17040 51972
rect 17092 51960 17098 52012
rect 17954 51960 17960 52012
rect 18012 52000 18018 52012
rect 18877 52003 18935 52009
rect 18877 52000 18889 52003
rect 18012 51972 18889 52000
rect 18012 51960 18018 51972
rect 18877 51969 18889 51972
rect 18923 51969 18935 52003
rect 18877 51963 18935 51969
rect 20625 52003 20683 52009
rect 20625 51969 20637 52003
rect 20671 52000 20683 52003
rect 20714 52000 20720 52012
rect 20671 51972 20720 52000
rect 20671 51969 20683 51972
rect 20625 51963 20683 51969
rect 20714 51960 20720 51972
rect 20772 51960 20778 52012
rect 22922 51960 22928 52012
rect 22980 52000 22986 52012
rect 23293 52003 23351 52009
rect 23293 52000 23305 52003
rect 22980 51972 23305 52000
rect 22980 51960 22986 51972
rect 23293 51969 23305 51972
rect 23339 51969 23351 52003
rect 23293 51963 23351 51969
rect 25590 51960 25596 52012
rect 25648 52000 25654 52012
rect 25777 52003 25835 52009
rect 25777 52000 25789 52003
rect 25648 51972 25789 52000
rect 25648 51960 25654 51972
rect 25777 51969 25789 51972
rect 25823 51969 25835 52003
rect 27338 52000 27344 52012
rect 27299 51972 27344 52000
rect 25777 51963 25835 51969
rect 27338 51960 27344 51972
rect 27396 51960 27402 52012
rect 27448 52009 27476 52040
rect 28442 52028 28448 52080
rect 28500 52068 28506 52080
rect 28500 52040 29592 52068
rect 28500 52028 28506 52040
rect 27433 52003 27491 52009
rect 27433 51969 27445 52003
rect 27479 51969 27491 52003
rect 27433 51963 27491 51969
rect 27525 52003 27583 52009
rect 27525 51969 27537 52003
rect 27571 51969 27583 52003
rect 27706 52000 27712 52012
rect 27667 51972 27712 52000
rect 27525 51963 27583 51969
rect 12618 51932 12624 51944
rect 12579 51904 12624 51932
rect 12618 51892 12624 51904
rect 12676 51892 12682 51944
rect 12894 51932 12900 51944
rect 12855 51904 12900 51932
rect 12894 51892 12900 51904
rect 12952 51892 12958 51944
rect 14734 51932 14740 51944
rect 14695 51904 14740 51932
rect 14734 51892 14740 51904
rect 14792 51892 14798 51944
rect 18322 51932 18328 51944
rect 18283 51904 18328 51932
rect 18322 51892 18328 51904
rect 18380 51892 18386 51944
rect 21726 51892 21732 51944
rect 21784 51932 21790 51944
rect 22281 51935 22339 51941
rect 22281 51932 22293 51935
rect 21784 51904 22293 51932
rect 21784 51892 21790 51904
rect 22281 51901 22293 51904
rect 22327 51901 22339 51935
rect 22281 51895 22339 51901
rect 22465 51935 22523 51941
rect 22465 51901 22477 51935
rect 22511 51932 22523 51935
rect 22554 51932 22560 51944
rect 22511 51904 22560 51932
rect 22511 51901 22523 51904
rect 22465 51895 22523 51901
rect 22554 51892 22560 51904
rect 22612 51892 22618 51944
rect 23569 51935 23627 51941
rect 23569 51901 23581 51935
rect 23615 51932 23627 51935
rect 24394 51932 24400 51944
rect 23615 51904 24400 51932
rect 23615 51901 23627 51904
rect 23569 51895 23627 51901
rect 24394 51892 24400 51904
rect 24452 51892 24458 51944
rect 26602 51892 26608 51944
rect 26660 51932 26666 51944
rect 27540 51932 27568 51963
rect 27706 51960 27712 51972
rect 27764 51960 27770 52012
rect 28169 52003 28227 52009
rect 28169 52000 28181 52003
rect 27908 51972 28181 52000
rect 26660 51904 27568 51932
rect 26660 51892 26666 51904
rect 17773 51867 17831 51873
rect 17773 51833 17785 51867
rect 17819 51864 17831 51867
rect 19150 51864 19156 51876
rect 17819 51836 19156 51864
rect 17819 51833 17831 51836
rect 17773 51827 17831 51833
rect 19150 51824 19156 51836
rect 19208 51824 19214 51876
rect 24210 51864 24216 51876
rect 19306 51836 24216 51864
rect 15746 51756 15752 51808
rect 15804 51796 15810 51808
rect 16117 51799 16175 51805
rect 16117 51796 16129 51799
rect 15804 51768 16129 51796
rect 15804 51756 15810 51768
rect 16117 51765 16129 51768
rect 16163 51796 16175 51799
rect 19306 51796 19334 51836
rect 24210 51824 24216 51836
rect 24268 51824 24274 51876
rect 25406 51824 25412 51876
rect 25464 51864 25470 51876
rect 25593 51867 25651 51873
rect 25593 51864 25605 51867
rect 25464 51836 25605 51864
rect 25464 51824 25470 51836
rect 25593 51833 25605 51836
rect 25639 51833 25651 51867
rect 25593 51827 25651 51833
rect 26970 51824 26976 51876
rect 27028 51864 27034 51876
rect 27908 51864 27936 51972
rect 28169 51969 28181 51972
rect 28215 51969 28227 52003
rect 28169 51963 28227 51969
rect 28353 52003 28411 52009
rect 28353 51969 28365 52003
rect 28399 52000 28411 52003
rect 28460 52000 28488 52028
rect 28399 51972 28488 52000
rect 28721 52003 28779 52009
rect 28399 51969 28411 51972
rect 28353 51963 28411 51969
rect 28721 51969 28733 52003
rect 28767 52000 28779 52003
rect 29178 52000 29184 52012
rect 28767 51972 29184 52000
rect 28767 51969 28779 51972
rect 28721 51963 28779 51969
rect 29178 51960 29184 51972
rect 29236 51960 29242 52012
rect 29564 52009 29592 52040
rect 29638 52028 29644 52080
rect 29696 52068 29702 52080
rect 29696 52040 29960 52068
rect 29696 52028 29702 52040
rect 29932 52009 29960 52040
rect 30006 52028 30012 52080
rect 30064 52068 30070 52080
rect 30466 52068 30472 52080
rect 30064 52040 30472 52068
rect 30064 52028 30070 52040
rect 30466 52028 30472 52040
rect 30524 52028 30530 52080
rect 29365 52003 29423 52009
rect 29365 51969 29377 52003
rect 29411 51969 29423 52003
rect 29365 51963 29423 51969
rect 29549 52003 29607 52009
rect 29549 51969 29561 52003
rect 29595 51969 29607 52003
rect 29549 51963 29607 51969
rect 29917 52003 29975 52009
rect 29917 51969 29929 52003
rect 29963 51969 29975 52003
rect 29917 51963 29975 51969
rect 28445 51935 28503 51941
rect 28445 51932 28457 51935
rect 27028 51836 27936 51864
rect 28205 51904 28457 51932
rect 27028 51824 27034 51836
rect 16163 51768 19334 51796
rect 16163 51765 16175 51768
rect 16117 51759 16175 51765
rect 23842 51756 23848 51808
rect 23900 51796 23906 51808
rect 28205 51796 28233 51904
rect 28445 51901 28457 51904
rect 28491 51901 28503 51935
rect 28445 51895 28503 51901
rect 28537 51935 28595 51941
rect 28537 51901 28549 51935
rect 28583 51932 28595 51935
rect 28902 51932 28908 51944
rect 28583 51904 28908 51932
rect 28583 51901 28595 51904
rect 28537 51895 28595 51901
rect 28902 51892 28908 51904
rect 28960 51892 28966 51944
rect 29270 51892 29276 51944
rect 29328 51932 29334 51944
rect 29380 51932 29408 51963
rect 29638 51932 29644 51944
rect 29328 51904 29408 51932
rect 29599 51904 29644 51932
rect 29328 51892 29334 51904
rect 29638 51892 29644 51904
rect 29696 51892 29702 51944
rect 29733 51935 29791 51941
rect 29733 51901 29745 51935
rect 29779 51901 29791 51935
rect 29733 51895 29791 51901
rect 29748 51864 29776 51895
rect 29656 51836 29776 51864
rect 23900 51768 28233 51796
rect 28905 51799 28963 51805
rect 23900 51756 23906 51768
rect 28905 51765 28917 51799
rect 28951 51796 28963 51799
rect 29086 51796 29092 51808
rect 28951 51768 29092 51796
rect 28951 51765 28963 51768
rect 28905 51759 28963 51765
rect 29086 51756 29092 51768
rect 29144 51756 29150 51808
rect 29454 51756 29460 51808
rect 29512 51796 29518 51808
rect 29656 51796 29684 51836
rect 29512 51768 29684 51796
rect 29512 51756 29518 51768
rect 1104 51706 30820 51728
rect 1104 51654 5915 51706
rect 5967 51654 5979 51706
rect 6031 51654 6043 51706
rect 6095 51654 6107 51706
rect 6159 51654 6171 51706
rect 6223 51654 15846 51706
rect 15898 51654 15910 51706
rect 15962 51654 15974 51706
rect 16026 51654 16038 51706
rect 16090 51654 16102 51706
rect 16154 51654 25776 51706
rect 25828 51654 25840 51706
rect 25892 51654 25904 51706
rect 25956 51654 25968 51706
rect 26020 51654 26032 51706
rect 26084 51654 30820 51706
rect 1104 51632 30820 51654
rect 12618 51552 12624 51604
rect 12676 51592 12682 51604
rect 12989 51595 13047 51601
rect 12989 51592 13001 51595
rect 12676 51564 13001 51592
rect 12676 51552 12682 51564
rect 12989 51561 13001 51564
rect 13035 51561 13047 51595
rect 14458 51592 14464 51604
rect 14419 51564 14464 51592
rect 12989 51555 13047 51561
rect 14458 51552 14464 51564
rect 14516 51552 14522 51604
rect 14734 51552 14740 51604
rect 14792 51592 14798 51604
rect 15749 51595 15807 51601
rect 15749 51592 15761 51595
rect 14792 51564 15761 51592
rect 14792 51552 14798 51564
rect 15749 51561 15761 51564
rect 15795 51561 15807 51595
rect 17954 51592 17960 51604
rect 17915 51564 17960 51592
rect 15749 51555 15807 51561
rect 17954 51552 17960 51564
rect 18012 51552 18018 51604
rect 19334 51592 19340 51604
rect 19295 51564 19340 51592
rect 19334 51552 19340 51564
rect 19392 51552 19398 51604
rect 19518 51552 19524 51604
rect 19576 51592 19582 51604
rect 20533 51595 20591 51601
rect 20533 51592 20545 51595
rect 19576 51564 20545 51592
rect 19576 51552 19582 51564
rect 20533 51561 20545 51564
rect 20579 51561 20591 51595
rect 20533 51555 20591 51561
rect 22186 51552 22192 51604
rect 22244 51592 22250 51604
rect 22281 51595 22339 51601
rect 22281 51592 22293 51595
rect 22244 51564 22293 51592
rect 22244 51552 22250 51564
rect 22281 51561 22293 51564
rect 22327 51561 22339 51595
rect 22281 51555 22339 51561
rect 27614 51552 27620 51604
rect 27672 51592 27678 51604
rect 29638 51592 29644 51604
rect 27672 51564 29644 51592
rect 27672 51552 27678 51564
rect 29638 51552 29644 51564
rect 29696 51552 29702 51604
rect 25314 51484 25320 51536
rect 25372 51524 25378 51536
rect 25958 51524 25964 51536
rect 25372 51496 25964 51524
rect 25372 51484 25378 51496
rect 25958 51484 25964 51496
rect 26016 51484 26022 51536
rect 29454 51484 29460 51536
rect 29512 51524 29518 51536
rect 30466 51524 30472 51536
rect 29512 51496 30472 51524
rect 29512 51484 29518 51496
rect 30466 51484 30472 51496
rect 30524 51484 30530 51536
rect 15746 51456 15752 51468
rect 14752 51428 15752 51456
rect 1394 51348 1400 51400
rect 1452 51388 1458 51400
rect 1581 51391 1639 51397
rect 1581 51388 1593 51391
rect 1452 51360 1593 51388
rect 1452 51348 1458 51360
rect 1581 51357 1593 51360
rect 1627 51357 1639 51391
rect 2222 51388 2228 51400
rect 2183 51360 2228 51388
rect 1581 51351 1639 51357
rect 2222 51348 2228 51360
rect 2280 51348 2286 51400
rect 12805 51391 12863 51397
rect 12805 51357 12817 51391
rect 12851 51388 12863 51391
rect 14642 51388 14648 51400
rect 12851 51360 14648 51388
rect 12851 51357 12863 51360
rect 12805 51351 12863 51357
rect 14642 51348 14648 51360
rect 14700 51348 14706 51400
rect 14752 51397 14780 51428
rect 15746 51416 15752 51428
rect 15804 51416 15810 51468
rect 18322 51416 18328 51468
rect 18380 51456 18386 51468
rect 18693 51459 18751 51465
rect 18693 51456 18705 51459
rect 18380 51428 18705 51456
rect 18380 51416 18386 51428
rect 18693 51425 18705 51428
rect 18739 51456 18751 51459
rect 19886 51456 19892 51468
rect 18739 51428 19892 51456
rect 18739 51425 18751 51428
rect 18693 51419 18751 51425
rect 19886 51416 19892 51428
rect 19944 51456 19950 51468
rect 21085 51459 21143 51465
rect 21085 51456 21097 51459
rect 19944 51428 21097 51456
rect 19944 51416 19950 51428
rect 21085 51425 21097 51428
rect 21131 51425 21143 51459
rect 23290 51456 23296 51468
rect 21085 51419 21143 51425
rect 22572 51428 23296 51456
rect 14737 51391 14795 51397
rect 14737 51357 14749 51391
rect 14783 51357 14795 51391
rect 14737 51351 14795 51357
rect 14829 51391 14887 51397
rect 14829 51357 14841 51391
rect 14875 51357 14887 51391
rect 14829 51351 14887 51357
rect 14366 51280 14372 51332
rect 14424 51320 14430 51332
rect 14844 51320 14872 51351
rect 14918 51348 14924 51400
rect 14976 51388 14982 51400
rect 15105 51391 15163 51397
rect 14976 51360 15021 51388
rect 14976 51348 14982 51360
rect 15105 51357 15117 51391
rect 15151 51357 15163 51391
rect 15105 51351 15163 51357
rect 14424 51292 14872 51320
rect 14424 51280 14430 51292
rect 1397 51255 1455 51261
rect 1397 51221 1409 51255
rect 1443 51252 1455 51255
rect 1762 51252 1768 51264
rect 1443 51224 1768 51252
rect 1443 51221 1455 51224
rect 1397 51215 1455 51221
rect 1762 51212 1768 51224
rect 1820 51212 1826 51264
rect 2038 51252 2044 51264
rect 1999 51224 2044 51252
rect 2038 51212 2044 51224
rect 2096 51212 2102 51264
rect 12618 51212 12624 51264
rect 12676 51252 12682 51264
rect 15120 51252 15148 51351
rect 15378 51348 15384 51400
rect 15436 51388 15442 51400
rect 15565 51391 15623 51397
rect 15565 51388 15577 51391
rect 15436 51360 15577 51388
rect 15436 51348 15442 51360
rect 15565 51357 15577 51360
rect 15611 51357 15623 51391
rect 15565 51351 15623 51357
rect 17678 51348 17684 51400
rect 17736 51388 17742 51400
rect 17773 51391 17831 51397
rect 17773 51388 17785 51391
rect 17736 51360 17785 51388
rect 17736 51348 17742 51360
rect 17773 51357 17785 51360
rect 17819 51357 17831 51391
rect 17773 51351 17831 51357
rect 19613 51391 19671 51397
rect 19613 51357 19625 51391
rect 19659 51388 19671 51391
rect 20622 51388 20628 51400
rect 19659 51360 20628 51388
rect 19659 51357 19671 51360
rect 19613 51351 19671 51357
rect 20622 51348 20628 51360
rect 20680 51388 20686 51400
rect 20809 51391 20867 51397
rect 20809 51388 20821 51391
rect 20680 51360 20821 51388
rect 20680 51348 20686 51360
rect 20809 51357 20821 51360
rect 20855 51357 20867 51391
rect 22462 51388 22468 51400
rect 22423 51360 22468 51388
rect 20809 51351 20867 51357
rect 22462 51348 22468 51360
rect 22520 51348 22526 51400
rect 22572 51397 22600 51428
rect 23290 51416 23296 51428
rect 23348 51416 23354 51468
rect 24026 51416 24032 51468
rect 24084 51456 24090 51468
rect 24394 51456 24400 51468
rect 24084 51428 24400 51456
rect 24084 51416 24090 51428
rect 24394 51416 24400 51428
rect 24452 51456 24458 51468
rect 25593 51459 25651 51465
rect 24452 51428 24716 51456
rect 24452 51416 24458 51428
rect 22557 51391 22615 51397
rect 22557 51357 22569 51391
rect 22603 51357 22615 51391
rect 22557 51351 22615 51357
rect 22646 51348 22652 51400
rect 22704 51388 22710 51400
rect 22741 51391 22799 51397
rect 22741 51388 22753 51391
rect 22704 51360 22753 51388
rect 22704 51348 22710 51360
rect 22741 51357 22753 51360
rect 22787 51357 22799 51391
rect 22741 51351 22799 51357
rect 22830 51348 22836 51400
rect 22888 51388 22894 51400
rect 24578 51388 24584 51400
rect 22888 51360 22933 51388
rect 24539 51360 24584 51388
rect 22888 51348 22894 51360
rect 24578 51348 24584 51360
rect 24636 51348 24642 51400
rect 24688 51388 24716 51428
rect 25593 51425 25605 51459
rect 25639 51456 25651 51459
rect 26142 51456 26148 51468
rect 25639 51428 26148 51456
rect 25639 51425 25651 51428
rect 25593 51419 25651 51425
rect 26142 51416 26148 51428
rect 26200 51416 26206 51468
rect 29362 51416 29368 51468
rect 29420 51416 29426 51468
rect 24688 51360 25268 51388
rect 17218 51280 17224 51332
rect 17276 51320 17282 51332
rect 18509 51323 18567 51329
rect 18509 51320 18521 51323
rect 17276 51292 18521 51320
rect 17276 51280 17282 51292
rect 18509 51289 18521 51292
rect 18555 51289 18567 51323
rect 19794 51320 19800 51332
rect 19755 51292 19800 51320
rect 18509 51283 18567 51289
rect 12676 51224 15148 51252
rect 18524 51252 18552 51283
rect 19794 51280 19800 51292
rect 19852 51280 19858 51332
rect 24394 51320 24400 51332
rect 24355 51292 24400 51320
rect 24394 51280 24400 51292
rect 24452 51280 24458 51332
rect 20622 51252 20628 51264
rect 18524 51224 20628 51252
rect 12676 51212 12682 51224
rect 20622 51212 20628 51224
rect 20680 51212 20686 51264
rect 20993 51255 21051 51261
rect 20993 51221 21005 51255
rect 21039 51252 21051 51255
rect 21358 51252 21364 51264
rect 21039 51224 21364 51252
rect 21039 51221 21051 51224
rect 20993 51215 21051 51221
rect 21358 51212 21364 51224
rect 21416 51212 21422 51264
rect 23382 51212 23388 51264
rect 23440 51252 23446 51264
rect 24486 51252 24492 51264
rect 23440 51224 24492 51252
rect 23440 51212 23446 51224
rect 24486 51212 24492 51224
rect 24544 51212 24550 51264
rect 24688 51261 24716 51360
rect 24946 51320 24952 51332
rect 24907 51292 24952 51320
rect 24946 51280 24952 51292
rect 25004 51280 25010 51332
rect 24673 51255 24731 51261
rect 24673 51221 24685 51255
rect 24719 51221 24731 51255
rect 24673 51215 24731 51221
rect 24762 51212 24768 51264
rect 24820 51252 24826 51264
rect 25240 51252 25268 51360
rect 25314 51348 25320 51400
rect 25372 51388 25378 51400
rect 28718 51388 28724 51400
rect 25372 51360 26188 51388
rect 28679 51360 28724 51388
rect 25372 51348 25378 51360
rect 25590 51280 25596 51332
rect 25648 51320 25654 51332
rect 25777 51323 25835 51329
rect 25777 51320 25789 51323
rect 25648 51292 25789 51320
rect 25648 51280 25654 51292
rect 25777 51289 25789 51292
rect 25823 51289 25835 51323
rect 26050 51320 26056 51332
rect 25777 51283 25835 51289
rect 25884 51292 26056 51320
rect 25884 51261 25912 51292
rect 26050 51280 26056 51292
rect 26108 51280 26114 51332
rect 26160 51329 26188 51360
rect 28718 51348 28724 51360
rect 28776 51348 28782 51400
rect 26145 51323 26203 51329
rect 26145 51289 26157 51323
rect 26191 51289 26203 51323
rect 26145 51283 26203 51289
rect 27614 51280 27620 51332
rect 27672 51320 27678 51332
rect 27798 51320 27804 51332
rect 27672 51292 27804 51320
rect 27672 51280 27678 51292
rect 27798 51280 27804 51292
rect 27856 51280 27862 51332
rect 25869 51255 25927 51261
rect 25869 51252 25881 51255
rect 24820 51224 24865 51252
rect 25240 51224 25881 51252
rect 24820 51212 24826 51224
rect 25869 51221 25881 51224
rect 25915 51221 25927 51255
rect 25869 51215 25927 51221
rect 25961 51255 26019 51261
rect 25961 51221 25973 51255
rect 26007 51252 26019 51255
rect 26326 51252 26332 51264
rect 26007 51224 26332 51252
rect 26007 51221 26019 51224
rect 25961 51215 26019 51221
rect 26326 51212 26332 51224
rect 26384 51212 26390 51264
rect 28902 51252 28908 51264
rect 28863 51224 28908 51252
rect 28902 51212 28908 51224
rect 28960 51212 28966 51264
rect 29086 51212 29092 51264
rect 29144 51252 29150 51264
rect 29380 51252 29408 51416
rect 29733 51323 29791 51329
rect 29733 51289 29745 51323
rect 29779 51320 29791 51323
rect 29914 51320 29920 51332
rect 29779 51292 29920 51320
rect 29779 51289 29791 51292
rect 29733 51283 29791 51289
rect 29914 51280 29920 51292
rect 29972 51280 29978 51332
rect 29825 51255 29883 51261
rect 29825 51252 29837 51255
rect 29144 51224 29837 51252
rect 29144 51212 29150 51224
rect 29825 51221 29837 51224
rect 29871 51221 29883 51255
rect 29825 51215 29883 51221
rect 30282 51212 30288 51264
rect 30340 51252 30346 51264
rect 30466 51252 30472 51264
rect 30340 51224 30472 51252
rect 30340 51212 30346 51224
rect 30466 51212 30472 51224
rect 30524 51212 30530 51264
rect 1104 51162 30820 51184
rect 1104 51110 10880 51162
rect 10932 51110 10944 51162
rect 10996 51110 11008 51162
rect 11060 51110 11072 51162
rect 11124 51110 11136 51162
rect 11188 51110 20811 51162
rect 20863 51110 20875 51162
rect 20927 51110 20939 51162
rect 20991 51110 21003 51162
rect 21055 51110 21067 51162
rect 21119 51110 30820 51162
rect 1104 51088 30820 51110
rect 14918 51008 14924 51060
rect 14976 51048 14982 51060
rect 17497 51051 17555 51057
rect 14976 51020 15148 51048
rect 14976 51008 14982 51020
rect 14366 50940 14372 50992
rect 14424 50980 14430 50992
rect 14424 50952 15056 50980
rect 14424 50940 14430 50952
rect 1578 50912 1584 50924
rect 1539 50884 1584 50912
rect 1578 50872 1584 50884
rect 1636 50872 1642 50924
rect 14918 50912 14924 50924
rect 14879 50884 14924 50912
rect 14918 50872 14924 50884
rect 14976 50872 14982 50924
rect 15028 50921 15056 50952
rect 15120 50924 15148 51020
rect 17497 51017 17509 51051
rect 17543 51048 17555 51051
rect 19702 51048 19708 51060
rect 17543 51020 19708 51048
rect 17543 51017 17555 51020
rect 17497 51011 17555 51017
rect 19702 51008 19708 51020
rect 19760 51048 19766 51060
rect 20346 51048 20352 51060
rect 19760 51020 20352 51048
rect 19760 51008 19766 51020
rect 20346 51008 20352 51020
rect 20404 51008 20410 51060
rect 22370 51048 22376 51060
rect 21376 51020 22376 51048
rect 19426 50980 19432 50992
rect 15396 50952 19432 50980
rect 15013 50915 15071 50921
rect 15013 50881 15025 50915
rect 15059 50881 15071 50915
rect 15013 50875 15071 50881
rect 15102 50872 15108 50924
rect 15160 50912 15166 50924
rect 15289 50915 15347 50921
rect 15160 50884 15205 50912
rect 15160 50872 15166 50884
rect 15289 50881 15301 50915
rect 15335 50881 15347 50915
rect 15289 50875 15347 50881
rect 13722 50804 13728 50856
rect 13780 50844 13786 50856
rect 15304 50844 15332 50875
rect 13780 50816 15332 50844
rect 13780 50804 13786 50816
rect 1854 50736 1860 50788
rect 1912 50776 1918 50788
rect 15396 50776 15424 50952
rect 19426 50940 19432 50952
rect 19484 50940 19490 50992
rect 20073 50983 20131 50989
rect 20073 50949 20085 50983
rect 20119 50980 20131 50983
rect 21266 50980 21272 50992
rect 20119 50952 21272 50980
rect 20119 50949 20131 50952
rect 20073 50943 20131 50949
rect 21266 50940 21272 50952
rect 21324 50940 21330 50992
rect 17310 50912 17316 50924
rect 17271 50884 17316 50912
rect 17310 50872 17316 50884
rect 17368 50872 17374 50924
rect 15470 50804 15476 50856
rect 15528 50844 15534 50856
rect 21376 50844 21404 51020
rect 22370 51008 22376 51020
rect 22428 51008 22434 51060
rect 22462 51008 22468 51060
rect 22520 51048 22526 51060
rect 22649 51051 22707 51057
rect 22649 51048 22661 51051
rect 22520 51020 22661 51048
rect 22520 51008 22526 51020
rect 22649 51017 22661 51020
rect 22695 51017 22707 51051
rect 22649 51011 22707 51017
rect 23934 51008 23940 51060
rect 23992 51048 23998 51060
rect 24210 51048 24216 51060
rect 23992 51020 24216 51048
rect 23992 51008 23998 51020
rect 24210 51008 24216 51020
rect 24268 51008 24274 51060
rect 24489 51051 24547 51057
rect 24489 51017 24501 51051
rect 24535 51017 24547 51051
rect 24673 51051 24731 51057
rect 24673 51048 24685 51051
rect 24489 51011 24547 51017
rect 24596 51020 24685 51048
rect 22094 50940 22100 50992
rect 22152 50980 22158 50992
rect 22152 50952 22197 50980
rect 22152 50940 22158 50952
rect 23290 50940 23296 50992
rect 23348 50980 23354 50992
rect 24504 50980 24532 51011
rect 23348 50952 24532 50980
rect 23348 50940 23354 50952
rect 21913 50915 21971 50921
rect 21913 50881 21925 50915
rect 21959 50912 21971 50915
rect 22278 50912 22284 50924
rect 21959 50884 22284 50912
rect 21959 50881 21971 50884
rect 21913 50875 21971 50881
rect 22278 50872 22284 50884
rect 22336 50872 22342 50924
rect 22557 50915 22615 50921
rect 22557 50881 22569 50915
rect 22603 50881 22615 50915
rect 22557 50875 22615 50881
rect 15528 50816 21404 50844
rect 15528 50804 15534 50816
rect 22186 50804 22192 50856
rect 22244 50844 22250 50856
rect 22572 50844 22600 50875
rect 22244 50816 22600 50844
rect 22244 50804 22250 50816
rect 1912 50748 15424 50776
rect 1912 50736 1918 50748
rect 15562 50736 15568 50788
rect 15620 50776 15626 50788
rect 21910 50776 21916 50788
rect 15620 50748 21916 50776
rect 15620 50736 15626 50748
rect 21910 50736 21916 50748
rect 21968 50736 21974 50788
rect 22002 50736 22008 50788
rect 22060 50776 22066 50788
rect 23308 50776 23336 50940
rect 23474 50872 23480 50924
rect 23532 50912 23538 50924
rect 24305 50915 24363 50921
rect 23532 50910 24256 50912
rect 24305 50910 24317 50915
rect 23532 50884 24317 50910
rect 23532 50872 23538 50884
rect 24228 50882 24317 50884
rect 24305 50881 24317 50882
rect 24351 50881 24363 50915
rect 24305 50875 24363 50881
rect 24486 50872 24492 50924
rect 24544 50912 24550 50924
rect 24596 50912 24624 51020
rect 24673 51017 24685 51020
rect 24719 51017 24731 51051
rect 24673 51011 24731 51017
rect 25501 51051 25559 51057
rect 25501 51017 25513 51051
rect 25547 51017 25559 51051
rect 25501 51011 25559 51017
rect 25593 51051 25651 51057
rect 25593 51017 25605 51051
rect 25639 51048 25651 51051
rect 25774 51048 25780 51060
rect 25639 51020 25780 51048
rect 25639 51017 25651 51020
rect 25593 51011 25651 51017
rect 25516 50980 25544 51011
rect 25774 51008 25780 51020
rect 25832 51008 25838 51060
rect 25958 51008 25964 51060
rect 26016 51048 26022 51060
rect 26418 51048 26424 51060
rect 26016 51020 26424 51048
rect 26016 51008 26022 51020
rect 26418 51008 26424 51020
rect 26476 51008 26482 51060
rect 29546 51048 29552 51060
rect 29012 51020 29552 51048
rect 26050 50980 26056 50992
rect 25516 50952 26056 50980
rect 26050 50940 26056 50952
rect 26108 50940 26114 50992
rect 25409 50915 25467 50921
rect 25409 50912 25421 50915
rect 24544 50884 24624 50912
rect 24688 50884 25421 50912
rect 24544 50872 24550 50884
rect 23382 50804 23388 50856
rect 23440 50844 23446 50856
rect 24397 50847 24455 50853
rect 24397 50844 24409 50847
rect 23440 50816 24409 50844
rect 23440 50804 23446 50816
rect 24397 50813 24409 50816
rect 24443 50813 24455 50847
rect 24397 50807 24455 50813
rect 22060 50748 23336 50776
rect 22060 50736 22066 50748
rect 23750 50736 23756 50788
rect 23808 50776 23814 50788
rect 24688 50776 24716 50884
rect 25409 50881 25421 50884
rect 25455 50881 25467 50915
rect 25409 50875 25467 50881
rect 25498 50872 25504 50924
rect 25556 50912 25562 50924
rect 25777 50915 25835 50921
rect 25777 50912 25789 50915
rect 25556 50884 25789 50912
rect 25556 50872 25562 50884
rect 25777 50881 25789 50884
rect 25823 50881 25835 50915
rect 25777 50875 25835 50881
rect 28810 50872 28816 50924
rect 28868 50912 28874 50924
rect 28905 50915 28963 50921
rect 28905 50912 28917 50915
rect 28868 50884 28917 50912
rect 28868 50872 28874 50884
rect 28905 50881 28917 50884
rect 28951 50881 28963 50915
rect 28905 50875 28963 50881
rect 29012 50856 29040 51020
rect 29546 51008 29552 51020
rect 29604 51008 29610 51060
rect 30834 51008 30840 51060
rect 30892 51048 30898 51060
rect 30892 51020 31892 51048
rect 30892 51008 30898 51020
rect 29638 50940 29644 50992
rect 29696 50980 29702 50992
rect 29822 50980 29828 50992
rect 29696 50952 29828 50980
rect 29696 50940 29702 50952
rect 29822 50940 29828 50952
rect 29880 50940 29886 50992
rect 29733 50915 29791 50921
rect 29733 50881 29745 50915
rect 29779 50912 29791 50915
rect 29779 50884 30328 50912
rect 29779 50881 29791 50884
rect 29733 50875 29791 50881
rect 24765 50847 24823 50853
rect 24765 50813 24777 50847
rect 24811 50844 24823 50847
rect 24854 50844 24860 50856
rect 24811 50816 24860 50844
rect 24811 50813 24823 50816
rect 24765 50807 24823 50813
rect 24854 50804 24860 50816
rect 24912 50804 24918 50856
rect 28994 50804 29000 50856
rect 29052 50804 29058 50856
rect 30300 50844 30328 50884
rect 31864 50856 31892 51020
rect 30926 50844 30932 50856
rect 30300 50816 30932 50844
rect 30926 50804 30932 50816
rect 30984 50804 30990 50856
rect 31846 50804 31852 50856
rect 31904 50804 31910 50856
rect 23808 50748 24716 50776
rect 23808 50736 23814 50748
rect 24946 50736 24952 50788
rect 25004 50736 25010 50788
rect 25225 50779 25283 50785
rect 25225 50745 25237 50779
rect 25271 50776 25283 50779
rect 25774 50776 25780 50788
rect 25271 50748 25780 50776
rect 25271 50745 25283 50748
rect 25225 50739 25283 50745
rect 25774 50736 25780 50748
rect 25832 50736 25838 50788
rect 30098 50736 30104 50788
rect 30156 50736 30162 50788
rect 1397 50711 1455 50717
rect 1397 50677 1409 50711
rect 1443 50708 1455 50711
rect 1670 50708 1676 50720
rect 1443 50680 1676 50708
rect 1443 50677 1455 50680
rect 1397 50671 1455 50677
rect 1670 50668 1676 50680
rect 1728 50668 1734 50720
rect 14645 50711 14703 50717
rect 14645 50677 14657 50711
rect 14691 50708 14703 50711
rect 15746 50708 15752 50720
rect 14691 50680 15752 50708
rect 14691 50677 14703 50680
rect 14645 50671 14703 50677
rect 15746 50668 15752 50680
rect 15804 50668 15810 50720
rect 20162 50708 20168 50720
rect 20123 50680 20168 50708
rect 20162 50668 20168 50680
rect 20220 50668 20226 50720
rect 22094 50668 22100 50720
rect 22152 50708 22158 50720
rect 22738 50708 22744 50720
rect 22152 50680 22744 50708
rect 22152 50668 22158 50680
rect 22738 50668 22744 50680
rect 22796 50668 22802 50720
rect 24121 50711 24179 50717
rect 24121 50677 24133 50711
rect 24167 50708 24179 50711
rect 24964 50708 24992 50736
rect 29086 50708 29092 50720
rect 24167 50680 24992 50708
rect 29047 50680 29092 50708
rect 24167 50677 24179 50680
rect 24121 50671 24179 50677
rect 29086 50668 29092 50680
rect 29144 50668 29150 50720
rect 29822 50708 29828 50720
rect 29783 50680 29828 50708
rect 29822 50668 29828 50680
rect 29880 50668 29886 50720
rect 29914 50668 29920 50720
rect 29972 50708 29978 50720
rect 30116 50708 30144 50736
rect 29972 50680 30144 50708
rect 29972 50668 29978 50680
rect 1104 50618 30820 50640
rect 1104 50566 5915 50618
rect 5967 50566 5979 50618
rect 6031 50566 6043 50618
rect 6095 50566 6107 50618
rect 6159 50566 6171 50618
rect 6223 50566 15846 50618
rect 15898 50566 15910 50618
rect 15962 50566 15974 50618
rect 16026 50566 16038 50618
rect 16090 50566 16102 50618
rect 16154 50566 25776 50618
rect 25828 50566 25840 50618
rect 25892 50566 25904 50618
rect 25956 50566 25968 50618
rect 26020 50566 26032 50618
rect 26084 50566 30820 50618
rect 1104 50544 30820 50566
rect 2682 50504 2688 50516
rect 2643 50476 2688 50504
rect 2682 50464 2688 50476
rect 2740 50464 2746 50516
rect 19889 50507 19947 50513
rect 19889 50473 19901 50507
rect 19935 50504 19947 50507
rect 21450 50504 21456 50516
rect 19935 50476 21456 50504
rect 19935 50473 19947 50476
rect 19889 50467 19947 50473
rect 21450 50464 21456 50476
rect 21508 50464 21514 50516
rect 21726 50504 21732 50516
rect 21687 50476 21732 50504
rect 21726 50464 21732 50476
rect 21784 50464 21790 50516
rect 22370 50464 22376 50516
rect 22428 50504 22434 50516
rect 22428 50476 24440 50504
rect 22428 50464 22434 50476
rect 21634 50396 21640 50448
rect 21692 50436 21698 50448
rect 21692 50408 22692 50436
rect 21692 50396 21698 50408
rect 22066 50340 22600 50368
rect 1486 50260 1492 50312
rect 1544 50300 1550 50312
rect 1765 50303 1823 50309
rect 1765 50300 1777 50303
rect 1544 50272 1777 50300
rect 1544 50260 1550 50272
rect 1765 50269 1777 50272
rect 1811 50269 1823 50303
rect 1765 50263 1823 50269
rect 2038 50260 2044 50312
rect 2096 50300 2102 50312
rect 2593 50303 2651 50309
rect 2593 50300 2605 50303
rect 2096 50272 2605 50300
rect 2096 50260 2102 50272
rect 2593 50269 2605 50272
rect 2639 50269 2651 50303
rect 2593 50263 2651 50269
rect 11793 50303 11851 50309
rect 11793 50269 11805 50303
rect 11839 50300 11851 50303
rect 11882 50300 11888 50312
rect 11839 50272 11888 50300
rect 11839 50269 11851 50272
rect 11793 50263 11851 50269
rect 11882 50260 11888 50272
rect 11940 50260 11946 50312
rect 15470 50300 15476 50312
rect 11992 50272 15476 50300
rect 1581 50235 1639 50241
rect 1581 50201 1593 50235
rect 1627 50201 1639 50235
rect 1581 50195 1639 50201
rect 1486 50124 1492 50176
rect 1544 50164 1550 50176
rect 1596 50164 1624 50195
rect 1854 50192 1860 50244
rect 1912 50232 1918 50244
rect 1949 50235 2007 50241
rect 1949 50232 1961 50235
rect 1912 50204 1961 50232
rect 1912 50192 1918 50204
rect 1949 50201 1961 50204
rect 1995 50201 2007 50235
rect 1949 50195 2007 50201
rect 2409 50235 2467 50241
rect 2409 50201 2421 50235
rect 2455 50201 2467 50235
rect 2409 50195 2467 50201
rect 2424 50164 2452 50195
rect 10502 50192 10508 50244
rect 10560 50232 10566 50244
rect 11992 50232 12020 50272
rect 15470 50260 15476 50272
rect 15528 50260 15534 50312
rect 15565 50303 15623 50309
rect 15565 50269 15577 50303
rect 15611 50300 15623 50303
rect 15654 50300 15660 50312
rect 15611 50272 15660 50300
rect 15611 50269 15623 50272
rect 15565 50263 15623 50269
rect 15654 50260 15660 50272
rect 15712 50260 15718 50312
rect 15838 50309 15844 50312
rect 15832 50300 15844 50309
rect 15799 50272 15844 50300
rect 15832 50263 15844 50272
rect 15838 50260 15844 50263
rect 15896 50260 15902 50312
rect 19702 50300 19708 50312
rect 19663 50272 19708 50300
rect 19702 50260 19708 50272
rect 19760 50260 19766 50312
rect 19978 50260 19984 50312
rect 20036 50300 20042 50312
rect 20349 50303 20407 50309
rect 20349 50300 20361 50303
rect 20036 50272 20361 50300
rect 20036 50260 20042 50272
rect 20349 50269 20361 50272
rect 20395 50269 20407 50303
rect 21082 50300 21088 50312
rect 20349 50263 20407 50269
rect 20456 50272 21088 50300
rect 10560 50204 12020 50232
rect 12060 50235 12118 50241
rect 10560 50192 10566 50204
rect 12060 50201 12072 50235
rect 12106 50232 12118 50235
rect 12250 50232 12256 50244
rect 12106 50204 12256 50232
rect 12106 50201 12118 50204
rect 12060 50195 12118 50201
rect 12250 50192 12256 50204
rect 12308 50192 12314 50244
rect 20456 50232 20484 50272
rect 21082 50260 21088 50272
rect 21140 50260 21146 50312
rect 21634 50260 21640 50312
rect 21692 50300 21698 50312
rect 22066 50300 22094 50340
rect 22462 50300 22468 50312
rect 21692 50272 22094 50300
rect 22423 50272 22468 50300
rect 21692 50260 21698 50272
rect 22462 50260 22468 50272
rect 22520 50260 22526 50312
rect 22572 50309 22600 50340
rect 22664 50309 22692 50408
rect 23014 50396 23020 50448
rect 23072 50436 23078 50448
rect 23934 50436 23940 50448
rect 23072 50408 23940 50436
rect 23072 50396 23078 50408
rect 22557 50303 22615 50309
rect 22557 50269 22569 50303
rect 22603 50269 22615 50303
rect 22557 50263 22615 50269
rect 22649 50303 22707 50309
rect 22649 50269 22661 50303
rect 22695 50269 22707 50303
rect 22649 50263 22707 50269
rect 22833 50303 22891 50309
rect 22833 50269 22845 50303
rect 22879 50300 22891 50303
rect 23014 50300 23020 50312
rect 22879 50272 23020 50300
rect 22879 50269 22891 50272
rect 22833 50263 22891 50269
rect 23014 50260 23020 50272
rect 23072 50260 23078 50312
rect 13188 50204 20484 50232
rect 20616 50235 20674 50241
rect 1544 50136 2452 50164
rect 1544 50124 1550 50136
rect 13078 50124 13084 50176
rect 13136 50164 13142 50176
rect 13188 50173 13216 50204
rect 20616 50201 20628 50235
rect 20662 50232 20674 50235
rect 22189 50235 22247 50241
rect 22189 50232 22201 50235
rect 20662 50204 22201 50232
rect 20662 50201 20674 50204
rect 20616 50195 20674 50201
rect 22189 50201 22201 50204
rect 22235 50201 22247 50235
rect 23400 50232 23428 50408
rect 23934 50396 23940 50408
rect 23992 50396 23998 50448
rect 24412 50445 24440 50476
rect 24762 50464 24768 50516
rect 24820 50504 24826 50516
rect 25222 50504 25228 50516
rect 24820 50476 25228 50504
rect 24820 50464 24826 50476
rect 25222 50464 25228 50476
rect 25280 50464 25286 50516
rect 24397 50439 24455 50445
rect 24397 50405 24409 50439
rect 24443 50405 24455 50439
rect 24397 50399 24455 50405
rect 24578 50396 24584 50448
rect 24636 50436 24642 50448
rect 24946 50436 24952 50448
rect 24636 50408 24952 50436
rect 24636 50396 24642 50408
rect 24946 50396 24952 50408
rect 25004 50396 25010 50448
rect 27890 50396 27896 50448
rect 27948 50436 27954 50448
rect 28166 50436 28172 50448
rect 27948 50408 28172 50436
rect 27948 50396 27954 50408
rect 28166 50396 28172 50408
rect 28224 50396 28230 50448
rect 23750 50368 23756 50380
rect 23492 50340 23756 50368
rect 23492 50309 23520 50340
rect 23750 50328 23756 50340
rect 23808 50368 23814 50380
rect 23808 50340 24624 50368
rect 23808 50328 23814 50340
rect 23477 50303 23535 50309
rect 23477 50269 23489 50303
rect 23523 50269 23535 50303
rect 23845 50303 23903 50309
rect 23845 50300 23857 50303
rect 23768 50288 23857 50300
rect 23477 50263 23535 50269
rect 23750 50236 23756 50288
rect 23808 50272 23857 50288
rect 23808 50236 23814 50272
rect 23845 50269 23857 50272
rect 23891 50269 23903 50303
rect 23845 50263 23903 50269
rect 24026 50260 24032 50312
rect 24084 50260 24090 50312
rect 24596 50309 24624 50340
rect 24581 50303 24639 50309
rect 24581 50269 24593 50303
rect 24627 50269 24639 50303
rect 24581 50263 24639 50269
rect 24670 50260 24676 50312
rect 24728 50300 24734 50312
rect 24805 50303 24863 50309
rect 24805 50300 24817 50303
rect 24728 50272 24817 50300
rect 24728 50260 24734 50272
rect 24805 50269 24817 50272
rect 24851 50269 24863 50303
rect 27982 50300 27988 50312
rect 27943 50272 27988 50300
rect 24805 50263 24863 50269
rect 27982 50260 27988 50272
rect 28040 50260 28046 50312
rect 24044 50232 24072 50260
rect 24949 50235 25007 50241
rect 23400 50204 23612 50232
rect 24044 50204 24716 50232
rect 22189 50195 22247 50201
rect 13173 50167 13231 50173
rect 13173 50164 13185 50167
rect 13136 50136 13185 50164
rect 13136 50124 13142 50136
rect 13173 50133 13185 50136
rect 13219 50133 13231 50167
rect 13173 50127 13231 50133
rect 14918 50124 14924 50176
rect 14976 50164 14982 50176
rect 16945 50167 17003 50173
rect 16945 50164 16957 50167
rect 14976 50136 16957 50164
rect 14976 50124 14982 50136
rect 16945 50133 16957 50136
rect 16991 50164 17003 50167
rect 21542 50164 21548 50176
rect 16991 50136 21548 50164
rect 16991 50133 17003 50136
rect 16945 50127 17003 50133
rect 21542 50124 21548 50136
rect 21600 50124 21606 50176
rect 22646 50124 22652 50176
rect 22704 50164 22710 50176
rect 23584 50173 23612 50204
rect 23385 50167 23443 50173
rect 23385 50164 23397 50167
rect 22704 50136 23397 50164
rect 22704 50124 22710 50136
rect 23385 50133 23397 50136
rect 23431 50133 23443 50167
rect 23385 50127 23443 50133
rect 23569 50167 23627 50173
rect 23569 50133 23581 50167
rect 23615 50133 23627 50167
rect 23569 50127 23627 50133
rect 23658 50124 23664 50176
rect 23716 50164 23722 50176
rect 24688 50173 24716 50204
rect 24949 50201 24961 50235
rect 24995 50232 25007 50235
rect 25222 50232 25228 50244
rect 24995 50204 25228 50232
rect 24995 50201 25007 50204
rect 24949 50195 25007 50201
rect 25222 50192 25228 50204
rect 25280 50192 25286 50244
rect 27890 50192 27896 50244
rect 27948 50232 27954 50244
rect 28534 50232 28540 50244
rect 27948 50204 28540 50232
rect 27948 50192 27954 50204
rect 28534 50192 28540 50204
rect 28592 50192 28598 50244
rect 28718 50192 28724 50244
rect 28776 50232 28782 50244
rect 28813 50235 28871 50241
rect 28813 50232 28825 50235
rect 28776 50204 28825 50232
rect 28776 50192 28782 50204
rect 28813 50201 28825 50204
rect 28859 50201 28871 50235
rect 28994 50232 29000 50244
rect 28955 50204 29000 50232
rect 28813 50195 28871 50201
rect 28994 50192 29000 50204
rect 29052 50192 29058 50244
rect 29730 50232 29736 50244
rect 29691 50204 29736 50232
rect 29730 50192 29736 50204
rect 29788 50192 29794 50244
rect 24673 50167 24731 50173
rect 23716 50136 23761 50164
rect 23716 50124 23722 50136
rect 24673 50133 24685 50167
rect 24719 50133 24731 50167
rect 24673 50127 24731 50133
rect 27246 50124 27252 50176
rect 27304 50164 27310 50176
rect 28169 50167 28227 50173
rect 28169 50164 28181 50167
rect 27304 50136 28181 50164
rect 27304 50124 27310 50136
rect 28169 50133 28181 50136
rect 28215 50133 28227 50167
rect 29822 50164 29828 50176
rect 29783 50136 29828 50164
rect 28169 50127 28227 50133
rect 29822 50124 29828 50136
rect 29880 50124 29886 50176
rect 1104 50074 30820 50096
rect 1104 50022 10880 50074
rect 10932 50022 10944 50074
rect 10996 50022 11008 50074
rect 11060 50022 11072 50074
rect 11124 50022 11136 50074
rect 11188 50022 20811 50074
rect 20863 50022 20875 50074
rect 20927 50022 20939 50074
rect 20991 50022 21003 50074
rect 21055 50022 21067 50074
rect 21119 50022 30820 50074
rect 1104 50000 30820 50022
rect 11882 49960 11888 49972
rect 11843 49932 11888 49960
rect 11882 49920 11888 49932
rect 11940 49920 11946 49972
rect 15654 49960 15660 49972
rect 15615 49932 15660 49960
rect 15654 49920 15660 49932
rect 15712 49920 15718 49972
rect 19978 49960 19984 49972
rect 19939 49932 19984 49960
rect 19978 49920 19984 49932
rect 20036 49920 20042 49972
rect 23014 49960 23020 49972
rect 22975 49932 23020 49960
rect 23014 49920 23020 49932
rect 23072 49920 23078 49972
rect 23750 49920 23756 49972
rect 23808 49960 23814 49972
rect 24213 49963 24271 49969
rect 23808 49932 23853 49960
rect 23808 49920 23814 49932
rect 24213 49929 24225 49963
rect 24259 49960 24271 49963
rect 24762 49960 24768 49972
rect 24259 49932 24768 49960
rect 24259 49929 24271 49932
rect 24213 49923 24271 49929
rect 24762 49920 24768 49932
rect 24820 49920 24826 49972
rect 24857 49963 24915 49969
rect 24857 49929 24869 49963
rect 24903 49929 24915 49963
rect 24857 49923 24915 49929
rect 25317 49963 25375 49969
rect 25317 49929 25329 49963
rect 25363 49960 25375 49963
rect 25774 49960 25780 49972
rect 25363 49932 25780 49960
rect 25363 49929 25375 49932
rect 25317 49923 25375 49929
rect 1486 49852 1492 49904
rect 1544 49892 1550 49904
rect 1581 49895 1639 49901
rect 1581 49892 1593 49895
rect 1544 49864 1593 49892
rect 1544 49852 1550 49864
rect 1581 49861 1593 49864
rect 1627 49861 1639 49895
rect 1762 49892 1768 49904
rect 1723 49864 1768 49892
rect 1581 49855 1639 49861
rect 1762 49852 1768 49864
rect 1820 49852 1826 49904
rect 24872 49892 24900 49923
rect 25222 49892 25228 49904
rect 23952 49864 24716 49892
rect 24872 49864 25228 49892
rect 2593 49827 2651 49833
rect 2593 49793 2605 49827
rect 2639 49824 2651 49827
rect 2774 49824 2780 49836
rect 2639 49796 2780 49824
rect 2639 49793 2651 49796
rect 2593 49787 2651 49793
rect 2774 49784 2780 49796
rect 2832 49784 2838 49836
rect 11698 49824 11704 49836
rect 11659 49796 11704 49824
rect 11698 49784 11704 49796
rect 11756 49784 11762 49836
rect 12989 49827 13047 49833
rect 12989 49793 13001 49827
rect 13035 49824 13047 49827
rect 14274 49824 14280 49836
rect 13035 49796 14280 49824
rect 13035 49793 13047 49796
rect 12989 49787 13047 49793
rect 14274 49784 14280 49796
rect 14332 49784 14338 49836
rect 15470 49824 15476 49836
rect 15431 49796 15476 49824
rect 15470 49784 15476 49796
rect 15528 49784 15534 49836
rect 19518 49784 19524 49836
rect 19576 49824 19582 49836
rect 19797 49827 19855 49833
rect 19797 49824 19809 49827
rect 19576 49796 19809 49824
rect 19576 49784 19582 49796
rect 19797 49793 19809 49796
rect 19843 49793 19855 49827
rect 19797 49787 19855 49793
rect 20346 49784 20352 49836
rect 20404 49824 20410 49836
rect 20441 49827 20499 49833
rect 20441 49824 20453 49827
rect 20404 49796 20453 49824
rect 20404 49784 20410 49796
rect 20441 49793 20453 49796
rect 20487 49793 20499 49827
rect 22370 49824 22376 49836
rect 22331 49796 22376 49824
rect 20441 49787 20499 49793
rect 22370 49784 22376 49796
rect 22428 49784 22434 49836
rect 1949 49759 2007 49765
rect 1949 49725 1961 49759
rect 1995 49756 2007 49759
rect 2498 49756 2504 49768
rect 1995 49728 2504 49756
rect 1995 49725 2007 49728
rect 1949 49719 2007 49725
rect 2498 49716 2504 49728
rect 2556 49716 2562 49768
rect 12526 49716 12532 49768
rect 12584 49756 12590 49768
rect 13265 49759 13323 49765
rect 13265 49756 13277 49759
rect 12584 49728 13277 49756
rect 12584 49716 12590 49728
rect 13265 49725 13277 49728
rect 13311 49725 13323 49759
rect 13265 49719 13323 49725
rect 14182 49716 14188 49768
rect 14240 49756 14246 49768
rect 14369 49759 14427 49765
rect 14369 49756 14381 49759
rect 14240 49728 14381 49756
rect 14240 49716 14246 49728
rect 14369 49725 14381 49728
rect 14415 49756 14427 49759
rect 14550 49756 14556 49768
rect 14415 49728 14556 49756
rect 14415 49725 14427 49728
rect 14369 49719 14427 49725
rect 14550 49716 14556 49728
rect 14608 49716 14614 49768
rect 17126 49716 17132 49768
rect 17184 49756 17190 49768
rect 17184 49728 23244 49756
rect 17184 49716 17190 49728
rect 14090 49648 14096 49700
rect 14148 49688 14154 49700
rect 22002 49688 22008 49700
rect 14148 49660 22008 49688
rect 14148 49648 14154 49660
rect 22002 49648 22008 49660
rect 22060 49648 22066 49700
rect 2130 49580 2136 49632
rect 2188 49620 2194 49632
rect 2409 49623 2467 49629
rect 2409 49620 2421 49623
rect 2188 49592 2421 49620
rect 2188 49580 2194 49592
rect 2409 49589 2421 49592
rect 2455 49589 2467 49623
rect 2409 49583 2467 49589
rect 20625 49623 20683 49629
rect 20625 49589 20637 49623
rect 20671 49620 20683 49623
rect 21542 49620 21548 49632
rect 20671 49592 21548 49620
rect 20671 49589 20683 49592
rect 20625 49583 20683 49589
rect 21542 49580 21548 49592
rect 21600 49580 21606 49632
rect 23216 49620 23244 49728
rect 23474 49716 23480 49768
rect 23532 49756 23538 49768
rect 23750 49756 23756 49768
rect 23532 49728 23756 49756
rect 23532 49716 23538 49728
rect 23750 49716 23756 49728
rect 23808 49756 23814 49768
rect 23952 49765 23980 49864
rect 24397 49827 24455 49833
rect 24397 49793 24409 49827
rect 24443 49824 24455 49827
rect 24578 49824 24584 49836
rect 24443 49796 24584 49824
rect 24443 49793 24455 49796
rect 24397 49787 24455 49793
rect 24578 49784 24584 49796
rect 24636 49784 24642 49836
rect 23937 49759 23995 49765
rect 23937 49756 23949 49759
rect 23808 49728 23949 49756
rect 23808 49716 23814 49728
rect 23937 49725 23949 49728
rect 23983 49725 23995 49759
rect 23937 49719 23995 49725
rect 24029 49759 24087 49765
rect 24029 49725 24041 49759
rect 24075 49725 24087 49759
rect 24029 49719 24087 49725
rect 24305 49759 24363 49765
rect 24305 49725 24317 49759
rect 24351 49756 24363 49759
rect 24486 49756 24492 49768
rect 24351 49728 24492 49756
rect 24351 49725 24363 49728
rect 24305 49719 24363 49725
rect 23290 49648 23296 49700
rect 23348 49688 23354 49700
rect 24044 49688 24072 49719
rect 24486 49716 24492 49728
rect 24544 49716 24550 49768
rect 24688 49756 24716 49864
rect 25222 49852 25228 49864
rect 25280 49852 25286 49904
rect 24762 49784 24768 49836
rect 24820 49824 24826 49836
rect 24820 49796 25176 49824
rect 24820 49784 24826 49796
rect 25148 49765 25176 49796
rect 25041 49759 25099 49765
rect 25041 49756 25053 49759
rect 24688 49728 25053 49756
rect 25041 49725 25053 49728
rect 25087 49725 25099 49759
rect 25041 49719 25099 49725
rect 25133 49759 25191 49765
rect 25133 49725 25145 49759
rect 25179 49725 25191 49759
rect 25133 49719 25191 49725
rect 24762 49688 24768 49700
rect 23348 49660 24768 49688
rect 23348 49648 23354 49660
rect 24762 49648 24768 49660
rect 24820 49648 24826 49700
rect 25332 49688 25360 49923
rect 25774 49920 25780 49932
rect 25832 49920 25838 49972
rect 30926 49960 30932 49972
rect 29748 49932 30932 49960
rect 28534 49852 28540 49904
rect 28592 49892 28598 49904
rect 28721 49895 28779 49901
rect 28721 49892 28733 49895
rect 28592 49864 28733 49892
rect 28592 49852 28598 49864
rect 28721 49861 28733 49864
rect 28767 49861 28779 49895
rect 28721 49855 28779 49861
rect 29086 49852 29092 49904
rect 29144 49892 29150 49904
rect 29748 49901 29776 49932
rect 30926 49920 30932 49932
rect 30984 49920 30990 49972
rect 29733 49895 29791 49901
rect 29733 49892 29745 49895
rect 29144 49864 29745 49892
rect 29144 49852 29150 49864
rect 29733 49861 29745 49864
rect 29779 49861 29791 49895
rect 29733 49855 29791 49861
rect 29822 49852 29828 49904
rect 29880 49892 29886 49904
rect 29917 49895 29975 49901
rect 29917 49892 29929 49895
rect 29880 49864 29929 49892
rect 29880 49852 29886 49864
rect 29917 49861 29929 49864
rect 29963 49861 29975 49895
rect 29917 49855 29975 49861
rect 25409 49827 25467 49833
rect 25409 49793 25421 49827
rect 25455 49824 25467 49827
rect 26326 49824 26332 49836
rect 25455 49796 26332 49824
rect 25455 49793 25467 49796
rect 25409 49787 25467 49793
rect 26326 49784 26332 49796
rect 26384 49784 26390 49836
rect 27246 49784 27252 49836
rect 27304 49824 27310 49836
rect 28813 49827 28871 49833
rect 27304 49796 28764 49824
rect 27304 49784 27310 49796
rect 25501 49759 25559 49765
rect 25501 49725 25513 49759
rect 25547 49725 25559 49759
rect 25501 49719 25559 49725
rect 24872 49660 25360 49688
rect 24872 49620 24900 49660
rect 23216 49592 24900 49620
rect 25222 49580 25228 49632
rect 25280 49620 25286 49632
rect 25516 49620 25544 49719
rect 25866 49716 25872 49768
rect 25924 49756 25930 49768
rect 28736 49765 28764 49796
rect 28813 49793 28825 49827
rect 28859 49824 28871 49827
rect 28994 49824 29000 49836
rect 28859 49796 29000 49824
rect 28859 49793 28871 49796
rect 28813 49787 28871 49793
rect 28994 49784 29000 49796
rect 29052 49824 29058 49836
rect 29052 49796 30052 49824
rect 29052 49784 29058 49796
rect 30024 49768 30052 49796
rect 28721 49759 28779 49765
rect 25924 49728 28396 49756
rect 25924 49716 25930 49728
rect 27430 49648 27436 49700
rect 27488 49688 27494 49700
rect 28261 49691 28319 49697
rect 28261 49688 28273 49691
rect 27488 49660 28273 49688
rect 27488 49648 27494 49660
rect 28261 49657 28273 49660
rect 28307 49657 28319 49691
rect 28368 49688 28396 49728
rect 28721 49725 28733 49759
rect 28767 49756 28779 49759
rect 29730 49756 29736 49768
rect 28767 49728 29736 49756
rect 28767 49725 28779 49728
rect 28721 49719 28779 49725
rect 29730 49716 29736 49728
rect 29788 49716 29794 49768
rect 30006 49756 30012 49768
rect 29967 49728 30012 49756
rect 30006 49716 30012 49728
rect 30064 49716 30070 49768
rect 29457 49691 29515 49697
rect 29457 49688 29469 49691
rect 28368 49660 29469 49688
rect 28261 49651 28319 49657
rect 29457 49657 29469 49660
rect 29503 49657 29515 49691
rect 29457 49651 29515 49657
rect 25280 49592 25544 49620
rect 25280 49580 25286 49592
rect 1104 49530 30820 49552
rect 1104 49478 5915 49530
rect 5967 49478 5979 49530
rect 6031 49478 6043 49530
rect 6095 49478 6107 49530
rect 6159 49478 6171 49530
rect 6223 49478 15846 49530
rect 15898 49478 15910 49530
rect 15962 49478 15974 49530
rect 16026 49478 16038 49530
rect 16090 49478 16102 49530
rect 16154 49478 25776 49530
rect 25828 49478 25840 49530
rect 25892 49478 25904 49530
rect 25956 49478 25968 49530
rect 26020 49478 26032 49530
rect 26084 49478 30820 49530
rect 1104 49456 30820 49478
rect 1949 49419 2007 49425
rect 1949 49385 1961 49419
rect 1995 49416 2007 49419
rect 1995 49388 10916 49416
rect 1995 49385 2007 49388
rect 1949 49379 2007 49385
rect 10888 49348 10916 49388
rect 10962 49376 10968 49428
rect 11020 49416 11026 49428
rect 14090 49416 14096 49428
rect 11020 49388 14096 49416
rect 11020 49376 11026 49388
rect 14090 49376 14096 49388
rect 14148 49376 14154 49428
rect 14274 49416 14280 49428
rect 14235 49388 14280 49416
rect 14274 49376 14280 49388
rect 14332 49376 14338 49428
rect 19613 49419 19671 49425
rect 19613 49385 19625 49419
rect 19659 49416 19671 49419
rect 19702 49416 19708 49428
rect 19659 49388 19708 49416
rect 19659 49385 19671 49388
rect 19613 49379 19671 49385
rect 19702 49376 19708 49388
rect 19760 49376 19766 49428
rect 21821 49419 21879 49425
rect 21821 49385 21833 49419
rect 21867 49416 21879 49419
rect 22370 49416 22376 49428
rect 21867 49388 22376 49416
rect 21867 49385 21879 49388
rect 21821 49379 21879 49385
rect 22370 49376 22376 49388
rect 22428 49376 22434 49428
rect 25409 49419 25467 49425
rect 25409 49385 25421 49419
rect 25455 49416 25467 49419
rect 25498 49416 25504 49428
rect 25455 49388 25504 49416
rect 25455 49385 25467 49388
rect 25409 49379 25467 49385
rect 25498 49376 25504 49388
rect 25556 49376 25562 49428
rect 26694 49416 26700 49428
rect 26655 49388 26700 49416
rect 26694 49376 26700 49388
rect 26752 49376 26758 49428
rect 27614 49416 27620 49428
rect 27575 49388 27620 49416
rect 27614 49376 27620 49388
rect 27672 49376 27678 49428
rect 17770 49348 17776 49360
rect 10888 49320 17776 49348
rect 17770 49308 17776 49320
rect 17828 49308 17834 49360
rect 20622 49308 20628 49360
rect 20680 49348 20686 49360
rect 23201 49351 23259 49357
rect 23201 49348 23213 49351
rect 20680 49320 23213 49348
rect 20680 49308 20686 49320
rect 23201 49317 23213 49320
rect 23247 49348 23259 49351
rect 23382 49348 23388 49360
rect 23247 49320 23388 49348
rect 23247 49317 23259 49320
rect 23201 49311 23259 49317
rect 23382 49308 23388 49320
rect 23440 49308 23446 49360
rect 25222 49308 25228 49360
rect 25280 49348 25286 49360
rect 25280 49320 26096 49348
rect 25280 49308 25286 49320
rect 2777 49283 2835 49289
rect 2777 49249 2789 49283
rect 2823 49280 2835 49283
rect 2823 49252 10088 49280
rect 2823 49249 2835 49252
rect 2777 49243 2835 49249
rect 1486 49172 1492 49224
rect 1544 49212 1550 49224
rect 1581 49215 1639 49221
rect 1581 49212 1593 49215
rect 1544 49184 1593 49212
rect 1544 49172 1550 49184
rect 1581 49181 1593 49184
rect 1627 49181 1639 49215
rect 1581 49175 1639 49181
rect 1670 49172 1676 49224
rect 1728 49212 1734 49224
rect 1765 49215 1823 49221
rect 1765 49212 1777 49215
rect 1728 49184 1777 49212
rect 1728 49172 1734 49184
rect 1765 49181 1777 49184
rect 1811 49181 1823 49215
rect 9950 49212 9956 49224
rect 9911 49184 9956 49212
rect 1765 49175 1823 49181
rect 9950 49172 9956 49184
rect 10008 49172 10014 49224
rect 10060 49212 10088 49252
rect 12066 49240 12072 49292
rect 12124 49280 12130 49292
rect 12437 49283 12495 49289
rect 12437 49280 12449 49283
rect 12124 49252 12449 49280
rect 12124 49240 12130 49252
rect 12437 49249 12449 49252
rect 12483 49280 12495 49283
rect 13357 49283 13415 49289
rect 13357 49280 13369 49283
rect 12483 49252 13369 49280
rect 12483 49249 12495 49252
rect 12437 49243 12495 49249
rect 13357 49249 13369 49252
rect 13403 49249 13415 49283
rect 13357 49243 13415 49249
rect 19794 49240 19800 49292
rect 19852 49280 19858 49292
rect 20073 49283 20131 49289
rect 20073 49280 20085 49283
rect 19852 49252 20085 49280
rect 19852 49240 19858 49252
rect 20073 49249 20085 49252
rect 20119 49280 20131 49283
rect 20993 49283 21051 49289
rect 20993 49280 21005 49283
rect 20119 49252 21005 49280
rect 20119 49249 20131 49252
rect 20073 49243 20131 49249
rect 20993 49249 21005 49252
rect 21039 49249 21051 49283
rect 20993 49243 21051 49249
rect 25593 49283 25651 49289
rect 25593 49249 25605 49283
rect 25639 49280 25651 49283
rect 25774 49280 25780 49292
rect 25639 49252 25780 49280
rect 25639 49249 25651 49252
rect 25593 49243 25651 49249
rect 25774 49240 25780 49252
rect 25832 49240 25838 49292
rect 26068 49289 26096 49320
rect 27154 49308 27160 49360
rect 27212 49308 27218 49360
rect 27430 49308 27436 49360
rect 27488 49348 27494 49360
rect 27488 49320 28286 49348
rect 27488 49308 27494 49320
rect 26053 49283 26111 49289
rect 26053 49249 26065 49283
rect 26099 49280 26111 49283
rect 26694 49280 26700 49292
rect 26099 49252 26700 49280
rect 26099 49249 26111 49252
rect 26053 49243 26111 49249
rect 26694 49240 26700 49252
rect 26752 49240 26758 49292
rect 27172 49280 27200 49308
rect 27172 49252 27844 49280
rect 12618 49212 12624 49224
rect 10060 49184 12624 49212
rect 12618 49172 12624 49184
rect 12676 49172 12682 49224
rect 14090 49212 14096 49224
rect 14051 49184 14096 49212
rect 14090 49172 14096 49184
rect 14148 49172 14154 49224
rect 21726 49172 21732 49224
rect 21784 49212 21790 49224
rect 22005 49215 22063 49221
rect 22005 49212 22017 49215
rect 21784 49184 22017 49212
rect 21784 49172 21790 49184
rect 22005 49181 22017 49184
rect 22051 49181 22063 49215
rect 22278 49212 22284 49224
rect 22239 49184 22284 49212
rect 22005 49175 22063 49181
rect 22278 49172 22284 49184
rect 22336 49172 22342 49224
rect 23017 49215 23075 49221
rect 23017 49181 23029 49215
rect 23063 49212 23075 49215
rect 23290 49212 23296 49224
rect 23063 49184 23296 49212
rect 23063 49181 23075 49184
rect 23017 49175 23075 49181
rect 23290 49172 23296 49184
rect 23348 49172 23354 49224
rect 25222 49172 25228 49224
rect 25280 49212 25286 49224
rect 25685 49215 25743 49221
rect 25685 49212 25697 49215
rect 25280 49184 25697 49212
rect 25280 49172 25286 49184
rect 25685 49181 25697 49184
rect 25731 49181 25743 49215
rect 25685 49175 25743 49181
rect 25866 49172 25872 49224
rect 25924 49212 25930 49224
rect 26418 49212 26424 49224
rect 25924 49184 26424 49212
rect 25924 49172 25930 49184
rect 26418 49172 26424 49184
rect 26476 49172 26482 49224
rect 26510 49172 26516 49224
rect 26568 49212 26574 49224
rect 26881 49215 26939 49221
rect 26881 49212 26893 49215
rect 26568 49184 26893 49212
rect 26568 49172 26574 49184
rect 26881 49181 26893 49184
rect 26927 49181 26939 49215
rect 26881 49175 26939 49181
rect 27157 49215 27215 49221
rect 27157 49181 27169 49215
rect 27203 49212 27215 49215
rect 27430 49212 27436 49224
rect 27203 49184 27436 49212
rect 27203 49181 27215 49184
rect 27157 49175 27215 49181
rect 27430 49172 27436 49184
rect 27488 49172 27494 49224
rect 27816 49221 27844 49252
rect 27890 49240 27896 49292
rect 27948 49280 27954 49292
rect 28166 49280 28172 49292
rect 27948 49252 28172 49280
rect 27948 49240 27954 49252
rect 28166 49240 28172 49252
rect 28224 49240 28230 49292
rect 27801 49215 27859 49221
rect 27801 49181 27813 49215
rect 27847 49181 27859 49215
rect 27801 49175 27859 49181
rect 28077 49215 28135 49221
rect 28077 49181 28089 49215
rect 28123 49212 28135 49215
rect 28258 49212 28286 49320
rect 28123 49184 28286 49212
rect 28629 49215 28687 49221
rect 28123 49181 28135 49184
rect 28077 49175 28135 49181
rect 28629 49181 28641 49215
rect 28675 49212 28687 49215
rect 28718 49212 28724 49224
rect 28675 49184 28724 49212
rect 28675 49181 28687 49184
rect 28629 49175 28687 49181
rect 28718 49172 28724 49184
rect 28776 49172 28782 49224
rect 2314 49104 2320 49156
rect 2372 49144 2378 49156
rect 2409 49147 2467 49153
rect 2409 49144 2421 49147
rect 2372 49116 2421 49144
rect 2372 49104 2378 49116
rect 2409 49113 2421 49116
rect 2455 49113 2467 49147
rect 2409 49107 2467 49113
rect 2593 49147 2651 49153
rect 2593 49113 2605 49147
rect 2639 49144 2651 49147
rect 3234 49144 3240 49156
rect 2639 49116 3240 49144
rect 2639 49113 2651 49116
rect 2593 49107 2651 49113
rect 3234 49104 3240 49116
rect 3292 49104 3298 49156
rect 9582 49104 9588 49156
rect 9640 49144 9646 49156
rect 10198 49147 10256 49153
rect 10198 49144 10210 49147
rect 9640 49116 10210 49144
rect 9640 49104 9646 49116
rect 10198 49113 10210 49116
rect 10244 49113 10256 49147
rect 10198 49107 10256 49113
rect 10962 49104 10968 49156
rect 11020 49104 11026 49156
rect 12342 49104 12348 49156
rect 12400 49144 12406 49156
rect 12529 49147 12587 49153
rect 12529 49144 12541 49147
rect 12400 49116 12541 49144
rect 12400 49104 12406 49116
rect 12529 49113 12541 49116
rect 12575 49113 12587 49147
rect 13170 49144 13176 49156
rect 13131 49116 13176 49144
rect 12529 49107 12587 49113
rect 13170 49104 13176 49116
rect 13228 49104 13234 49156
rect 20165 49147 20223 49153
rect 20165 49113 20177 49147
rect 20211 49144 20223 49147
rect 20346 49144 20352 49156
rect 20211 49116 20352 49144
rect 20211 49113 20223 49116
rect 20165 49107 20223 49113
rect 20346 49104 20352 49116
rect 20404 49104 20410 49156
rect 20809 49147 20867 49153
rect 20809 49113 20821 49147
rect 20855 49144 20867 49147
rect 21266 49144 21272 49156
rect 20855 49116 21272 49144
rect 20855 49113 20867 49116
rect 20809 49107 20867 49113
rect 21266 49104 21272 49116
rect 21324 49104 21330 49156
rect 22189 49147 22247 49153
rect 22189 49113 22201 49147
rect 22235 49144 22247 49147
rect 22462 49144 22468 49156
rect 22235 49116 22468 49144
rect 22235 49113 22247 49116
rect 22189 49107 22247 49113
rect 22462 49104 22468 49116
rect 22520 49104 22526 49156
rect 27065 49147 27123 49153
rect 27065 49144 27077 49147
rect 25792 49116 27077 49144
rect 9858 49036 9864 49088
rect 9916 49076 9922 49088
rect 10980 49076 11008 49104
rect 11333 49079 11391 49085
rect 11333 49076 11345 49079
rect 9916 49048 11345 49076
rect 9916 49036 9922 49048
rect 11333 49045 11345 49048
rect 11379 49045 11391 49079
rect 11333 49039 11391 49045
rect 11422 49036 11428 49088
rect 11480 49076 11486 49088
rect 11959 49079 12017 49085
rect 11959 49076 11971 49079
rect 11480 49048 11971 49076
rect 11480 49036 11486 49048
rect 11959 49045 11971 49048
rect 12005 49045 12017 49079
rect 11959 49039 12017 49045
rect 12158 49036 12164 49088
rect 12216 49076 12222 49088
rect 12437 49079 12495 49085
rect 12437 49076 12449 49079
rect 12216 49048 12449 49076
rect 12216 49036 12222 49048
rect 12437 49045 12449 49048
rect 12483 49045 12495 49079
rect 20070 49076 20076 49088
rect 20031 49048 20076 49076
rect 12437 49039 12495 49045
rect 20070 49036 20076 49048
rect 20128 49036 20134 49088
rect 20714 49036 20720 49088
rect 20772 49076 20778 49088
rect 22922 49076 22928 49088
rect 20772 49048 22928 49076
rect 20772 49036 20778 49048
rect 22922 49036 22928 49048
rect 22980 49036 22986 49088
rect 25498 49036 25504 49088
rect 25556 49076 25562 49088
rect 25792 49085 25820 49116
rect 27065 49113 27077 49116
rect 27111 49113 27123 49147
rect 27065 49107 27123 49113
rect 28166 49104 28172 49156
rect 28224 49144 28230 49156
rect 28350 49144 28356 49156
rect 28224 49116 28356 49144
rect 28224 49104 28230 49116
rect 28350 49104 28356 49116
rect 28408 49104 28414 49156
rect 29730 49144 29736 49156
rect 29691 49116 29736 49144
rect 29730 49104 29736 49116
rect 29788 49104 29794 49156
rect 30101 49147 30159 49153
rect 30101 49113 30113 49147
rect 30147 49144 30159 49147
rect 30926 49144 30932 49156
rect 30147 49116 30932 49144
rect 30147 49113 30159 49116
rect 30101 49107 30159 49113
rect 30926 49104 30932 49116
rect 30984 49104 30990 49156
rect 25777 49079 25835 49085
rect 25777 49076 25789 49079
rect 25556 49048 25789 49076
rect 25556 49036 25562 49048
rect 25777 49045 25789 49048
rect 25823 49045 25835 49079
rect 25777 49039 25835 49045
rect 25961 49079 26019 49085
rect 25961 49045 25973 49079
rect 26007 49076 26019 49079
rect 26418 49076 26424 49088
rect 26007 49048 26424 49076
rect 26007 49045 26019 49048
rect 25961 49039 26019 49045
rect 26418 49036 26424 49048
rect 26476 49036 26482 49088
rect 26970 49036 26976 49088
rect 27028 49076 27034 49088
rect 27522 49076 27528 49088
rect 27028 49048 27528 49076
rect 27028 49036 27034 49048
rect 27522 49036 27528 49048
rect 27580 49036 27586 49088
rect 27614 49036 27620 49088
rect 27672 49076 27678 49088
rect 27985 49079 28043 49085
rect 27985 49076 27997 49079
rect 27672 49048 27997 49076
rect 27672 49036 27678 49048
rect 27985 49045 27997 49048
rect 28031 49045 28043 49079
rect 27985 49039 28043 49045
rect 28905 49079 28963 49085
rect 28905 49045 28917 49079
rect 28951 49076 28963 49079
rect 28951 49048 30880 49076
rect 28951 49045 28963 49048
rect 28905 49039 28963 49045
rect 1104 48986 30820 49008
rect 1104 48934 10880 48986
rect 10932 48934 10944 48986
rect 10996 48934 11008 48986
rect 11060 48934 11072 48986
rect 11124 48934 11136 48986
rect 11188 48934 20811 48986
rect 20863 48934 20875 48986
rect 20927 48934 20939 48986
rect 20991 48934 21003 48986
rect 21055 48934 21067 48986
rect 21119 48934 30820 48986
rect 1104 48912 30820 48934
rect 3234 48872 3240 48884
rect 3195 48844 3240 48872
rect 3234 48832 3240 48844
rect 3292 48832 3298 48884
rect 9950 48832 9956 48884
rect 10008 48872 10014 48884
rect 10413 48875 10471 48881
rect 10413 48872 10425 48875
rect 10008 48844 10425 48872
rect 10008 48832 10014 48844
rect 10413 48841 10425 48844
rect 10459 48841 10471 48875
rect 13722 48872 13728 48884
rect 10413 48835 10471 48841
rect 10520 48844 13728 48872
rect 1486 48764 1492 48816
rect 1544 48804 1550 48816
rect 1581 48807 1639 48813
rect 1581 48804 1593 48807
rect 1544 48776 1593 48804
rect 1544 48764 1550 48776
rect 1581 48773 1593 48776
rect 1627 48773 1639 48807
rect 1581 48767 1639 48773
rect 1765 48807 1823 48813
rect 1765 48773 1777 48807
rect 1811 48804 1823 48807
rect 2130 48804 2136 48816
rect 1811 48776 2136 48804
rect 1811 48773 1823 48776
rect 1765 48767 1823 48773
rect 2130 48764 2136 48776
rect 2188 48764 2194 48816
rect 2777 48807 2835 48813
rect 2777 48773 2789 48807
rect 2823 48804 2835 48807
rect 10520 48804 10548 48844
rect 13722 48832 13728 48844
rect 13780 48832 13786 48884
rect 15194 48832 15200 48884
rect 15252 48872 15258 48884
rect 15252 48844 22784 48872
rect 15252 48832 15258 48844
rect 2823 48776 10548 48804
rect 2823 48773 2835 48776
rect 2777 48767 2835 48773
rect 11974 48764 11980 48816
rect 12032 48804 12038 48816
rect 12069 48807 12127 48813
rect 12069 48804 12081 48807
rect 12032 48776 12081 48804
rect 12032 48764 12038 48776
rect 12069 48773 12081 48776
rect 12115 48804 12127 48807
rect 12158 48804 12164 48816
rect 12115 48776 12164 48804
rect 12115 48773 12127 48776
rect 12069 48767 12127 48773
rect 12158 48764 12164 48776
rect 12216 48764 12222 48816
rect 18506 48804 18512 48816
rect 17411 48776 18512 48804
rect 2314 48696 2320 48748
rect 2372 48736 2378 48748
rect 2409 48739 2467 48745
rect 2409 48736 2421 48739
rect 2372 48708 2421 48736
rect 2372 48696 2378 48708
rect 2409 48705 2421 48708
rect 2455 48705 2467 48739
rect 2590 48736 2596 48748
rect 2551 48708 2596 48736
rect 2409 48699 2467 48705
rect 2590 48696 2596 48708
rect 2648 48696 2654 48748
rect 3418 48736 3424 48748
rect 3379 48708 3424 48736
rect 3418 48696 3424 48708
rect 3476 48696 3482 48748
rect 10229 48739 10287 48745
rect 10229 48705 10241 48739
rect 10275 48736 10287 48739
rect 11422 48736 11428 48748
rect 10275 48708 11428 48736
rect 10275 48705 10287 48708
rect 10229 48699 10287 48705
rect 11422 48696 11428 48708
rect 11480 48696 11486 48748
rect 14553 48739 14611 48745
rect 14553 48705 14565 48739
rect 14599 48736 14611 48739
rect 15746 48736 15752 48748
rect 14599 48708 15752 48736
rect 14599 48705 14611 48708
rect 14553 48699 14611 48705
rect 15746 48696 15752 48708
rect 15804 48696 15810 48748
rect 17411 48745 17439 48776
rect 18506 48764 18512 48776
rect 18564 48764 18570 48816
rect 19794 48804 19800 48816
rect 19755 48776 19800 48804
rect 19794 48764 19800 48776
rect 19852 48764 19858 48816
rect 19981 48807 20039 48813
rect 19981 48773 19993 48807
rect 20027 48804 20039 48807
rect 20162 48804 20168 48816
rect 20027 48776 20168 48804
rect 20027 48773 20039 48776
rect 19981 48767 20039 48773
rect 20162 48764 20168 48776
rect 20220 48764 20226 48816
rect 20714 48804 20720 48816
rect 20675 48776 20720 48804
rect 20714 48764 20720 48776
rect 20772 48764 20778 48816
rect 21542 48764 21548 48816
rect 21600 48804 21606 48816
rect 22370 48804 22376 48816
rect 21600 48776 22376 48804
rect 21600 48764 21606 48776
rect 22370 48764 22376 48776
rect 22428 48804 22434 48816
rect 22756 48804 22784 48844
rect 22922 48832 22928 48884
rect 22980 48872 22986 48884
rect 23569 48875 23627 48881
rect 23569 48872 23581 48875
rect 22980 48844 23581 48872
rect 22980 48832 22986 48844
rect 23569 48841 23581 48844
rect 23615 48841 23627 48875
rect 23569 48835 23627 48841
rect 24305 48875 24363 48881
rect 24305 48841 24317 48875
rect 24351 48872 24363 48875
rect 24486 48872 24492 48884
rect 24351 48844 24492 48872
rect 24351 48841 24363 48844
rect 24305 48835 24363 48841
rect 24486 48832 24492 48844
rect 24544 48832 24550 48884
rect 24578 48832 24584 48884
rect 24636 48872 24642 48884
rect 25133 48875 25191 48881
rect 25133 48872 25145 48875
rect 24636 48844 25145 48872
rect 24636 48832 24642 48844
rect 25133 48841 25145 48844
rect 25179 48841 25191 48875
rect 25682 48872 25688 48884
rect 25643 48844 25688 48872
rect 25133 48835 25191 48841
rect 25682 48832 25688 48844
rect 25740 48832 25746 48884
rect 25866 48832 25872 48884
rect 25924 48832 25930 48884
rect 25958 48832 25964 48884
rect 26016 48872 26022 48884
rect 26053 48875 26111 48881
rect 26053 48872 26065 48875
rect 26016 48844 26065 48872
rect 26016 48832 26022 48844
rect 26053 48841 26065 48844
rect 26099 48872 26111 48875
rect 26099 48844 26188 48872
rect 26099 48841 26111 48844
rect 26053 48835 26111 48841
rect 22428 48776 22692 48804
rect 22756 48776 24348 48804
rect 22428 48764 22434 48776
rect 17385 48739 17443 48745
rect 17385 48705 17397 48739
rect 17431 48705 17443 48739
rect 17494 48739 17552 48745
rect 17494 48736 17506 48739
rect 17385 48699 17443 48705
rect 17492 48705 17506 48736
rect 17540 48705 17552 48739
rect 17492 48699 17552 48705
rect 17589 48739 17647 48745
rect 17589 48705 17601 48739
rect 17635 48705 17647 48739
rect 17770 48736 17776 48748
rect 17731 48708 17776 48736
rect 17589 48699 17647 48705
rect 12066 48668 12072 48680
rect 12027 48640 12072 48668
rect 12066 48628 12072 48640
rect 12124 48628 12130 48680
rect 12158 48628 12164 48680
rect 12216 48668 12222 48680
rect 12342 48668 12348 48680
rect 12216 48640 12348 48668
rect 12216 48628 12222 48640
rect 12342 48628 12348 48640
rect 12400 48628 12406 48680
rect 11606 48600 11612 48612
rect 11567 48572 11612 48600
rect 11606 48560 11612 48572
rect 11664 48560 11670 48612
rect 14734 48600 14740 48612
rect 14695 48572 14740 48600
rect 14734 48560 14740 48572
rect 14792 48560 14798 48612
rect 17492 48600 17520 48699
rect 17604 48668 17632 48699
rect 17770 48696 17776 48708
rect 17828 48696 17834 48748
rect 22094 48696 22100 48748
rect 22152 48736 22158 48748
rect 22557 48739 22615 48745
rect 22557 48736 22569 48739
rect 22152 48708 22569 48736
rect 22152 48696 22158 48708
rect 22557 48705 22569 48708
rect 22603 48705 22615 48739
rect 22664 48736 22692 48776
rect 22833 48739 22891 48745
rect 22833 48736 22845 48739
rect 22664 48708 22845 48736
rect 22557 48699 22615 48705
rect 22833 48705 22845 48708
rect 22879 48705 22891 48739
rect 22833 48699 22891 48705
rect 23290 48696 23296 48748
rect 23348 48736 23354 48748
rect 23385 48739 23443 48745
rect 23385 48736 23397 48739
rect 23348 48708 23397 48736
rect 23348 48696 23354 48708
rect 23385 48705 23397 48708
rect 23431 48705 23443 48739
rect 23385 48699 23443 48705
rect 24213 48739 24271 48745
rect 24213 48705 24225 48739
rect 24259 48705 24271 48739
rect 24213 48699 24271 48705
rect 20073 48671 20131 48677
rect 17604 48640 17816 48668
rect 17788 48612 17816 48640
rect 20073 48637 20085 48671
rect 20119 48668 20131 48671
rect 20346 48668 20352 48680
rect 20119 48640 20352 48668
rect 20119 48637 20131 48640
rect 20073 48631 20131 48637
rect 20346 48628 20352 48640
rect 20404 48668 20410 48680
rect 23474 48668 23480 48680
rect 20404 48640 20668 48668
rect 20404 48628 20410 48640
rect 17586 48600 17592 48612
rect 17492 48572 17592 48600
rect 17586 48560 17592 48572
rect 17644 48560 17650 48612
rect 17770 48560 17776 48612
rect 17828 48560 17834 48612
rect 19518 48600 19524 48612
rect 19479 48572 19524 48600
rect 19518 48560 19524 48572
rect 19576 48560 19582 48612
rect 20640 48544 20668 48640
rect 22664 48640 23480 48668
rect 22664 48609 22692 48640
rect 23474 48628 23480 48640
rect 23532 48628 23538 48680
rect 22649 48603 22707 48609
rect 22649 48569 22661 48603
rect 22695 48569 22707 48603
rect 22649 48563 22707 48569
rect 22741 48603 22799 48609
rect 22741 48569 22753 48603
rect 22787 48569 22799 48603
rect 22741 48563 22799 48569
rect 1946 48532 1952 48544
rect 1907 48504 1952 48532
rect 1946 48492 1952 48504
rect 2004 48492 2010 48544
rect 17129 48535 17187 48541
rect 17129 48501 17141 48535
rect 17175 48532 17187 48535
rect 17402 48532 17408 48544
rect 17175 48504 17408 48532
rect 17175 48501 17187 48504
rect 17129 48495 17187 48501
rect 17402 48492 17408 48504
rect 17460 48492 17466 48544
rect 20622 48492 20628 48544
rect 20680 48532 20686 48544
rect 20809 48535 20867 48541
rect 20809 48532 20821 48535
rect 20680 48504 20821 48532
rect 20680 48492 20686 48504
rect 20809 48501 20821 48504
rect 20855 48501 20867 48535
rect 20809 48495 20867 48501
rect 22094 48492 22100 48544
rect 22152 48532 22158 48544
rect 22373 48535 22431 48541
rect 22373 48532 22385 48535
rect 22152 48504 22385 48532
rect 22152 48492 22158 48504
rect 22373 48501 22385 48504
rect 22419 48501 22431 48535
rect 22756 48532 22784 48563
rect 22922 48560 22928 48612
rect 22980 48600 22986 48612
rect 24228 48600 24256 48699
rect 22980 48572 24256 48600
rect 22980 48560 22986 48572
rect 23014 48532 23020 48544
rect 22756 48504 23020 48532
rect 22373 48495 22431 48501
rect 23014 48492 23020 48504
rect 23072 48492 23078 48544
rect 24320 48532 24348 48776
rect 25498 48764 25504 48816
rect 25556 48804 25562 48816
rect 25884 48804 25912 48832
rect 25556 48776 25912 48804
rect 26160 48804 26188 48844
rect 26970 48832 26976 48884
rect 27028 48872 27034 48884
rect 27157 48875 27215 48881
rect 27157 48872 27169 48875
rect 27028 48844 27169 48872
rect 27028 48832 27034 48844
rect 27157 48841 27169 48844
rect 27203 48841 27215 48875
rect 27157 48835 27215 48841
rect 27525 48875 27583 48881
rect 27525 48841 27537 48875
rect 27571 48841 27583 48875
rect 27525 48835 27583 48841
rect 27540 48804 27568 48835
rect 28258 48832 28264 48884
rect 28316 48872 28322 48884
rect 28629 48875 28687 48881
rect 28629 48872 28641 48875
rect 28316 48844 28641 48872
rect 28316 48832 28322 48844
rect 28629 48841 28641 48844
rect 28675 48872 28687 48875
rect 28994 48872 29000 48884
rect 28675 48844 29000 48872
rect 28675 48841 28687 48844
rect 28629 48835 28687 48841
rect 28994 48832 29000 48844
rect 29052 48832 29058 48884
rect 26160 48776 27568 48804
rect 25556 48764 25562 48776
rect 29546 48764 29552 48816
rect 29604 48804 29610 48816
rect 29917 48807 29975 48813
rect 29917 48804 29929 48807
rect 29604 48776 29929 48804
rect 29604 48764 29610 48776
rect 29917 48773 29929 48776
rect 29963 48773 29975 48807
rect 29917 48767 29975 48773
rect 24762 48696 24768 48748
rect 24820 48736 24826 48748
rect 25041 48739 25099 48745
rect 25041 48736 25053 48739
rect 24820 48708 25053 48736
rect 24820 48696 24826 48708
rect 25041 48705 25053 48708
rect 25087 48705 25099 48739
rect 25041 48699 25099 48705
rect 25222 48696 25228 48748
rect 25280 48736 25286 48748
rect 25961 48742 26019 48745
rect 25884 48739 26019 48742
rect 25884 48736 25973 48739
rect 25280 48714 25973 48736
rect 25280 48708 25912 48714
rect 25280 48696 25286 48708
rect 25961 48705 25973 48714
rect 26007 48705 26019 48739
rect 26418 48736 26424 48748
rect 25961 48699 26019 48705
rect 26252 48708 26424 48736
rect 25774 48628 25780 48680
rect 25832 48668 25838 48680
rect 25869 48671 25927 48677
rect 25869 48668 25881 48671
rect 25832 48640 25881 48668
rect 25832 48628 25838 48640
rect 25869 48637 25881 48640
rect 25915 48637 25927 48671
rect 25869 48631 25927 48637
rect 26142 48628 26148 48680
rect 26200 48668 26206 48680
rect 26252 48677 26280 48708
rect 26418 48696 26424 48708
rect 26476 48696 26482 48748
rect 26878 48696 26884 48748
rect 26936 48736 26942 48748
rect 27154 48736 27160 48748
rect 26936 48708 27160 48736
rect 26936 48696 26942 48708
rect 27154 48696 27160 48708
rect 27212 48736 27218 48748
rect 27341 48739 27399 48745
rect 27341 48736 27353 48739
rect 27212 48708 27353 48736
rect 27212 48696 27218 48708
rect 27341 48705 27353 48708
rect 27387 48705 27399 48739
rect 27341 48699 27399 48705
rect 27522 48696 27528 48748
rect 27580 48736 27586 48748
rect 27617 48739 27675 48745
rect 27617 48736 27629 48739
rect 27580 48708 27629 48736
rect 27580 48696 27586 48708
rect 27617 48705 27629 48708
rect 27663 48705 27675 48739
rect 27617 48699 27675 48705
rect 28258 48696 28264 48748
rect 28316 48736 28322 48748
rect 28537 48739 28595 48745
rect 28537 48736 28549 48739
rect 28316 48708 28549 48736
rect 28316 48696 28322 48708
rect 28537 48705 28549 48708
rect 28583 48705 28595 48739
rect 28537 48699 28595 48705
rect 29086 48696 29092 48748
rect 29144 48736 29150 48748
rect 29733 48739 29791 48745
rect 29733 48736 29745 48739
rect 29144 48708 29745 48736
rect 29144 48696 29150 48708
rect 29733 48705 29745 48708
rect 29779 48705 29791 48739
rect 29733 48699 29791 48705
rect 26237 48671 26295 48677
rect 26237 48668 26249 48671
rect 26200 48640 26249 48668
rect 26200 48628 26206 48640
rect 26237 48637 26249 48640
rect 26283 48637 26295 48671
rect 26237 48631 26295 48637
rect 26329 48671 26387 48677
rect 26329 48637 26341 48671
rect 26375 48668 26387 48671
rect 26694 48668 26700 48680
rect 26375 48640 26700 48668
rect 26375 48637 26387 48640
rect 26329 48631 26387 48637
rect 26694 48628 26700 48640
rect 26752 48628 26758 48680
rect 28813 48671 28871 48677
rect 28813 48637 28825 48671
rect 28859 48637 28871 48671
rect 30006 48668 30012 48680
rect 29967 48640 30012 48668
rect 28813 48631 28871 48637
rect 28828 48600 28856 48631
rect 30006 48628 30012 48640
rect 30064 48628 30070 48680
rect 30024 48600 30052 48628
rect 26114 48572 28396 48600
rect 28828 48572 30052 48600
rect 26114 48532 26142 48572
rect 24320 48504 26142 48532
rect 26510 48492 26516 48544
rect 26568 48532 26574 48544
rect 26878 48532 26884 48544
rect 26568 48504 26884 48532
rect 26568 48492 26574 48504
rect 26878 48492 26884 48504
rect 26936 48492 26942 48544
rect 28169 48535 28227 48541
rect 28169 48501 28181 48535
rect 28215 48532 28227 48535
rect 28258 48532 28264 48544
rect 28215 48504 28264 48532
rect 28215 48501 28227 48504
rect 28169 48495 28227 48501
rect 28258 48492 28264 48504
rect 28316 48492 28322 48544
rect 28368 48532 28396 48572
rect 29457 48535 29515 48541
rect 29457 48532 29469 48535
rect 28368 48504 29469 48532
rect 29457 48501 29469 48504
rect 29503 48501 29515 48535
rect 29457 48495 29515 48501
rect 1104 48442 30820 48464
rect 1104 48390 5915 48442
rect 5967 48390 5979 48442
rect 6031 48390 6043 48442
rect 6095 48390 6107 48442
rect 6159 48390 6171 48442
rect 6223 48390 15846 48442
rect 15898 48390 15910 48442
rect 15962 48390 15974 48442
rect 16026 48390 16038 48442
rect 16090 48390 16102 48442
rect 16154 48390 25776 48442
rect 25828 48390 25840 48442
rect 25892 48390 25904 48442
rect 25956 48390 25968 48442
rect 26020 48390 26032 48442
rect 26084 48390 30820 48442
rect 1104 48368 30820 48390
rect 1486 48288 1492 48340
rect 1544 48328 1550 48340
rect 1673 48331 1731 48337
rect 1673 48328 1685 48331
rect 1544 48300 1685 48328
rect 1544 48288 1550 48300
rect 1673 48297 1685 48300
rect 1719 48297 1731 48331
rect 1673 48291 1731 48297
rect 1946 48288 1952 48340
rect 2004 48328 2010 48340
rect 18506 48328 18512 48340
rect 2004 48300 12434 48328
rect 18467 48300 18512 48328
rect 2004 48288 2010 48300
rect 2685 48263 2743 48269
rect 2685 48229 2697 48263
rect 2731 48260 2743 48263
rect 2866 48260 2872 48272
rect 2731 48232 2872 48260
rect 2731 48229 2743 48232
rect 2685 48223 2743 48229
rect 2866 48220 2872 48232
rect 2924 48220 2930 48272
rect 11698 48220 11704 48272
rect 11756 48260 11762 48272
rect 11885 48263 11943 48269
rect 11885 48260 11897 48263
rect 11756 48232 11897 48260
rect 11756 48220 11762 48232
rect 11885 48229 11897 48232
rect 11931 48229 11943 48263
rect 11885 48223 11943 48229
rect 12406 48192 12434 48300
rect 18506 48288 18512 48300
rect 18564 48328 18570 48340
rect 18966 48328 18972 48340
rect 18564 48300 18972 48328
rect 18564 48288 18570 48300
rect 18966 48288 18972 48300
rect 19024 48288 19030 48340
rect 26234 48328 26240 48340
rect 26068 48300 26240 48328
rect 19518 48220 19524 48272
rect 19576 48260 19582 48272
rect 20533 48263 20591 48269
rect 20533 48260 20545 48263
rect 19576 48232 20545 48260
rect 19576 48220 19582 48232
rect 20533 48229 20545 48232
rect 20579 48229 20591 48263
rect 20533 48223 20591 48229
rect 21913 48263 21971 48269
rect 21913 48229 21925 48263
rect 21959 48260 21971 48263
rect 22462 48260 22468 48272
rect 21959 48232 22468 48260
rect 21959 48229 21971 48232
rect 21913 48223 21971 48229
rect 12406 48164 14964 48192
rect 1857 48127 1915 48133
rect 1857 48093 1869 48127
rect 1903 48124 1915 48127
rect 2406 48124 2412 48136
rect 1903 48096 2412 48124
rect 1903 48093 1915 48096
rect 1857 48087 1915 48093
rect 2406 48084 2412 48096
rect 2464 48084 2470 48136
rect 12066 48084 12072 48136
rect 12124 48124 12130 48136
rect 12161 48127 12219 48133
rect 12161 48124 12173 48127
rect 12124 48096 12173 48124
rect 12124 48084 12130 48096
rect 12161 48093 12173 48096
rect 12207 48093 12219 48127
rect 12161 48087 12219 48093
rect 14274 48084 14280 48136
rect 14332 48084 14338 48136
rect 14366 48084 14372 48136
rect 14424 48124 14430 48136
rect 14936 48133 14964 48164
rect 19426 48152 19432 48204
rect 19484 48192 19490 48204
rect 19794 48192 19800 48204
rect 19484 48164 19800 48192
rect 19484 48152 19490 48164
rect 19794 48152 19800 48164
rect 19852 48152 19858 48204
rect 20548 48192 20576 48223
rect 22462 48220 22468 48232
rect 22520 48220 22526 48272
rect 25314 48220 25320 48272
rect 25372 48260 25378 48272
rect 25685 48263 25743 48269
rect 25685 48260 25697 48263
rect 25372 48232 25697 48260
rect 25372 48220 25378 48232
rect 25685 48229 25697 48232
rect 25731 48229 25743 48263
rect 25685 48223 25743 48229
rect 26068 48192 26096 48300
rect 26234 48288 26240 48300
rect 26292 48288 26298 48340
rect 26418 48288 26424 48340
rect 26476 48288 26482 48340
rect 26510 48288 26516 48340
rect 26568 48288 26574 48340
rect 30852 48328 30880 49048
rect 30852 48300 31248 48328
rect 26142 48220 26148 48272
rect 26200 48260 26206 48272
rect 26436 48260 26464 48288
rect 26200 48232 26464 48260
rect 26200 48220 26206 48232
rect 26237 48195 26295 48201
rect 26237 48192 26249 48195
rect 20548 48164 23612 48192
rect 14553 48127 14611 48133
rect 14553 48124 14565 48127
rect 14424 48096 14565 48124
rect 14424 48084 14430 48096
rect 14553 48093 14565 48096
rect 14599 48093 14611 48127
rect 14553 48087 14611 48093
rect 14645 48127 14703 48133
rect 14645 48093 14657 48127
rect 14691 48093 14703 48127
rect 14645 48087 14703 48093
rect 14737 48127 14795 48133
rect 14737 48093 14749 48127
rect 14783 48093 14795 48127
rect 14737 48087 14795 48093
rect 14921 48127 14979 48133
rect 14921 48093 14933 48127
rect 14967 48093 14979 48127
rect 14921 48087 14979 48093
rect 17129 48127 17187 48133
rect 17129 48093 17141 48127
rect 17175 48124 17187 48127
rect 18506 48124 18512 48136
rect 17175 48096 18512 48124
rect 17175 48093 17187 48096
rect 17129 48087 17187 48093
rect 2314 48056 2320 48068
rect 2275 48028 2320 48056
rect 2314 48016 2320 48028
rect 2372 48016 2378 48068
rect 2501 48059 2559 48065
rect 2501 48025 2513 48059
rect 2547 48025 2559 48059
rect 12437 48059 12495 48065
rect 12437 48056 12449 48059
rect 2501 48019 2559 48025
rect 12176 48028 12449 48056
rect 1762 47948 1768 48000
rect 1820 47988 1826 48000
rect 2516 47988 2544 48019
rect 12176 48000 12204 48028
rect 12437 48025 12449 48028
rect 12483 48025 12495 48059
rect 13354 48056 13360 48068
rect 13315 48028 13360 48056
rect 12437 48019 12495 48025
rect 13354 48016 13360 48028
rect 13412 48016 13418 48068
rect 14292 48056 14320 48084
rect 14660 48056 14688 48087
rect 14292 48028 14688 48056
rect 14752 48056 14780 48087
rect 18506 48084 18512 48096
rect 18564 48084 18570 48136
rect 19242 48124 19248 48136
rect 19203 48096 19248 48124
rect 19242 48084 19248 48096
rect 19300 48084 19306 48136
rect 20346 48124 20352 48136
rect 20307 48096 20352 48124
rect 20346 48084 20352 48096
rect 20404 48084 20410 48136
rect 20714 48084 20720 48136
rect 20772 48124 20778 48136
rect 21177 48127 21235 48133
rect 21177 48124 21189 48127
rect 20772 48096 21189 48124
rect 20772 48084 20778 48096
rect 21177 48093 21189 48096
rect 21223 48093 21235 48127
rect 21177 48087 21235 48093
rect 21726 48084 21732 48136
rect 21784 48124 21790 48136
rect 21821 48127 21879 48133
rect 21821 48124 21833 48127
rect 21784 48096 21833 48124
rect 21784 48084 21790 48096
rect 21821 48093 21833 48096
rect 21867 48093 21879 48127
rect 21821 48087 21879 48093
rect 15102 48056 15108 48068
rect 14752 48028 15108 48056
rect 15102 48016 15108 48028
rect 15160 48016 15166 48068
rect 17402 48065 17408 48068
rect 16117 48059 16175 48065
rect 16117 48025 16129 48059
rect 16163 48056 16175 48059
rect 16163 48028 17356 48056
rect 16163 48025 16175 48028
rect 16117 48019 16175 48025
rect 1820 47960 2544 47988
rect 1820 47948 1826 47960
rect 12158 47948 12164 48000
rect 12216 47948 12222 48000
rect 12345 47991 12403 47997
rect 12345 47957 12357 47991
rect 12391 47988 12403 47991
rect 13449 47991 13507 47997
rect 13449 47988 13461 47991
rect 12391 47960 13461 47988
rect 12391 47957 12403 47960
rect 12345 47951 12403 47957
rect 13449 47957 13461 47960
rect 13495 47988 13507 47991
rect 13906 47988 13912 48000
rect 13495 47960 13912 47988
rect 13495 47957 13507 47960
rect 13449 47951 13507 47957
rect 13906 47948 13912 47960
rect 13964 47948 13970 48000
rect 14277 47991 14335 47997
rect 14277 47957 14289 47991
rect 14323 47988 14335 47991
rect 14918 47988 14924 48000
rect 14323 47960 14924 47988
rect 14323 47957 14335 47960
rect 14277 47951 14335 47957
rect 14918 47948 14924 47960
rect 14976 47948 14982 48000
rect 16206 47988 16212 48000
rect 16167 47960 16212 47988
rect 16206 47948 16212 47960
rect 16264 47948 16270 48000
rect 17328 47988 17356 48028
rect 17396 48019 17408 48065
rect 17460 48056 17466 48068
rect 21361 48059 21419 48065
rect 21361 48056 21373 48059
rect 17460 48028 17496 48056
rect 20364 48028 21373 48056
rect 17402 48016 17408 48019
rect 17460 48016 17466 48028
rect 20364 48000 20392 48028
rect 21361 48025 21373 48028
rect 21407 48025 21419 48059
rect 23584 48056 23612 48164
rect 25332 48164 26249 48192
rect 25332 48136 25360 48164
rect 26237 48161 26249 48164
rect 26283 48161 26295 48195
rect 26528 48192 26556 48288
rect 27065 48263 27123 48269
rect 27065 48229 27077 48263
rect 27111 48260 27123 48263
rect 27890 48260 27896 48272
rect 27111 48232 27896 48260
rect 27111 48229 27123 48232
rect 27065 48223 27123 48229
rect 27890 48220 27896 48232
rect 27948 48220 27954 48272
rect 28350 48220 28356 48272
rect 28408 48260 28414 48272
rect 28537 48263 28595 48269
rect 28537 48260 28549 48263
rect 28408 48232 28549 48260
rect 28408 48220 28414 48232
rect 28537 48229 28549 48232
rect 28583 48229 28595 48263
rect 28537 48223 28595 48229
rect 29549 48263 29607 48269
rect 29549 48229 29561 48263
rect 29595 48260 29607 48263
rect 31110 48260 31116 48272
rect 29595 48232 31116 48260
rect 29595 48229 29607 48232
rect 29549 48223 29607 48229
rect 31110 48220 31116 48232
rect 31168 48220 31174 48272
rect 26528 48164 27936 48192
rect 26237 48155 26295 48161
rect 25314 48084 25320 48136
rect 25372 48084 25378 48136
rect 25682 48084 25688 48136
rect 25740 48124 25746 48136
rect 25869 48127 25927 48133
rect 25869 48124 25881 48127
rect 25740 48096 25881 48124
rect 25740 48084 25746 48096
rect 25869 48093 25881 48096
rect 25915 48093 25927 48127
rect 25869 48087 25927 48093
rect 25961 48127 26019 48133
rect 25961 48093 25973 48127
rect 26007 48093 26019 48127
rect 25961 48087 26019 48093
rect 25222 48056 25228 48068
rect 23584 48028 25228 48056
rect 21361 48019 21419 48025
rect 25222 48016 25228 48028
rect 25280 48056 25286 48068
rect 25976 48056 26004 48087
rect 26050 48084 26056 48136
rect 26108 48133 26114 48136
rect 26108 48127 26157 48133
rect 26108 48093 26111 48127
rect 26145 48124 26157 48127
rect 26329 48127 26387 48133
rect 26145 48096 26201 48124
rect 26145 48093 26157 48096
rect 26108 48087 26157 48093
rect 26329 48093 26341 48127
rect 26375 48124 26387 48127
rect 26694 48124 26700 48136
rect 26375 48096 26700 48124
rect 26375 48093 26387 48096
rect 26329 48087 26387 48093
rect 26108 48084 26114 48087
rect 26694 48084 26700 48096
rect 26752 48084 26758 48136
rect 27264 48133 27292 48164
rect 27908 48136 27936 48164
rect 29012 48164 30052 48192
rect 29012 48136 29040 48164
rect 27249 48127 27307 48133
rect 27249 48093 27261 48127
rect 27295 48124 27307 48127
rect 27522 48124 27528 48136
rect 27295 48096 27329 48124
rect 27483 48096 27528 48124
rect 27295 48093 27307 48096
rect 27249 48087 27307 48093
rect 27522 48084 27528 48096
rect 27580 48084 27586 48136
rect 27890 48084 27896 48136
rect 27948 48124 27954 48136
rect 28721 48127 28779 48133
rect 28721 48124 28733 48127
rect 27948 48096 28733 48124
rect 27948 48084 27954 48096
rect 28721 48093 28733 48096
rect 28767 48093 28779 48127
rect 28994 48124 29000 48136
rect 28955 48096 29000 48124
rect 28721 48087 28779 48093
rect 25280 48028 26004 48056
rect 26068 48056 26096 48084
rect 27433 48059 27491 48065
rect 27433 48056 27445 48059
rect 26068 48028 27445 48056
rect 25280 48016 25286 48028
rect 27433 48025 27445 48028
rect 27479 48025 27491 48059
rect 28736 48056 28764 48087
rect 28994 48084 29000 48096
rect 29052 48084 29058 48136
rect 30024 48133 30052 48164
rect 29733 48127 29791 48133
rect 29733 48093 29745 48127
rect 29779 48093 29791 48127
rect 29733 48087 29791 48093
rect 30009 48127 30067 48133
rect 30009 48093 30021 48127
rect 30055 48093 30067 48127
rect 30009 48087 30067 48093
rect 29748 48056 29776 48087
rect 31110 48084 31116 48136
rect 31168 48124 31174 48136
rect 31220 48124 31248 48300
rect 31168 48096 31248 48124
rect 31168 48084 31174 48096
rect 28736 48028 29776 48056
rect 27433 48019 27491 48025
rect 18414 47988 18420 48000
rect 17328 47960 18420 47988
rect 18414 47948 18420 47960
rect 18472 47948 18478 48000
rect 19426 47988 19432 48000
rect 19387 47960 19432 47988
rect 19426 47948 19432 47960
rect 19484 47948 19490 48000
rect 20346 47948 20352 48000
rect 20404 47948 20410 48000
rect 20530 47948 20536 48000
rect 20588 47988 20594 48000
rect 28905 47991 28963 47997
rect 28905 47988 28917 47991
rect 20588 47960 28917 47988
rect 20588 47948 20594 47960
rect 28905 47957 28917 47960
rect 28951 47988 28963 47991
rect 28994 47988 29000 48000
rect 28951 47960 29000 47988
rect 28951 47957 28963 47960
rect 28905 47951 28963 47957
rect 28994 47948 29000 47960
rect 29052 47948 29058 48000
rect 29917 47991 29975 47997
rect 29917 47957 29929 47991
rect 29963 47988 29975 47991
rect 30282 47988 30288 48000
rect 29963 47960 30288 47988
rect 29963 47957 29975 47960
rect 29917 47951 29975 47957
rect 30282 47948 30288 47960
rect 30340 47948 30346 48000
rect 1104 47898 30820 47920
rect 1104 47846 10880 47898
rect 10932 47846 10944 47898
rect 10996 47846 11008 47898
rect 11060 47846 11072 47898
rect 11124 47846 11136 47898
rect 11188 47846 20811 47898
rect 20863 47846 20875 47898
rect 20927 47846 20939 47898
rect 20991 47846 21003 47898
rect 21055 47846 21067 47898
rect 21119 47846 30820 47898
rect 1104 47824 30820 47846
rect 1397 47787 1455 47793
rect 1397 47753 1409 47787
rect 1443 47784 1455 47787
rect 1762 47784 1768 47796
rect 1443 47756 1768 47784
rect 1443 47753 1455 47756
rect 1397 47747 1455 47753
rect 1762 47744 1768 47756
rect 1820 47744 1826 47796
rect 2041 47787 2099 47793
rect 2041 47753 2053 47787
rect 2087 47784 2099 47787
rect 2590 47784 2596 47796
rect 2087 47756 2596 47784
rect 2087 47753 2099 47756
rect 2041 47747 2099 47753
rect 2590 47744 2596 47756
rect 2648 47744 2654 47796
rect 13906 47784 13912 47796
rect 13867 47756 13912 47784
rect 13906 47744 13912 47756
rect 13964 47784 13970 47796
rect 15105 47787 15163 47793
rect 15105 47784 15117 47787
rect 13964 47756 15117 47784
rect 13964 47744 13970 47756
rect 15105 47753 15117 47756
rect 15151 47753 15163 47787
rect 15105 47747 15163 47753
rect 16025 47787 16083 47793
rect 16025 47753 16037 47787
rect 16071 47784 16083 47787
rect 17678 47784 17684 47796
rect 16071 47756 17684 47784
rect 16071 47753 16083 47756
rect 16025 47747 16083 47753
rect 17678 47744 17684 47756
rect 17736 47744 17742 47796
rect 17862 47744 17868 47796
rect 17920 47784 17926 47796
rect 18506 47784 18512 47796
rect 17920 47756 18184 47784
rect 18467 47756 18512 47784
rect 17920 47744 17926 47756
rect 2498 47676 2504 47728
rect 2556 47716 2562 47728
rect 2556 47688 2774 47716
rect 2556 47676 2562 47688
rect 1578 47648 1584 47660
rect 1539 47620 1584 47648
rect 1578 47608 1584 47620
rect 1636 47608 1642 47660
rect 2222 47648 2228 47660
rect 2183 47620 2228 47648
rect 2222 47608 2228 47620
rect 2280 47608 2286 47660
rect 2746 47444 2774 47688
rect 14734 47676 14740 47728
rect 14792 47716 14798 47728
rect 14921 47719 14979 47725
rect 14921 47716 14933 47719
rect 14792 47688 14933 47716
rect 14792 47676 14798 47688
rect 14921 47685 14933 47688
rect 14967 47685 14979 47719
rect 18156 47716 18184 47756
rect 18506 47744 18512 47756
rect 18564 47744 18570 47796
rect 25958 47784 25964 47796
rect 25919 47756 25964 47784
rect 25958 47744 25964 47756
rect 26016 47744 26022 47796
rect 26050 47716 26056 47728
rect 18156 47688 26056 47716
rect 14921 47679 14979 47685
rect 26050 47676 26056 47688
rect 26108 47676 26114 47728
rect 28994 47676 29000 47728
rect 29052 47716 29058 47728
rect 29917 47719 29975 47725
rect 29917 47716 29929 47719
rect 29052 47688 29929 47716
rect 29052 47676 29058 47688
rect 29917 47685 29929 47688
rect 29963 47685 29975 47719
rect 29917 47679 29975 47685
rect 30006 47676 30012 47728
rect 30064 47716 30070 47728
rect 30064 47688 30109 47716
rect 30064 47676 30070 47688
rect 14458 47648 14464 47660
rect 13924 47620 14464 47648
rect 13924 47589 13952 47620
rect 14458 47608 14464 47620
rect 14516 47648 14522 47660
rect 14752 47648 14780 47676
rect 14516 47620 14780 47648
rect 15933 47651 15991 47657
rect 14516 47608 14522 47620
rect 15933 47617 15945 47651
rect 15979 47648 15991 47651
rect 16758 47648 16764 47660
rect 15979 47620 16764 47648
rect 15979 47617 15991 47620
rect 15933 47611 15991 47617
rect 16758 47608 16764 47620
rect 16816 47608 16822 47660
rect 17310 47648 17316 47660
rect 17236 47620 17316 47648
rect 13909 47583 13967 47589
rect 13909 47549 13921 47583
rect 13955 47549 13967 47583
rect 13909 47543 13967 47549
rect 14001 47583 14059 47589
rect 14001 47549 14013 47583
rect 14047 47580 14059 47583
rect 14550 47580 14556 47592
rect 14047 47552 14556 47580
rect 14047 47549 14059 47552
rect 14001 47543 14059 47549
rect 14550 47540 14556 47552
rect 14608 47580 14614 47592
rect 17236 47589 17264 47620
rect 17310 47608 17316 47620
rect 17368 47608 17374 47660
rect 17474 47608 17480 47660
rect 17532 47657 17538 47660
rect 17702 47657 17760 47663
rect 17532 47651 17555 47657
rect 17543 47617 17555 47651
rect 17589 47651 17647 47657
rect 17589 47632 17601 47651
rect 17532 47611 17555 47617
rect 17585 47617 17601 47632
rect 17635 47617 17647 47651
rect 17702 47623 17714 47657
rect 17748 47654 17760 47657
rect 17748 47626 17816 47654
rect 17748 47623 17760 47626
rect 17702 47617 17760 47623
rect 17585 47611 17647 47617
rect 17532 47608 17538 47611
rect 17585 47604 17623 47611
rect 15197 47583 15255 47589
rect 15197 47580 15209 47583
rect 14608 47552 15209 47580
rect 14608 47540 14614 47552
rect 15197 47549 15209 47552
rect 15243 47549 15255 47583
rect 15197 47543 15255 47549
rect 17221 47583 17279 47589
rect 17221 47549 17233 47583
rect 17267 47549 17279 47583
rect 17221 47543 17279 47549
rect 17585 47524 17613 47604
rect 17788 47580 17816 47626
rect 17865 47651 17923 47657
rect 17865 47617 17877 47651
rect 17911 47617 17923 47651
rect 18322 47648 18328 47660
rect 18283 47620 18328 47648
rect 17865 47611 17923 47617
rect 17696 47552 17816 47580
rect 17696 47524 17724 47552
rect 13449 47515 13507 47521
rect 13449 47481 13461 47515
rect 13495 47512 13507 47515
rect 14090 47512 14096 47524
rect 13495 47484 14096 47512
rect 13495 47481 13507 47484
rect 13449 47475 13507 47481
rect 14090 47472 14096 47484
rect 14148 47472 14154 47524
rect 14642 47512 14648 47524
rect 14603 47484 14648 47512
rect 14642 47472 14648 47484
rect 14700 47472 14706 47524
rect 17585 47484 17592 47524
rect 17586 47472 17592 47484
rect 17644 47472 17650 47524
rect 17678 47472 17684 47524
rect 17736 47472 17742 47524
rect 17880 47444 17908 47611
rect 18322 47608 18328 47620
rect 18380 47608 18386 47660
rect 18969 47651 19027 47657
rect 18969 47617 18981 47651
rect 19015 47617 19027 47651
rect 18969 47611 19027 47617
rect 17954 47540 17960 47592
rect 18012 47580 18018 47592
rect 18984 47580 19012 47611
rect 19978 47608 19984 47660
rect 20036 47648 20042 47660
rect 20257 47651 20315 47657
rect 20257 47648 20269 47651
rect 20036 47620 20269 47648
rect 20036 47608 20042 47620
rect 20257 47617 20269 47620
rect 20303 47617 20315 47651
rect 26142 47648 26148 47660
rect 26103 47620 26148 47648
rect 20257 47611 20315 47617
rect 26142 47608 26148 47620
rect 26200 47608 26206 47660
rect 26329 47651 26387 47657
rect 26329 47617 26341 47651
rect 26375 47617 26387 47651
rect 26329 47611 26387 47617
rect 26421 47651 26479 47657
rect 26421 47617 26433 47651
rect 26467 47648 26479 47651
rect 26467 47620 27568 47648
rect 26467 47617 26479 47620
rect 26421 47611 26479 47617
rect 18012 47552 19012 47580
rect 18012 47540 18018 47552
rect 25222 47540 25228 47592
rect 25280 47580 25286 47592
rect 26344 47580 26372 47611
rect 27540 47592 27568 47620
rect 25280 47552 26372 47580
rect 25280 47540 25286 47552
rect 27246 47540 27252 47592
rect 27304 47580 27310 47592
rect 27433 47583 27491 47589
rect 27433 47580 27445 47583
rect 27304 47552 27445 47580
rect 27304 47540 27310 47552
rect 27433 47549 27445 47552
rect 27479 47549 27491 47583
rect 27433 47543 27491 47549
rect 27522 47540 27528 47592
rect 27580 47580 27586 47592
rect 27709 47583 27767 47589
rect 27709 47580 27721 47583
rect 27580 47552 27721 47580
rect 27580 47540 27586 47552
rect 27709 47549 27721 47552
rect 27755 47549 27767 47583
rect 29825 47583 29883 47589
rect 29825 47580 29837 47583
rect 27709 47543 27767 47549
rect 29564 47552 29837 47580
rect 19794 47472 19800 47524
rect 19852 47512 19858 47524
rect 29457 47515 29515 47521
rect 29457 47512 29469 47515
rect 19852 47484 29469 47512
rect 19852 47472 19858 47484
rect 29457 47481 29469 47484
rect 29503 47481 29515 47515
rect 29457 47475 29515 47481
rect 19150 47444 19156 47456
rect 2746 47416 17908 47444
rect 19111 47416 19156 47444
rect 19150 47404 19156 47416
rect 19208 47404 19214 47456
rect 20441 47447 20499 47453
rect 20441 47413 20453 47447
rect 20487 47444 20499 47447
rect 20714 47444 20720 47456
rect 20487 47416 20720 47444
rect 20487 47413 20499 47416
rect 20441 47407 20499 47413
rect 20714 47404 20720 47416
rect 20772 47404 20778 47456
rect 25498 47404 25504 47456
rect 25556 47444 25562 47456
rect 26418 47444 26424 47456
rect 25556 47416 26424 47444
rect 25556 47404 25562 47416
rect 26418 47404 26424 47416
rect 26476 47404 26482 47456
rect 28350 47404 28356 47456
rect 28408 47444 28414 47456
rect 29564 47444 29592 47552
rect 29825 47549 29837 47552
rect 29871 47549 29883 47583
rect 29825 47543 29883 47549
rect 28408 47416 29592 47444
rect 28408 47404 28414 47416
rect 1104 47354 30820 47376
rect 1104 47302 5915 47354
rect 5967 47302 5979 47354
rect 6031 47302 6043 47354
rect 6095 47302 6107 47354
rect 6159 47302 6171 47354
rect 6223 47302 15846 47354
rect 15898 47302 15910 47354
rect 15962 47302 15974 47354
rect 16026 47302 16038 47354
rect 16090 47302 16102 47354
rect 16154 47302 25776 47354
rect 25828 47302 25840 47354
rect 25892 47302 25904 47354
rect 25956 47302 25968 47354
rect 26020 47302 26032 47354
rect 26084 47302 30820 47354
rect 1104 47280 30820 47302
rect 14366 47200 14372 47252
rect 14424 47240 14430 47252
rect 14424 47212 16068 47240
rect 14424 47200 14430 47212
rect 1578 47036 1584 47048
rect 1539 47008 1584 47036
rect 1578 46996 1584 47008
rect 1636 46996 1642 47048
rect 2406 46996 2412 47048
rect 2464 47036 2470 47048
rect 2593 47039 2651 47045
rect 2593 47036 2605 47039
rect 2464 47008 2605 47036
rect 2464 46996 2470 47008
rect 2593 47005 2605 47008
rect 2639 47005 2651 47039
rect 2593 46999 2651 47005
rect 13357 47039 13415 47045
rect 13357 47005 13369 47039
rect 13403 47036 13415 47039
rect 14366 47036 14372 47048
rect 13403 47008 14372 47036
rect 13403 47005 13415 47008
rect 13357 46999 13415 47005
rect 14366 46996 14372 47008
rect 14424 46996 14430 47048
rect 14642 47036 14648 47048
rect 14603 47008 14648 47036
rect 14642 46996 14648 47008
rect 14700 46996 14706 47048
rect 14918 47045 14924 47048
rect 14912 47036 14924 47045
rect 14879 47008 14924 47036
rect 14912 46999 14924 47008
rect 14918 46996 14924 46999
rect 14976 46996 14982 47048
rect 13541 46971 13599 46977
rect 13541 46937 13553 46971
rect 13587 46968 13599 46971
rect 14734 46968 14740 46980
rect 13587 46940 14740 46968
rect 13587 46937 13599 46940
rect 13541 46931 13599 46937
rect 14734 46928 14740 46940
rect 14792 46928 14798 46980
rect 16040 46968 16068 47212
rect 17494 47200 17500 47252
rect 17552 47240 17558 47252
rect 18693 47243 18751 47249
rect 18693 47240 18705 47243
rect 17552 47212 18705 47240
rect 17552 47200 17558 47212
rect 18693 47209 18705 47212
rect 18739 47240 18751 47243
rect 20530 47240 20536 47252
rect 18739 47212 20536 47240
rect 18739 47209 18751 47212
rect 18693 47203 18751 47209
rect 20530 47200 20536 47212
rect 20588 47200 20594 47252
rect 23474 47240 23480 47252
rect 23435 47212 23480 47240
rect 23474 47200 23480 47212
rect 23532 47200 23538 47252
rect 24026 47200 24032 47252
rect 24084 47240 24090 47252
rect 24949 47243 25007 47249
rect 24949 47240 24961 47243
rect 24084 47212 24961 47240
rect 24084 47200 24090 47212
rect 24949 47209 24961 47212
rect 24995 47209 25007 47243
rect 24949 47203 25007 47209
rect 26513 47243 26571 47249
rect 26513 47209 26525 47243
rect 26559 47240 26571 47243
rect 26602 47240 26608 47252
rect 26559 47212 26608 47240
rect 26559 47209 26571 47212
rect 26513 47203 26571 47209
rect 26602 47200 26608 47212
rect 26660 47200 26666 47252
rect 16853 47175 16911 47181
rect 16853 47141 16865 47175
rect 16899 47172 16911 47175
rect 17034 47172 17040 47184
rect 16899 47144 17040 47172
rect 16899 47141 16911 47144
rect 16853 47135 16911 47141
rect 17034 47132 17040 47144
rect 17092 47132 17098 47184
rect 19242 47132 19248 47184
rect 19300 47132 19306 47184
rect 19429 47175 19487 47181
rect 19429 47141 19441 47175
rect 19475 47172 19487 47175
rect 19610 47172 19616 47184
rect 19475 47144 19616 47172
rect 19475 47141 19487 47144
rect 19429 47135 19487 47141
rect 19610 47132 19616 47144
rect 19668 47132 19674 47184
rect 22554 47132 22560 47184
rect 22612 47172 22618 47184
rect 22925 47175 22983 47181
rect 22925 47172 22937 47175
rect 22612 47144 22937 47172
rect 22612 47132 22618 47144
rect 22925 47141 22937 47144
rect 22971 47141 22983 47175
rect 22925 47135 22983 47141
rect 24762 47132 24768 47184
rect 24820 47172 24826 47184
rect 26050 47172 26056 47184
rect 24820 47144 26056 47172
rect 24820 47132 24826 47144
rect 26050 47132 26056 47144
rect 26108 47132 26114 47184
rect 27246 47172 27252 47184
rect 26620 47144 27252 47172
rect 17310 47104 17316 47116
rect 17271 47076 17316 47104
rect 17310 47064 17316 47076
rect 17368 47064 17374 47116
rect 19260 47104 19288 47132
rect 22572 47104 22600 47132
rect 26620 47116 26648 47144
rect 27246 47132 27252 47144
rect 27304 47132 27310 47184
rect 19260 47076 19932 47104
rect 16669 47039 16727 47045
rect 16669 47005 16681 47039
rect 16715 47036 16727 47039
rect 18138 47036 18144 47048
rect 16715 47008 18144 47036
rect 16715 47005 16727 47008
rect 16669 46999 16727 47005
rect 18138 46996 18144 47008
rect 18196 46996 18202 47048
rect 19245 47039 19303 47045
rect 19245 47005 19257 47039
rect 19291 47036 19303 47039
rect 19334 47036 19340 47048
rect 19291 47008 19340 47036
rect 19291 47005 19303 47008
rect 19245 46999 19303 47005
rect 19334 46996 19340 47008
rect 19392 46996 19398 47048
rect 19904 47045 19932 47076
rect 22296 47076 22600 47104
rect 22296 47048 22324 47076
rect 26142 47064 26148 47116
rect 26200 47064 26206 47116
rect 26602 47064 26608 47116
rect 26660 47064 26666 47116
rect 27154 47064 27160 47116
rect 27212 47104 27218 47116
rect 27433 47107 27491 47113
rect 27433 47104 27445 47107
rect 27212 47076 27445 47104
rect 27212 47064 27218 47076
rect 27433 47073 27445 47076
rect 27479 47073 27491 47107
rect 27433 47067 27491 47073
rect 27709 47107 27767 47113
rect 27709 47073 27721 47107
rect 27755 47104 27767 47107
rect 27890 47104 27896 47116
rect 27755 47076 27896 47104
rect 27755 47073 27767 47076
rect 27709 47067 27767 47073
rect 27890 47064 27896 47076
rect 27948 47064 27954 47116
rect 30742 47064 30748 47116
rect 30800 47104 30806 47116
rect 30926 47104 30932 47116
rect 30800 47076 30932 47104
rect 30800 47064 30806 47076
rect 30926 47064 30932 47076
rect 30984 47064 30990 47116
rect 19889 47039 19947 47045
rect 19889 47005 19901 47039
rect 19935 47005 19947 47039
rect 22278 47036 22284 47048
rect 19889 46999 19947 47005
rect 19996 47008 22094 47036
rect 22191 47008 22284 47036
rect 16040 46940 17172 46968
rect 1397 46903 1455 46909
rect 1397 46869 1409 46903
rect 1443 46900 1455 46903
rect 2222 46900 2228 46912
rect 1443 46872 2228 46900
rect 1443 46869 1455 46872
rect 1397 46863 1455 46869
rect 2222 46860 2228 46872
rect 2280 46860 2286 46912
rect 2314 46860 2320 46912
rect 2372 46900 2378 46912
rect 16040 46909 16068 46940
rect 2409 46903 2467 46909
rect 2409 46900 2421 46903
rect 2372 46872 2421 46900
rect 2372 46860 2378 46872
rect 2409 46869 2421 46872
rect 2455 46869 2467 46903
rect 2409 46863 2467 46869
rect 16025 46903 16083 46909
rect 16025 46869 16037 46903
rect 16071 46869 16083 46903
rect 17144 46900 17172 46940
rect 17218 46928 17224 46980
rect 17276 46968 17282 46980
rect 17558 46971 17616 46977
rect 17558 46968 17570 46971
rect 17276 46940 17570 46968
rect 17276 46928 17282 46940
rect 17558 46937 17570 46940
rect 17604 46937 17616 46971
rect 19996 46968 20024 47008
rect 17558 46931 17616 46937
rect 17696 46940 20024 46968
rect 17696 46900 17724 46940
rect 20530 46928 20536 46980
rect 20588 46968 20594 46980
rect 20625 46971 20683 46977
rect 20625 46968 20637 46971
rect 20588 46940 20637 46968
rect 20588 46928 20594 46940
rect 20625 46937 20637 46940
rect 20671 46937 20683 46971
rect 20625 46931 20683 46937
rect 20809 46971 20867 46977
rect 20809 46937 20821 46971
rect 20855 46968 20867 46971
rect 21174 46968 21180 46980
rect 20855 46940 21180 46968
rect 20855 46937 20867 46940
rect 20809 46931 20867 46937
rect 21174 46928 21180 46940
rect 21232 46928 21238 46980
rect 22066 46968 22094 47008
rect 22278 46996 22284 47008
rect 22336 46996 22342 47048
rect 22465 47039 22523 47045
rect 22465 47005 22477 47039
rect 22511 47036 22523 47039
rect 22554 47036 22560 47048
rect 22511 47008 22560 47036
rect 22511 47005 22523 47008
rect 22465 46999 22523 47005
rect 22554 46996 22560 47008
rect 22612 47036 22618 47048
rect 22738 47036 22744 47048
rect 22612 47008 22744 47036
rect 22612 46996 22618 47008
rect 22738 46996 22744 47008
rect 22796 46996 22802 47048
rect 23106 46996 23112 47048
rect 23164 47036 23170 47048
rect 23201 47039 23259 47045
rect 23201 47036 23213 47039
rect 23164 47008 23213 47036
rect 23164 46996 23170 47008
rect 23201 47005 23213 47008
rect 23247 47005 23259 47039
rect 26160 47036 26188 47064
rect 26697 47039 26755 47045
rect 26697 47036 26709 47039
rect 26160 47008 26709 47036
rect 23201 46999 23259 47005
rect 26697 47005 26709 47008
rect 26743 47005 26755 47039
rect 26697 46999 26755 47005
rect 26973 47039 27031 47045
rect 26973 47005 26985 47039
rect 27019 47036 27031 47039
rect 27522 47036 27528 47048
rect 27019 47008 27528 47036
rect 27019 47005 27031 47008
rect 26973 46999 27031 47005
rect 27522 46996 27528 47008
rect 27580 46996 27586 47048
rect 28718 47036 28724 47048
rect 28679 47008 28724 47036
rect 28718 46996 28724 47008
rect 28776 46996 28782 47048
rect 22066 46940 24716 46968
rect 20070 46900 20076 46912
rect 17144 46872 17724 46900
rect 20031 46872 20076 46900
rect 16025 46863 16083 46869
rect 20070 46860 20076 46872
rect 20128 46860 20134 46912
rect 22370 46900 22376 46912
rect 22331 46872 22376 46900
rect 22370 46860 22376 46872
rect 22428 46860 22434 46912
rect 23014 46860 23020 46912
rect 23072 46900 23078 46912
rect 23109 46903 23167 46909
rect 23109 46900 23121 46903
rect 23072 46872 23121 46900
rect 23072 46860 23078 46872
rect 23109 46869 23121 46872
rect 23155 46869 23167 46903
rect 23109 46863 23167 46869
rect 23293 46903 23351 46909
rect 23293 46869 23305 46903
rect 23339 46900 23351 46903
rect 23382 46900 23388 46912
rect 23339 46872 23388 46900
rect 23339 46869 23351 46872
rect 23293 46863 23351 46869
rect 23382 46860 23388 46872
rect 23440 46860 23446 46912
rect 24688 46900 24716 46940
rect 24762 46928 24768 46980
rect 24820 46968 24826 46980
rect 24857 46971 24915 46977
rect 24857 46968 24869 46971
rect 24820 46940 24869 46968
rect 24820 46928 24826 46940
rect 24857 46937 24869 46940
rect 24903 46937 24915 46971
rect 24857 46931 24915 46937
rect 26142 46928 26148 46980
rect 26200 46968 26206 46980
rect 26881 46971 26939 46977
rect 26881 46968 26893 46971
rect 26200 46940 26893 46968
rect 26200 46928 26206 46940
rect 26881 46937 26893 46940
rect 26927 46937 26939 46971
rect 29730 46968 29736 46980
rect 29691 46940 29736 46968
rect 26881 46931 26939 46937
rect 29730 46928 29736 46940
rect 29788 46928 29794 46980
rect 30101 46971 30159 46977
rect 30101 46937 30113 46971
rect 30147 46968 30159 46971
rect 30742 46968 30748 46980
rect 30147 46940 30748 46968
rect 30147 46937 30159 46940
rect 30101 46931 30159 46937
rect 30742 46928 30748 46940
rect 30800 46928 30806 46980
rect 26510 46900 26516 46912
rect 24688 46872 26516 46900
rect 26510 46860 26516 46872
rect 26568 46860 26574 46912
rect 27522 46860 27528 46912
rect 27580 46900 27586 46912
rect 28350 46900 28356 46912
rect 27580 46872 28356 46900
rect 27580 46860 27586 46872
rect 28350 46860 28356 46872
rect 28408 46900 28414 46912
rect 28905 46903 28963 46909
rect 28905 46900 28917 46903
rect 28408 46872 28917 46900
rect 28408 46860 28414 46872
rect 28905 46869 28917 46872
rect 28951 46869 28963 46903
rect 28905 46863 28963 46869
rect 1104 46810 30820 46832
rect 1104 46758 10880 46810
rect 10932 46758 10944 46810
rect 10996 46758 11008 46810
rect 11060 46758 11072 46810
rect 11124 46758 11136 46810
rect 11188 46758 20811 46810
rect 20863 46758 20875 46810
rect 20927 46758 20939 46810
rect 20991 46758 21003 46810
rect 21055 46758 21067 46810
rect 21119 46758 30820 46810
rect 1104 46736 30820 46758
rect 13170 46696 13176 46708
rect 13131 46668 13176 46696
rect 13170 46656 13176 46668
rect 13228 46656 13234 46708
rect 14182 46656 14188 46708
rect 14240 46696 14246 46708
rect 16482 46696 16488 46708
rect 14240 46668 16488 46696
rect 14240 46656 14246 46668
rect 16482 46656 16488 46668
rect 16540 46656 16546 46708
rect 19058 46696 19064 46708
rect 19019 46668 19064 46696
rect 19058 46656 19064 46668
rect 19116 46656 19122 46708
rect 24946 46656 24952 46708
rect 25004 46696 25010 46708
rect 25225 46699 25283 46705
rect 25225 46696 25237 46699
rect 25004 46668 25237 46696
rect 25004 46656 25010 46668
rect 25225 46665 25237 46668
rect 25271 46665 25283 46699
rect 25225 46659 25283 46665
rect 25685 46699 25743 46705
rect 25685 46665 25697 46699
rect 25731 46696 25743 46699
rect 26510 46696 26516 46708
rect 25731 46668 26516 46696
rect 25731 46665 25743 46668
rect 25685 46659 25743 46665
rect 26510 46656 26516 46668
rect 26568 46656 26574 46708
rect 28718 46656 28724 46708
rect 28776 46696 28782 46708
rect 28902 46696 28908 46708
rect 28776 46668 28908 46696
rect 28776 46656 28782 46668
rect 28902 46656 28908 46668
rect 28960 46656 28966 46708
rect 12802 46588 12808 46640
rect 12860 46628 12866 46640
rect 14200 46628 14228 46656
rect 14458 46628 14464 46640
rect 12860 46600 14228 46628
rect 14419 46600 14464 46628
rect 12860 46588 12866 46600
rect 14458 46588 14464 46600
rect 14516 46588 14522 46640
rect 14645 46631 14703 46637
rect 14645 46597 14657 46631
rect 14691 46628 14703 46631
rect 14734 46628 14740 46640
rect 14691 46600 14740 46628
rect 14691 46597 14703 46600
rect 14645 46591 14703 46597
rect 14734 46588 14740 46600
rect 14792 46588 14798 46640
rect 15562 46588 15568 46640
rect 15620 46628 15626 46640
rect 15933 46631 15991 46637
rect 15933 46628 15945 46631
rect 15620 46600 15945 46628
rect 15620 46588 15626 46600
rect 15933 46597 15945 46600
rect 15979 46628 15991 46631
rect 17221 46631 17279 46637
rect 17221 46628 17233 46631
rect 15979 46600 17233 46628
rect 15979 46597 15991 46600
rect 15933 46591 15991 46597
rect 17221 46597 17233 46600
rect 17267 46628 17279 46631
rect 18141 46631 18199 46637
rect 18141 46628 18153 46631
rect 17267 46600 18153 46628
rect 17267 46597 17279 46600
rect 17221 46591 17279 46597
rect 18141 46597 18153 46600
rect 18187 46597 18199 46631
rect 18141 46591 18199 46597
rect 19426 46588 19432 46640
rect 19484 46628 19490 46640
rect 19521 46631 19579 46637
rect 19521 46628 19533 46631
rect 19484 46600 19533 46628
rect 19484 46588 19490 46600
rect 19521 46597 19533 46600
rect 19567 46597 19579 46631
rect 21266 46628 21272 46640
rect 21227 46600 21272 46628
rect 19521 46591 19579 46597
rect 21266 46588 21272 46600
rect 21324 46588 21330 46640
rect 23382 46628 23388 46640
rect 22020 46600 23388 46628
rect 1394 46520 1400 46572
rect 1452 46560 1458 46572
rect 1581 46563 1639 46569
rect 1581 46560 1593 46563
rect 1452 46532 1593 46560
rect 1452 46520 1458 46532
rect 1581 46529 1593 46532
rect 1627 46529 1639 46563
rect 11882 46560 11888 46572
rect 11843 46532 11888 46560
rect 1581 46523 1639 46529
rect 11882 46520 11888 46532
rect 11940 46520 11946 46572
rect 15654 46520 15660 46572
rect 15712 46560 15718 46572
rect 15749 46563 15807 46569
rect 15749 46560 15761 46563
rect 15712 46532 15761 46560
rect 15712 46520 15718 46532
rect 15749 46529 15761 46532
rect 15795 46560 15807 46563
rect 16206 46560 16212 46572
rect 15795 46532 16212 46560
rect 15795 46529 15807 46532
rect 15749 46523 15807 46529
rect 16206 46520 16212 46532
rect 16264 46560 16270 46572
rect 17037 46563 17095 46569
rect 17037 46560 17049 46563
rect 16264 46532 17049 46560
rect 16264 46520 16270 46532
rect 17037 46529 17049 46532
rect 17083 46529 17095 46563
rect 17954 46560 17960 46572
rect 17915 46532 17960 46560
rect 17037 46523 17095 46529
rect 17954 46520 17960 46532
rect 18012 46520 18018 46572
rect 18874 46560 18880 46572
rect 18835 46532 18880 46560
rect 18874 46520 18880 46532
rect 18932 46520 18938 46572
rect 22020 46569 22048 46600
rect 23382 46588 23388 46600
rect 23440 46588 23446 46640
rect 22005 46563 22063 46569
rect 22005 46529 22017 46563
rect 22051 46529 22063 46563
rect 22005 46523 22063 46529
rect 22097 46563 22155 46569
rect 22097 46529 22109 46563
rect 22143 46560 22155 46563
rect 22370 46560 22376 46572
rect 22143 46532 22376 46560
rect 22143 46529 22155 46532
rect 22097 46523 22155 46529
rect 22370 46520 22376 46532
rect 22428 46520 22434 46572
rect 22738 46520 22744 46572
rect 22796 46560 22802 46572
rect 22922 46560 22928 46572
rect 22796 46532 22928 46560
rect 22796 46520 22802 46532
rect 22922 46520 22928 46532
rect 22980 46520 22986 46572
rect 23106 46520 23112 46572
rect 23164 46560 23170 46572
rect 23293 46563 23351 46569
rect 23293 46560 23305 46563
rect 23164 46532 23305 46560
rect 23164 46520 23170 46532
rect 23293 46529 23305 46532
rect 23339 46529 23351 46563
rect 23474 46560 23480 46572
rect 23435 46532 23480 46560
rect 23293 46523 23351 46529
rect 23474 46520 23480 46532
rect 23532 46520 23538 46572
rect 28810 46520 28816 46572
rect 28868 46560 28874 46572
rect 28905 46563 28963 46569
rect 28905 46560 28917 46563
rect 28868 46532 28917 46560
rect 28868 46520 28874 46532
rect 28905 46529 28917 46532
rect 28951 46529 28963 46563
rect 29730 46560 29736 46572
rect 29691 46532 29736 46560
rect 28905 46523 28963 46529
rect 29730 46520 29736 46532
rect 29788 46520 29794 46572
rect 14550 46452 14556 46504
rect 14608 46492 14614 46504
rect 14737 46495 14795 46501
rect 14737 46492 14749 46495
rect 14608 46464 14749 46492
rect 14608 46452 14614 46464
rect 14737 46461 14749 46464
rect 14783 46461 14795 46495
rect 14737 46455 14795 46461
rect 16025 46495 16083 46501
rect 16025 46461 16037 46495
rect 16071 46492 16083 46495
rect 16298 46492 16304 46504
rect 16071 46464 16304 46492
rect 16071 46461 16083 46464
rect 16025 46455 16083 46461
rect 16298 46452 16304 46464
rect 16356 46492 16362 46504
rect 17313 46495 17371 46501
rect 17313 46492 17325 46495
rect 16356 46464 17325 46492
rect 16356 46452 16362 46464
rect 17313 46461 17325 46464
rect 17359 46461 17371 46495
rect 17313 46455 17371 46461
rect 22281 46495 22339 46501
rect 22281 46461 22293 46495
rect 22327 46492 22339 46495
rect 22462 46492 22468 46504
rect 22327 46464 22468 46492
rect 22327 46461 22339 46464
rect 22281 46455 22339 46461
rect 22462 46452 22468 46464
rect 22520 46452 22526 46504
rect 25409 46495 25467 46501
rect 25409 46461 25421 46495
rect 25455 46461 25467 46495
rect 25409 46455 25467 46461
rect 14185 46427 14243 46433
rect 14185 46393 14197 46427
rect 14231 46424 14243 46427
rect 14826 46424 14832 46436
rect 14231 46396 14832 46424
rect 14231 46393 14243 46396
rect 14185 46387 14243 46393
rect 14826 46384 14832 46396
rect 14884 46384 14890 46436
rect 15470 46424 15476 46436
rect 15431 46396 15476 46424
rect 15470 46384 15476 46396
rect 15528 46384 15534 46436
rect 16761 46427 16819 46433
rect 16761 46393 16773 46427
rect 16807 46424 16819 46427
rect 18322 46424 18328 46436
rect 16807 46396 18328 46424
rect 16807 46393 16819 46396
rect 16761 46387 16819 46393
rect 18322 46384 18328 46396
rect 18380 46384 18386 46436
rect 23106 46384 23112 46436
rect 23164 46424 23170 46436
rect 23290 46424 23296 46436
rect 23164 46396 23296 46424
rect 23164 46384 23170 46396
rect 23290 46384 23296 46396
rect 23348 46384 23354 46436
rect 25424 46424 25452 46455
rect 25498 46452 25504 46504
rect 25556 46492 25562 46504
rect 25774 46492 25780 46504
rect 25556 46464 25601 46492
rect 25735 46464 25780 46492
rect 25556 46452 25562 46464
rect 25774 46452 25780 46464
rect 25832 46452 25838 46504
rect 25869 46495 25927 46501
rect 25869 46461 25881 46495
rect 25915 46492 25927 46495
rect 26050 46492 26056 46504
rect 25915 46464 26056 46492
rect 25915 46461 25927 46464
rect 25869 46455 25927 46461
rect 26050 46452 26056 46464
rect 26108 46492 26114 46504
rect 26510 46492 26516 46504
rect 26108 46464 26516 46492
rect 26108 46452 26114 46464
rect 26510 46452 26516 46464
rect 26568 46452 26574 46504
rect 25424 46396 25544 46424
rect 25516 46368 25544 46396
rect 1397 46359 1455 46365
rect 1397 46325 1409 46359
rect 1443 46356 1455 46359
rect 2406 46356 2412 46368
rect 1443 46328 2412 46356
rect 1443 46325 1455 46328
rect 1397 46319 1455 46325
rect 2406 46316 2412 46328
rect 2464 46316 2470 46368
rect 13814 46316 13820 46368
rect 13872 46356 13878 46368
rect 13998 46356 14004 46368
rect 13872 46328 14004 46356
rect 13872 46316 13878 46328
rect 13998 46316 14004 46328
rect 14056 46356 14062 46368
rect 21450 46356 21456 46368
rect 14056 46328 21456 46356
rect 14056 46316 14062 46328
rect 21450 46316 21456 46328
rect 21508 46316 21514 46368
rect 22186 46316 22192 46368
rect 22244 46356 22250 46368
rect 22244 46328 22289 46356
rect 22244 46316 22250 46328
rect 23014 46316 23020 46368
rect 23072 46356 23078 46368
rect 23385 46359 23443 46365
rect 23385 46356 23397 46359
rect 23072 46328 23397 46356
rect 23072 46316 23078 46328
rect 23385 46325 23397 46328
rect 23431 46325 23443 46359
rect 23385 46319 23443 46325
rect 25498 46316 25504 46368
rect 25556 46316 25562 46368
rect 29086 46356 29092 46368
rect 29047 46328 29092 46356
rect 29086 46316 29092 46328
rect 29144 46316 29150 46368
rect 30009 46359 30067 46365
rect 30009 46325 30021 46359
rect 30055 46356 30067 46359
rect 31110 46356 31116 46368
rect 30055 46328 31116 46356
rect 30055 46325 30067 46328
rect 30009 46319 30067 46325
rect 31110 46316 31116 46328
rect 31168 46316 31174 46368
rect 1104 46266 30820 46288
rect 1104 46214 5915 46266
rect 5967 46214 5979 46266
rect 6031 46214 6043 46266
rect 6095 46214 6107 46266
rect 6159 46214 6171 46266
rect 6223 46214 15846 46266
rect 15898 46214 15910 46266
rect 15962 46214 15974 46266
rect 16026 46214 16038 46266
rect 16090 46214 16102 46266
rect 16154 46214 25776 46266
rect 25828 46214 25840 46266
rect 25892 46214 25904 46266
rect 25956 46214 25968 46266
rect 26020 46214 26032 46266
rect 26084 46214 30820 46266
rect 30926 46248 30932 46300
rect 30984 46288 30990 46300
rect 31386 46288 31392 46300
rect 30984 46260 31392 46288
rect 30984 46248 30990 46260
rect 31386 46248 31392 46260
rect 31444 46248 31450 46300
rect 1104 46192 30820 46214
rect 12713 46155 12771 46161
rect 12713 46121 12725 46155
rect 12759 46152 12771 46155
rect 12894 46152 12900 46164
rect 12759 46124 12900 46152
rect 12759 46121 12771 46124
rect 12713 46115 12771 46121
rect 12894 46112 12900 46124
rect 12952 46112 12958 46164
rect 14642 46152 14648 46164
rect 14603 46124 14648 46152
rect 14642 46112 14648 46124
rect 14700 46112 14706 46164
rect 19886 46112 19892 46164
rect 19944 46152 19950 46164
rect 19981 46155 20039 46161
rect 19981 46152 19993 46155
rect 19944 46124 19993 46152
rect 19944 46112 19950 46124
rect 19981 46121 19993 46124
rect 20027 46121 20039 46155
rect 22278 46152 22284 46164
rect 22239 46124 22284 46152
rect 19981 46115 20039 46121
rect 22278 46112 22284 46124
rect 22336 46152 22342 46164
rect 22336 46124 22784 46152
rect 22336 46112 22342 46124
rect 11609 46087 11667 46093
rect 11609 46053 11621 46087
rect 11655 46053 11667 46087
rect 11609 46047 11667 46053
rect 1486 45908 1492 45960
rect 1544 45948 1550 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 1544 45920 1593 45948
rect 1544 45908 1550 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 2222 45908 2228 45960
rect 2280 45948 2286 45960
rect 2501 45951 2559 45957
rect 2501 45948 2513 45951
rect 2280 45920 2513 45948
rect 2280 45908 2286 45920
rect 2501 45917 2513 45920
rect 2547 45917 2559 45951
rect 2501 45911 2559 45917
rect 10321 45951 10379 45957
rect 10321 45917 10333 45951
rect 10367 45948 10379 45951
rect 11624 45948 11652 46047
rect 12618 46044 12624 46096
rect 12676 46084 12682 46096
rect 13262 46084 13268 46096
rect 12676 46056 13268 46084
rect 12676 46044 12682 46056
rect 13262 46044 13268 46056
rect 13320 46044 13326 46096
rect 14366 46044 14372 46096
rect 14424 46084 14430 46096
rect 17037 46087 17095 46093
rect 17037 46084 17049 46087
rect 14424 46056 17049 46084
rect 14424 46044 14430 46056
rect 17037 46053 17049 46056
rect 17083 46084 17095 46087
rect 17954 46084 17960 46096
rect 17083 46056 17960 46084
rect 17083 46053 17095 46056
rect 17037 46047 17095 46053
rect 17954 46044 17960 46056
rect 18012 46044 18018 46096
rect 22756 46093 22784 46124
rect 22830 46112 22836 46164
rect 22888 46152 22894 46164
rect 23382 46152 23388 46164
rect 22888 46124 23388 46152
rect 22888 46112 22894 46124
rect 23382 46112 23388 46124
rect 23440 46112 23446 46164
rect 26878 46112 26884 46164
rect 26936 46152 26942 46164
rect 27246 46152 27252 46164
rect 26936 46124 27252 46152
rect 26936 46112 26942 46124
rect 27246 46112 27252 46124
rect 27304 46112 27310 46164
rect 29362 46112 29368 46164
rect 29420 46152 29426 46164
rect 29549 46155 29607 46161
rect 29549 46152 29561 46155
rect 29420 46124 29561 46152
rect 29420 46112 29426 46124
rect 29549 46121 29561 46124
rect 29595 46121 29607 46155
rect 31754 46152 31760 46164
rect 29549 46115 29607 46121
rect 31036 46124 31760 46152
rect 31036 46096 31064 46124
rect 31754 46112 31760 46124
rect 31812 46112 31818 46164
rect 22741 46087 22799 46093
rect 22741 46053 22753 46087
rect 22787 46053 22799 46087
rect 22741 46047 22799 46053
rect 25222 46044 25228 46096
rect 25280 46084 25286 46096
rect 25406 46084 25412 46096
rect 25280 46056 25412 46084
rect 25280 46044 25286 46056
rect 25406 46044 25412 46056
rect 25464 46044 25470 46096
rect 31018 46044 31024 46096
rect 31076 46044 31082 46096
rect 31846 46044 31852 46096
rect 31904 46084 31910 46096
rect 31904 46056 31984 46084
rect 31904 46044 31910 46056
rect 12069 46019 12127 46025
rect 12069 45985 12081 46019
rect 12115 46016 12127 46019
rect 12434 46016 12440 46028
rect 12115 45988 12440 46016
rect 12115 45985 12127 45988
rect 12069 45979 12127 45985
rect 12434 45976 12440 45988
rect 12492 45976 12498 46028
rect 13814 46016 13820 46028
rect 13004 45988 13820 46016
rect 13004 45957 13032 45988
rect 13814 45976 13820 45988
rect 13872 45976 13878 46028
rect 18233 46019 18291 46025
rect 18233 46016 18245 46019
rect 15120 45988 18245 46016
rect 10367 45920 11652 45948
rect 12989 45951 13047 45957
rect 10367 45917 10379 45920
rect 10321 45911 10379 45917
rect 12989 45917 13001 45951
rect 13035 45917 13047 45951
rect 12989 45911 13047 45917
rect 13081 45951 13139 45957
rect 13081 45917 13093 45951
rect 13127 45917 13139 45951
rect 13081 45911 13139 45917
rect 13173 45951 13231 45957
rect 13173 45917 13185 45951
rect 13219 45917 13231 45951
rect 13173 45911 13231 45917
rect 2314 45880 2320 45892
rect 2275 45852 2320 45880
rect 2314 45840 2320 45852
rect 2372 45840 2378 45892
rect 11514 45840 11520 45892
rect 11572 45880 11578 45892
rect 12158 45880 12164 45892
rect 11572 45852 12164 45880
rect 11572 45840 11578 45852
rect 12158 45840 12164 45852
rect 12216 45840 12222 45892
rect 12710 45840 12716 45892
rect 12768 45880 12774 45892
rect 13096 45880 13124 45911
rect 12768 45852 13124 45880
rect 12768 45840 12774 45852
rect 1394 45812 1400 45824
rect 1355 45784 1400 45812
rect 1394 45772 1400 45784
rect 1452 45772 1458 45824
rect 2222 45772 2228 45824
rect 2280 45812 2286 45824
rect 2498 45812 2504 45824
rect 2280 45784 2504 45812
rect 2280 45772 2286 45784
rect 2498 45772 2504 45784
rect 2556 45772 2562 45824
rect 2682 45812 2688 45824
rect 2643 45784 2688 45812
rect 2682 45772 2688 45784
rect 2740 45772 2746 45824
rect 10042 45772 10048 45824
rect 10100 45812 10106 45824
rect 10505 45815 10563 45821
rect 10505 45812 10517 45815
rect 10100 45784 10517 45812
rect 10100 45772 10106 45784
rect 10505 45781 10517 45784
rect 10551 45781 10563 45815
rect 10505 45775 10563 45781
rect 11698 45772 11704 45824
rect 11756 45812 11762 45824
rect 11974 45812 11980 45824
rect 11756 45784 11980 45812
rect 11756 45772 11762 45784
rect 11974 45772 11980 45784
rect 12032 45812 12038 45824
rect 12069 45815 12127 45821
rect 12069 45812 12081 45815
rect 12032 45784 12081 45812
rect 12032 45772 12038 45784
rect 12069 45781 12081 45784
rect 12115 45781 12127 45815
rect 12069 45775 12127 45781
rect 12894 45772 12900 45824
rect 12952 45812 12958 45824
rect 13185 45812 13213 45911
rect 13262 45908 13268 45960
rect 13320 45948 13326 45960
rect 15120 45957 15148 45988
rect 18233 45985 18245 45988
rect 18279 46016 18291 46019
rect 18874 46016 18880 46028
rect 18279 45988 18880 46016
rect 18279 45985 18291 45988
rect 18233 45979 18291 45985
rect 18874 45976 18880 45988
rect 18932 45976 18938 46028
rect 20714 45976 20720 46028
rect 20772 46016 20778 46028
rect 20901 46019 20959 46025
rect 20901 46016 20913 46019
rect 20772 45988 20913 46016
rect 20772 45976 20778 45988
rect 20901 45985 20913 45988
rect 20947 45985 20959 46019
rect 20901 45979 20959 45985
rect 21910 45976 21916 46028
rect 21968 46016 21974 46028
rect 21968 45988 22416 46016
rect 21968 45976 21974 45988
rect 13357 45951 13415 45957
rect 13357 45948 13369 45951
rect 13320 45920 13369 45948
rect 13320 45908 13326 45920
rect 13357 45917 13369 45920
rect 13403 45917 13415 45951
rect 13357 45911 13415 45917
rect 14461 45951 14519 45957
rect 14461 45917 14473 45951
rect 14507 45917 14519 45951
rect 14461 45911 14519 45917
rect 15105 45951 15163 45957
rect 15105 45917 15117 45951
rect 15151 45917 15163 45951
rect 15105 45911 15163 45917
rect 21168 45951 21226 45957
rect 21168 45917 21180 45951
rect 21214 45948 21226 45951
rect 22186 45948 22192 45960
rect 21214 45920 22192 45948
rect 21214 45917 21226 45920
rect 21168 45911 21226 45917
rect 14476 45880 14504 45911
rect 22186 45908 22192 45920
rect 22244 45908 22250 45960
rect 15194 45880 15200 45892
rect 14476 45852 15200 45880
rect 15194 45840 15200 45852
rect 15252 45840 15258 45892
rect 15746 45880 15752 45892
rect 15707 45852 15752 45880
rect 15746 45840 15752 45852
rect 15804 45840 15810 45892
rect 18049 45883 18107 45889
rect 18049 45849 18061 45883
rect 18095 45880 18107 45883
rect 18230 45880 18236 45892
rect 18095 45852 18236 45880
rect 18095 45849 18107 45852
rect 18049 45843 18107 45849
rect 18230 45840 18236 45852
rect 18288 45840 18294 45892
rect 19886 45880 19892 45892
rect 19847 45852 19892 45880
rect 19886 45840 19892 45852
rect 19944 45840 19950 45892
rect 22388 45880 22416 45988
rect 22462 45976 22468 46028
rect 22520 46016 22526 46028
rect 22830 46016 22836 46028
rect 22520 45988 22836 46016
rect 22520 45976 22526 45988
rect 22830 45976 22836 45988
rect 22888 45976 22894 46028
rect 23293 46019 23351 46025
rect 23293 45985 23305 46019
rect 23339 45985 23351 46019
rect 23293 45979 23351 45985
rect 23014 45948 23020 45960
rect 22975 45920 23020 45948
rect 23014 45908 23020 45920
rect 23072 45908 23078 45960
rect 23308 45880 23336 45979
rect 25038 45976 25044 46028
rect 25096 46016 25102 46028
rect 25682 46016 25688 46028
rect 25096 45988 25688 46016
rect 25096 45976 25102 45988
rect 25682 45976 25688 45988
rect 25740 46016 25746 46028
rect 25777 46019 25835 46025
rect 25777 46016 25789 46019
rect 25740 45988 25789 46016
rect 25740 45976 25746 45988
rect 25777 45985 25789 45988
rect 25823 45985 25835 46019
rect 25777 45979 25835 45985
rect 25501 45951 25559 45957
rect 25501 45917 25513 45951
rect 25547 45917 25559 45951
rect 25501 45911 25559 45917
rect 21928 45852 22094 45880
rect 22388 45852 23336 45880
rect 24857 45883 24915 45889
rect 13262 45812 13268 45824
rect 12952 45784 13268 45812
rect 12952 45772 12958 45784
rect 13262 45772 13268 45784
rect 13320 45772 13326 45824
rect 15289 45815 15347 45821
rect 15289 45781 15301 45815
rect 15335 45812 15347 45815
rect 16942 45812 16948 45824
rect 15335 45784 16948 45812
rect 15335 45781 15347 45784
rect 15289 45775 15347 45781
rect 16942 45772 16948 45784
rect 17000 45772 17006 45824
rect 17402 45772 17408 45824
rect 17460 45812 17466 45824
rect 21928 45812 21956 45852
rect 17460 45784 21956 45812
rect 22066 45812 22094 45852
rect 24857 45849 24869 45883
rect 24903 45880 24915 45883
rect 25406 45880 25412 45892
rect 24903 45852 25412 45880
rect 24903 45849 24915 45852
rect 24857 45843 24915 45849
rect 25406 45840 25412 45852
rect 25464 45880 25470 45892
rect 25516 45880 25544 45911
rect 29178 45908 29184 45960
rect 29236 45948 29242 45960
rect 29362 45948 29368 45960
rect 29236 45920 29368 45948
rect 29236 45908 29242 45920
rect 29362 45908 29368 45920
rect 29420 45908 29426 45960
rect 29730 45948 29736 45960
rect 29691 45920 29736 45948
rect 29730 45908 29736 45920
rect 29788 45908 29794 45960
rect 30006 45948 30012 45960
rect 29967 45920 30012 45948
rect 30006 45908 30012 45920
rect 30064 45908 30070 45960
rect 25464 45852 25544 45880
rect 25464 45840 25470 45852
rect 28350 45840 28356 45892
rect 28408 45880 28414 45892
rect 29748 45880 29776 45908
rect 28408 45852 29776 45880
rect 28408 45840 28414 45852
rect 22925 45815 22983 45821
rect 22925 45812 22937 45815
rect 22066 45784 22937 45812
rect 17460 45772 17466 45784
rect 22925 45781 22937 45784
rect 22971 45812 22983 45815
rect 23014 45812 23020 45824
rect 22971 45784 23020 45812
rect 22971 45781 22983 45784
rect 22925 45775 22983 45781
rect 23014 45772 23020 45784
rect 23072 45772 23078 45824
rect 23109 45815 23167 45821
rect 23109 45781 23121 45815
rect 23155 45812 23167 45815
rect 23290 45812 23296 45824
rect 23155 45784 23296 45812
rect 23155 45781 23167 45784
rect 23109 45775 23167 45781
rect 23290 45772 23296 45784
rect 23348 45772 23354 45824
rect 23750 45772 23756 45824
rect 23808 45812 23814 45824
rect 24026 45812 24032 45824
rect 23808 45784 24032 45812
rect 23808 45772 23814 45784
rect 24026 45772 24032 45784
rect 24084 45812 24090 45824
rect 24949 45815 25007 45821
rect 24949 45812 24961 45815
rect 24084 45784 24961 45812
rect 24084 45772 24090 45784
rect 24949 45781 24961 45784
rect 24995 45781 25007 45815
rect 24949 45775 25007 45781
rect 25314 45772 25320 45824
rect 25372 45812 25378 45824
rect 25682 45812 25688 45824
rect 25372 45784 25688 45812
rect 25372 45772 25378 45784
rect 25682 45772 25688 45784
rect 25740 45772 25746 45824
rect 29178 45772 29184 45824
rect 29236 45812 29242 45824
rect 29917 45815 29975 45821
rect 29917 45812 29929 45815
rect 29236 45784 29929 45812
rect 29236 45772 29242 45784
rect 29917 45781 29929 45784
rect 29963 45781 29975 45815
rect 31956 45812 31984 46056
rect 29917 45775 29975 45781
rect 31772 45784 31984 45812
rect 1104 45722 30820 45744
rect 1104 45670 10880 45722
rect 10932 45670 10944 45722
rect 10996 45670 11008 45722
rect 11060 45670 11072 45722
rect 11124 45670 11136 45722
rect 11188 45670 20811 45722
rect 20863 45670 20875 45722
rect 20927 45670 20939 45722
rect 20991 45670 21003 45722
rect 21055 45670 21067 45722
rect 21119 45670 30820 45722
rect 1104 45648 30820 45670
rect 2682 45568 2688 45620
rect 2740 45608 2746 45620
rect 13998 45608 14004 45620
rect 2740 45580 14004 45608
rect 2740 45568 2746 45580
rect 13998 45568 14004 45580
rect 14056 45568 14062 45620
rect 15746 45568 15752 45620
rect 15804 45608 15810 45620
rect 16117 45611 16175 45617
rect 16117 45608 16129 45611
rect 15804 45580 16129 45608
rect 15804 45568 15810 45580
rect 16117 45577 16129 45580
rect 16163 45577 16175 45611
rect 16117 45571 16175 45577
rect 20346 45568 20352 45620
rect 20404 45568 20410 45620
rect 24305 45611 24363 45617
rect 24305 45577 24317 45611
rect 24351 45608 24363 45611
rect 24670 45608 24676 45620
rect 24351 45580 24676 45608
rect 24351 45577 24363 45580
rect 24305 45571 24363 45577
rect 24670 45568 24676 45580
rect 24728 45568 24734 45620
rect 25314 45608 25320 45620
rect 24872 45580 25320 45608
rect 2314 45540 2320 45552
rect 2275 45512 2320 45540
rect 2314 45500 2320 45512
rect 2372 45500 2378 45552
rect 2406 45500 2412 45552
rect 2464 45540 2470 45552
rect 2501 45543 2559 45549
rect 2501 45540 2513 45543
rect 2464 45512 2513 45540
rect 2464 45500 2470 45512
rect 2501 45509 2513 45512
rect 2547 45509 2559 45543
rect 12526 45540 12532 45552
rect 12487 45512 12532 45540
rect 2501 45503 2559 45509
rect 12526 45500 12532 45512
rect 12584 45500 12590 45552
rect 12802 45540 12808 45552
rect 12800 45500 12808 45540
rect 12860 45500 12866 45552
rect 13262 45540 13268 45552
rect 13096 45512 13268 45540
rect 1578 45472 1584 45484
rect 1539 45444 1584 45472
rect 1578 45432 1584 45444
rect 1636 45432 1642 45484
rect 12800 45481 12828 45500
rect 12759 45475 12828 45481
rect 12759 45441 12771 45475
rect 12805 45444 12828 45475
rect 12897 45475 12955 45481
rect 12805 45441 12817 45444
rect 12759 45435 12817 45441
rect 12897 45441 12909 45475
rect 12943 45441 12955 45475
rect 12897 45435 12955 45441
rect 13010 45475 13068 45481
rect 13010 45441 13022 45475
rect 13056 45472 13068 45475
rect 13096 45472 13124 45512
rect 13262 45500 13268 45512
rect 13320 45500 13326 45552
rect 16942 45500 16948 45552
rect 17000 45540 17006 45552
rect 17037 45543 17095 45549
rect 17037 45540 17049 45543
rect 17000 45512 17049 45540
rect 17000 45500 17006 45512
rect 17037 45509 17049 45512
rect 17083 45509 17095 45543
rect 17037 45503 17095 45509
rect 18414 45500 18420 45552
rect 18472 45540 18478 45552
rect 18601 45543 18659 45549
rect 18601 45540 18613 45543
rect 18472 45512 18613 45540
rect 18472 45500 18478 45512
rect 18601 45509 18613 45512
rect 18647 45509 18659 45543
rect 18601 45503 18659 45509
rect 13056 45444 13124 45472
rect 13173 45475 13231 45481
rect 13056 45441 13068 45444
rect 13010 45435 13068 45441
rect 13173 45441 13185 45475
rect 13219 45441 13231 45475
rect 13722 45472 13728 45484
rect 13683 45444 13728 45472
rect 13173 45435 13231 45441
rect 12526 45364 12532 45416
rect 12584 45404 12590 45416
rect 12912 45404 12940 45435
rect 12584 45376 12940 45404
rect 12584 45364 12590 45376
rect 7466 45296 7472 45348
rect 7524 45336 7530 45348
rect 13188 45336 13216 45435
rect 13722 45432 13728 45444
rect 13780 45432 13786 45484
rect 14182 45432 14188 45484
rect 14240 45472 14246 45484
rect 15933 45475 15991 45481
rect 15933 45472 15945 45475
rect 14240 45444 15945 45472
rect 14240 45432 14246 45444
rect 15933 45441 15945 45444
rect 15979 45441 15991 45475
rect 15933 45435 15991 45441
rect 18506 45432 18512 45484
rect 18564 45472 18570 45484
rect 19245 45475 19303 45481
rect 19245 45472 19257 45475
rect 18564 45444 19257 45472
rect 18564 45432 18570 45444
rect 19245 45441 19257 45444
rect 19291 45441 19303 45475
rect 19245 45435 19303 45441
rect 20257 45475 20315 45481
rect 20257 45441 20269 45475
rect 20303 45441 20315 45475
rect 20257 45435 20315 45441
rect 7524 45308 13216 45336
rect 7524 45296 7530 45308
rect 13354 45296 13360 45348
rect 13412 45336 13418 45348
rect 15013 45339 15071 45345
rect 15013 45336 15025 45339
rect 13412 45308 15025 45336
rect 13412 45296 13418 45308
rect 15013 45305 15025 45308
rect 15059 45305 15071 45339
rect 19978 45336 19984 45348
rect 19939 45308 19984 45336
rect 15013 45299 15071 45305
rect 19978 45296 19984 45308
rect 20036 45296 20042 45348
rect 20272 45336 20300 45435
rect 20364 45404 20392 45568
rect 20441 45543 20499 45549
rect 20441 45509 20453 45543
rect 20487 45540 20499 45543
rect 21174 45540 21180 45552
rect 20487 45512 21180 45540
rect 20487 45509 20499 45512
rect 20441 45503 20499 45509
rect 21174 45500 21180 45512
rect 21232 45500 21238 45552
rect 22094 45500 22100 45552
rect 22152 45540 22158 45552
rect 22646 45540 22652 45552
rect 22152 45512 22652 45540
rect 22152 45500 22158 45512
rect 22646 45500 22652 45512
rect 22704 45500 22710 45552
rect 24397 45543 24455 45549
rect 24397 45509 24409 45543
rect 24443 45540 24455 45543
rect 24762 45540 24768 45552
rect 24443 45512 24768 45540
rect 24443 45509 24455 45512
rect 24397 45503 24455 45509
rect 24762 45500 24768 45512
rect 24820 45540 24826 45552
rect 24872 45540 24900 45580
rect 25314 45568 25320 45580
rect 25372 45568 25378 45620
rect 25409 45611 25467 45617
rect 25409 45577 25421 45611
rect 25455 45608 25467 45611
rect 25455 45580 25636 45608
rect 25455 45577 25467 45580
rect 25409 45571 25467 45577
rect 24820 45512 24900 45540
rect 24820 45500 24826 45512
rect 24946 45500 24952 45552
rect 25004 45540 25010 45552
rect 25498 45540 25504 45552
rect 25004 45512 25504 45540
rect 25004 45500 25010 45512
rect 25498 45500 25504 45512
rect 25556 45500 25562 45552
rect 25608 45540 25636 45580
rect 28902 45568 28908 45620
rect 28960 45608 28966 45620
rect 29181 45611 29239 45617
rect 29181 45608 29193 45611
rect 28960 45580 29193 45608
rect 28960 45568 28966 45580
rect 29181 45577 29193 45580
rect 29227 45577 29239 45611
rect 29181 45571 29239 45577
rect 26418 45540 26424 45552
rect 25608 45512 26424 45540
rect 26418 45500 26424 45512
rect 26476 45500 26482 45552
rect 27798 45500 27804 45552
rect 27856 45540 27862 45552
rect 28629 45543 28687 45549
rect 28629 45540 28641 45543
rect 27856 45512 28641 45540
rect 27856 45500 27862 45512
rect 28629 45509 28641 45512
rect 28675 45509 28687 45543
rect 29730 45540 29736 45552
rect 28629 45503 28687 45509
rect 29380 45512 29736 45540
rect 20714 45432 20720 45484
rect 20772 45472 20778 45484
rect 21085 45475 21143 45481
rect 21085 45472 21097 45475
rect 20772 45444 21097 45472
rect 20772 45432 20778 45444
rect 21085 45441 21097 45444
rect 21131 45441 21143 45475
rect 21910 45472 21916 45484
rect 21871 45444 21916 45472
rect 21085 45435 21143 45441
rect 21910 45432 21916 45444
rect 21968 45432 21974 45484
rect 22462 45432 22468 45484
rect 22520 45472 22526 45484
rect 23750 45472 23756 45484
rect 22520 45444 23756 45472
rect 22520 45432 22526 45444
rect 23750 45432 23756 45444
rect 23808 45472 23814 45484
rect 24121 45475 24179 45481
rect 24121 45472 24133 45475
rect 23808 45444 24133 45472
rect 23808 45432 23814 45444
rect 24121 45441 24133 45444
rect 24167 45441 24179 45475
rect 25593 45475 25651 45481
rect 25593 45472 25605 45475
rect 24121 45435 24179 45441
rect 24780 45444 25605 45472
rect 20533 45407 20591 45413
rect 20533 45404 20545 45407
rect 20364 45376 20545 45404
rect 20533 45373 20545 45376
rect 20579 45404 20591 45407
rect 20898 45404 20904 45416
rect 20579 45376 20904 45404
rect 20579 45373 20591 45376
rect 20533 45367 20591 45373
rect 20898 45364 20904 45376
rect 20956 45364 20962 45416
rect 20990 45364 20996 45416
rect 21048 45404 21054 45416
rect 22097 45407 22155 45413
rect 22097 45404 22109 45407
rect 21048 45376 22109 45404
rect 21048 45364 21054 45376
rect 22097 45373 22109 45376
rect 22143 45373 22155 45407
rect 24026 45404 24032 45416
rect 23987 45376 24032 45404
rect 22097 45367 22155 45373
rect 24026 45364 24032 45376
rect 24084 45364 24090 45416
rect 21008 45336 21036 45364
rect 20272 45308 21036 45336
rect 24136 45336 24164 45435
rect 24780 45416 24808 45444
rect 25593 45441 25605 45444
rect 25639 45441 25651 45475
rect 25593 45435 25651 45441
rect 28350 45432 28356 45484
rect 28408 45472 28414 45484
rect 29380 45481 29408 45512
rect 29730 45500 29736 45512
rect 29788 45500 29794 45552
rect 28445 45475 28503 45481
rect 28445 45472 28457 45475
rect 28408 45444 28457 45472
rect 28408 45432 28414 45444
rect 28445 45441 28457 45444
rect 28491 45441 28503 45475
rect 28721 45475 28779 45481
rect 28721 45472 28733 45475
rect 28445 45435 28503 45441
rect 28552 45444 28733 45472
rect 28552 45416 28580 45444
rect 28721 45441 28733 45444
rect 28767 45441 28779 45475
rect 28721 45435 28779 45441
rect 29365 45475 29423 45481
rect 29365 45441 29377 45475
rect 29411 45441 29423 45475
rect 29546 45472 29552 45484
rect 29507 45444 29552 45472
rect 29365 45435 29423 45441
rect 29546 45432 29552 45444
rect 29604 45432 29610 45484
rect 29641 45475 29699 45481
rect 29641 45441 29653 45475
rect 29687 45441 29699 45475
rect 29641 45435 29699 45441
rect 24489 45407 24547 45413
rect 24489 45373 24501 45407
rect 24535 45404 24547 45407
rect 24762 45404 24768 45416
rect 24535 45376 24768 45404
rect 24535 45373 24547 45376
rect 24489 45367 24547 45373
rect 24762 45364 24768 45376
rect 24820 45364 24826 45416
rect 25038 45364 25044 45416
rect 25096 45404 25102 45416
rect 25133 45407 25191 45413
rect 25133 45404 25145 45407
rect 25096 45376 25145 45404
rect 25096 45364 25102 45376
rect 25133 45373 25145 45376
rect 25179 45373 25191 45407
rect 25133 45367 25191 45373
rect 25225 45407 25283 45413
rect 25225 45373 25237 45407
rect 25271 45373 25283 45407
rect 25225 45367 25283 45373
rect 25240 45336 25268 45367
rect 25314 45364 25320 45416
rect 25372 45404 25378 45416
rect 25501 45407 25559 45413
rect 25501 45404 25513 45407
rect 25372 45376 25513 45404
rect 25372 45364 25378 45376
rect 25501 45373 25513 45376
rect 25547 45373 25559 45407
rect 25501 45367 25559 45373
rect 28534 45364 28540 45416
rect 28592 45404 28598 45416
rect 29656 45404 29684 45435
rect 30006 45404 30012 45416
rect 28592 45376 30012 45404
rect 28592 45364 28598 45376
rect 30006 45364 30012 45376
rect 30064 45364 30070 45416
rect 29270 45336 29276 45348
rect 24136 45308 25268 45336
rect 28276 45308 29276 45336
rect 1397 45271 1455 45277
rect 1397 45237 1409 45271
rect 1443 45268 1455 45271
rect 1762 45268 1768 45280
rect 1443 45240 1768 45268
rect 1443 45237 1455 45240
rect 1397 45231 1455 45237
rect 1762 45228 1768 45240
rect 1820 45228 1826 45280
rect 2685 45271 2743 45277
rect 2685 45237 2697 45271
rect 2731 45268 2743 45271
rect 12618 45268 12624 45280
rect 2731 45240 12624 45268
rect 2731 45237 2743 45240
rect 2685 45231 2743 45237
rect 12618 45228 12624 45240
rect 12676 45228 12682 45280
rect 19429 45271 19487 45277
rect 19429 45237 19441 45271
rect 19475 45268 19487 45271
rect 19518 45268 19524 45280
rect 19475 45240 19524 45268
rect 19475 45237 19487 45240
rect 19429 45231 19487 45237
rect 19518 45228 19524 45240
rect 19576 45228 19582 45280
rect 21177 45271 21235 45277
rect 21177 45237 21189 45271
rect 21223 45268 21235 45271
rect 22462 45268 22468 45280
rect 21223 45240 22468 45268
rect 21223 45237 21235 45240
rect 21177 45231 21235 45237
rect 22462 45228 22468 45240
rect 22520 45228 22526 45280
rect 23845 45271 23903 45277
rect 23845 45237 23857 45271
rect 23891 45268 23903 45271
rect 24670 45268 24676 45280
rect 23891 45240 24676 45268
rect 23891 45237 23903 45240
rect 23845 45231 23903 45237
rect 24670 45228 24676 45240
rect 24728 45228 24734 45280
rect 24946 45268 24952 45280
rect 24907 45240 24952 45268
rect 24946 45228 24952 45240
rect 25004 45228 25010 45280
rect 28276 45277 28304 45308
rect 29270 45296 29276 45308
rect 29328 45296 29334 45348
rect 31772 45280 31800 45784
rect 31846 45704 31852 45756
rect 31904 45704 31910 45756
rect 28261 45271 28319 45277
rect 28261 45237 28273 45271
rect 28307 45237 28319 45271
rect 28261 45231 28319 45237
rect 28902 45228 28908 45280
rect 28960 45268 28966 45280
rect 29086 45268 29092 45280
rect 28960 45240 29092 45268
rect 28960 45228 28966 45240
rect 29086 45228 29092 45240
rect 29144 45228 29150 45280
rect 31754 45228 31760 45280
rect 31812 45228 31818 45280
rect 1104 45178 30820 45200
rect 1104 45126 5915 45178
rect 5967 45126 5979 45178
rect 6031 45126 6043 45178
rect 6095 45126 6107 45178
rect 6159 45126 6171 45178
rect 6223 45126 15846 45178
rect 15898 45126 15910 45178
rect 15962 45126 15974 45178
rect 16026 45126 16038 45178
rect 16090 45126 16102 45178
rect 16154 45126 25776 45178
rect 25828 45126 25840 45178
rect 25892 45126 25904 45178
rect 25956 45126 25968 45178
rect 26020 45126 26032 45178
rect 26084 45126 30820 45178
rect 1104 45104 30820 45126
rect 1949 45067 2007 45073
rect 1949 45033 1961 45067
rect 1995 45064 2007 45067
rect 7466 45064 7472 45076
rect 1995 45036 7472 45064
rect 1995 45033 2007 45036
rect 1949 45027 2007 45033
rect 7466 45024 7472 45036
rect 7524 45024 7530 45076
rect 11977 45067 12035 45073
rect 11977 45033 11989 45067
rect 12023 45064 12035 45067
rect 12250 45064 12256 45076
rect 12023 45036 12256 45064
rect 12023 45033 12035 45036
rect 11977 45027 12035 45033
rect 12250 45024 12256 45036
rect 12308 45024 12314 45076
rect 16758 45024 16764 45076
rect 16816 45064 16822 45076
rect 16942 45064 16948 45076
rect 16816 45036 16948 45064
rect 16816 45024 16822 45036
rect 16942 45024 16948 45036
rect 17000 45064 17006 45076
rect 18233 45067 18291 45073
rect 18233 45064 18245 45067
rect 17000 45036 18245 45064
rect 17000 45024 17006 45036
rect 18233 45033 18245 45036
rect 18279 45033 18291 45067
rect 18233 45027 18291 45033
rect 20533 45067 20591 45073
rect 20533 45033 20545 45067
rect 20579 45064 20591 45067
rect 22278 45064 22284 45076
rect 20579 45036 22284 45064
rect 20579 45033 20591 45036
rect 20533 45027 20591 45033
rect 22278 45024 22284 45036
rect 22336 45024 22342 45076
rect 28718 45024 28724 45076
rect 28776 45064 28782 45076
rect 29549 45067 29607 45073
rect 29549 45064 29561 45067
rect 28776 45036 29561 45064
rect 28776 45024 28782 45036
rect 29549 45033 29561 45036
rect 29595 45033 29607 45067
rect 29549 45027 29607 45033
rect 31864 45008 31892 45704
rect 13078 44996 13084 45008
rect 12084 44968 13084 44996
rect 10042 44928 10048 44940
rect 10003 44900 10048 44928
rect 10042 44888 10048 44900
rect 10100 44888 10106 44940
rect 1394 44820 1400 44872
rect 1452 44860 1458 44872
rect 1765 44863 1823 44869
rect 1765 44860 1777 44863
rect 1452 44832 1777 44860
rect 1452 44820 1458 44832
rect 1765 44829 1777 44832
rect 1811 44829 1823 44863
rect 12084 44860 12112 44968
rect 13078 44956 13084 44968
rect 13136 44956 13142 45008
rect 19337 44999 19395 45005
rect 19337 44965 19349 44999
rect 19383 44996 19395 44999
rect 19426 44996 19432 45008
rect 19383 44968 19432 44996
rect 19383 44965 19395 44968
rect 19337 44959 19395 44965
rect 19426 44956 19432 44968
rect 19484 44956 19490 45008
rect 20898 44956 20904 45008
rect 20956 44996 20962 45008
rect 20956 44968 21128 44996
rect 20956 44956 20962 44968
rect 12894 44928 12900 44940
rect 12452 44900 12900 44928
rect 12452 44869 12480 44900
rect 12894 44888 12900 44900
rect 12952 44888 12958 44940
rect 19794 44928 19800 44940
rect 19755 44900 19800 44928
rect 19794 44888 19800 44900
rect 19852 44888 19858 44940
rect 20990 44928 20996 44940
rect 20951 44900 20996 44928
rect 20990 44888 20996 44900
rect 21048 44888 21054 44940
rect 21100 44937 21128 44968
rect 24486 44956 24492 45008
rect 24544 44996 24550 45008
rect 26326 44996 26332 45008
rect 24544 44968 26332 44996
rect 24544 44956 24550 44968
rect 26326 44956 26332 44968
rect 26384 44956 26390 45008
rect 28077 44999 28135 45005
rect 28077 44965 28089 44999
rect 28123 44996 28135 44999
rect 29086 44996 29092 45008
rect 28123 44968 29092 44996
rect 28123 44965 28135 44968
rect 28077 44959 28135 44965
rect 29086 44956 29092 44968
rect 29144 44956 29150 45008
rect 29270 44956 29276 45008
rect 29328 44996 29334 45008
rect 29638 44996 29644 45008
rect 29328 44968 29644 44996
rect 29328 44956 29334 44968
rect 29638 44956 29644 44968
rect 29696 44956 29702 45008
rect 31846 44956 31852 45008
rect 31904 44956 31910 45008
rect 21085 44931 21143 44937
rect 21085 44897 21097 44931
rect 21131 44897 21143 44931
rect 25038 44928 25044 44940
rect 24999 44900 25044 44928
rect 21085 44891 21143 44897
rect 12207 44863 12265 44869
rect 12207 44860 12219 44863
rect 12084 44832 12219 44860
rect 1765 44823 1823 44829
rect 12207 44829 12219 44832
rect 12253 44829 12265 44863
rect 12207 44823 12265 44829
rect 12345 44863 12403 44869
rect 12345 44829 12357 44863
rect 12391 44829 12403 44863
rect 12345 44823 12403 44829
rect 12437 44863 12495 44869
rect 12437 44829 12449 44863
rect 12483 44829 12495 44863
rect 12437 44823 12495 44829
rect 12633 44863 12691 44869
rect 12633 44829 12645 44863
rect 12679 44860 12691 44863
rect 12986 44860 12992 44872
rect 12679 44832 12992 44860
rect 12679 44829 12691 44832
rect 12633 44823 12691 44829
rect 1581 44795 1639 44801
rect 1581 44761 1593 44795
rect 1627 44792 1639 44795
rect 1670 44792 1676 44804
rect 1627 44764 1676 44792
rect 1627 44761 1639 44764
rect 1581 44755 1639 44761
rect 1670 44752 1676 44764
rect 1728 44752 1734 44804
rect 9766 44752 9772 44804
rect 9824 44792 9830 44804
rect 10290 44795 10348 44801
rect 10290 44792 10302 44795
rect 9824 44764 10302 44792
rect 9824 44752 9830 44764
rect 10290 44761 10302 44764
rect 10336 44761 10348 44795
rect 12373 44792 12401 44823
rect 12986 44820 12992 44832
rect 13044 44820 13050 44872
rect 13354 44860 13360 44872
rect 13315 44832 13360 44860
rect 13354 44820 13360 44832
rect 13412 44820 13418 44872
rect 13906 44820 13912 44872
rect 13964 44860 13970 44872
rect 17126 44860 17132 44872
rect 13964 44832 17132 44860
rect 13964 44820 13970 44832
rect 17126 44820 17132 44832
rect 17184 44820 17190 44872
rect 19334 44820 19340 44872
rect 19392 44860 19398 44872
rect 21100 44860 21128 44891
rect 25038 44888 25044 44900
rect 25096 44888 25102 44940
rect 25314 44888 25320 44940
rect 25372 44928 25378 44940
rect 25409 44931 25467 44937
rect 25409 44928 25421 44931
rect 25372 44900 25421 44928
rect 25372 44888 25378 44900
rect 25409 44897 25421 44900
rect 25455 44897 25467 44931
rect 25409 44891 25467 44897
rect 28350 44888 28356 44940
rect 28408 44928 28414 44940
rect 28902 44928 28908 44940
rect 28408 44900 28908 44928
rect 28408 44888 28414 44900
rect 28902 44888 28908 44900
rect 28960 44888 28966 44940
rect 19392 44832 21128 44860
rect 21913 44863 21971 44869
rect 19392 44820 19398 44832
rect 21913 44829 21925 44863
rect 21959 44860 21971 44863
rect 22180 44863 22238 44869
rect 21959 44832 22094 44860
rect 21959 44829 21971 44832
rect 21913 44823 21971 44829
rect 12526 44792 12532 44804
rect 12373 44764 12532 44792
rect 10290 44755 10348 44761
rect 12526 44752 12532 44764
rect 12584 44752 12590 44804
rect 14461 44795 14519 44801
rect 14461 44761 14473 44795
rect 14507 44792 14519 44795
rect 15286 44792 15292 44804
rect 14507 44764 15292 44792
rect 14507 44761 14519 44764
rect 14461 44755 14519 44761
rect 15286 44752 15292 44764
rect 15344 44752 15350 44804
rect 16945 44795 17003 44801
rect 16945 44761 16957 44795
rect 16991 44792 17003 44795
rect 17862 44792 17868 44804
rect 16991 44764 17868 44792
rect 16991 44761 17003 44764
rect 16945 44755 17003 44761
rect 17862 44752 17868 44764
rect 17920 44752 17926 44804
rect 19889 44795 19947 44801
rect 19889 44761 19901 44795
rect 19935 44792 19947 44795
rect 19978 44792 19984 44804
rect 19935 44764 19984 44792
rect 19935 44761 19947 44764
rect 19889 44755 19947 44761
rect 19978 44752 19984 44764
rect 20036 44792 20042 44804
rect 20622 44792 20628 44804
rect 20036 44764 20628 44792
rect 20036 44752 20042 44764
rect 20622 44752 20628 44764
rect 20680 44752 20686 44804
rect 10410 44684 10416 44736
rect 10468 44724 10474 44736
rect 11425 44727 11483 44733
rect 11425 44724 11437 44727
rect 10468 44696 11437 44724
rect 10468 44684 10474 44696
rect 11425 44693 11437 44696
rect 11471 44724 11483 44727
rect 13262 44724 13268 44736
rect 11471 44696 13268 44724
rect 11471 44693 11483 44696
rect 11425 44687 11483 44693
rect 13262 44684 13268 44696
rect 13320 44684 13326 44736
rect 13449 44727 13507 44733
rect 13449 44693 13461 44727
rect 13495 44724 13507 44727
rect 14642 44724 14648 44736
rect 13495 44696 14648 44724
rect 13495 44693 13507 44696
rect 13449 44687 13507 44693
rect 14642 44684 14648 44696
rect 14700 44684 14706 44736
rect 15746 44724 15752 44736
rect 15707 44696 15752 44724
rect 15746 44684 15752 44696
rect 15804 44684 15810 44736
rect 19797 44727 19855 44733
rect 19797 44693 19809 44727
rect 19843 44724 19855 44727
rect 20993 44727 21051 44733
rect 20993 44724 21005 44727
rect 19843 44696 21005 44724
rect 19843 44693 19855 44696
rect 19797 44687 19855 44693
rect 20993 44693 21005 44696
rect 21039 44724 21051 44727
rect 21174 44724 21180 44736
rect 21039 44696 21180 44724
rect 21039 44693 21051 44696
rect 20993 44687 21051 44693
rect 21174 44684 21180 44696
rect 21232 44684 21238 44736
rect 22066 44724 22094 44832
rect 22180 44829 22192 44863
rect 22226 44860 22238 44863
rect 22646 44860 22652 44872
rect 22226 44832 22652 44860
rect 22226 44829 22238 44832
rect 22180 44823 22238 44829
rect 22646 44820 22652 44832
rect 22704 44820 22710 44872
rect 23658 44820 23664 44872
rect 23716 44820 23722 44872
rect 23750 44820 23756 44872
rect 23808 44860 23814 44872
rect 24486 44860 24492 44872
rect 23808 44832 24492 44860
rect 23808 44820 23814 44832
rect 24486 44820 24492 44832
rect 24544 44860 24550 44872
rect 25133 44863 25191 44869
rect 25133 44860 25145 44863
rect 24544 44832 25145 44860
rect 24544 44820 24550 44832
rect 25133 44829 25145 44832
rect 25179 44829 25191 44863
rect 25133 44823 25191 44829
rect 25501 44863 25559 44869
rect 25501 44829 25513 44863
rect 25547 44829 25559 44863
rect 27154 44860 27160 44872
rect 27115 44832 27160 44860
rect 25501 44823 25559 44829
rect 22370 44752 22376 44804
rect 22428 44792 22434 44804
rect 23676 44792 23704 44820
rect 22428 44764 23704 44792
rect 22428 44752 22434 44764
rect 24762 44752 24768 44804
rect 24820 44792 24826 44804
rect 25516 44792 25544 44823
rect 27154 44820 27160 44832
rect 27212 44820 27218 44872
rect 28258 44860 28264 44872
rect 28219 44832 28264 44860
rect 28258 44820 28264 44832
rect 28316 44820 28322 44872
rect 28718 44860 28724 44872
rect 28679 44832 28724 44860
rect 28718 44820 28724 44832
rect 28776 44820 28782 44872
rect 29730 44860 29736 44872
rect 29691 44832 29736 44860
rect 29730 44820 29736 44832
rect 29788 44820 29794 44872
rect 30006 44860 30012 44872
rect 29967 44832 30012 44860
rect 30006 44820 30012 44832
rect 30064 44820 30070 44872
rect 24820 44764 25544 44792
rect 24820 44752 24826 44764
rect 22646 44724 22652 44736
rect 22066 44696 22652 44724
rect 22646 44684 22652 44696
rect 22704 44684 22710 44736
rect 23293 44727 23351 44733
rect 23293 44693 23305 44727
rect 23339 44724 23351 44727
rect 23658 44724 23664 44736
rect 23339 44696 23664 44724
rect 23339 44693 23351 44696
rect 23293 44687 23351 44693
rect 23658 44684 23664 44696
rect 23716 44684 23722 44736
rect 24857 44727 24915 44733
rect 24857 44693 24869 44727
rect 24903 44724 24915 44727
rect 25038 44724 25044 44736
rect 24903 44696 25044 44724
rect 24903 44693 24915 44696
rect 24857 44687 24915 44693
rect 25038 44684 25044 44696
rect 25096 44684 25102 44736
rect 25130 44684 25136 44736
rect 25188 44724 25194 44736
rect 25225 44727 25283 44733
rect 25225 44724 25237 44727
rect 25188 44696 25237 44724
rect 25188 44684 25194 44696
rect 25225 44693 25237 44696
rect 25271 44693 25283 44727
rect 25225 44687 25283 44693
rect 26878 44684 26884 44736
rect 26936 44724 26942 44736
rect 27341 44727 27399 44733
rect 27341 44724 27353 44727
rect 26936 44696 27353 44724
rect 26936 44684 26942 44696
rect 27341 44693 27353 44696
rect 27387 44693 27399 44727
rect 28902 44724 28908 44736
rect 28863 44696 28908 44724
rect 27341 44687 27399 44693
rect 28902 44684 28908 44696
rect 28960 44684 28966 44736
rect 29638 44684 29644 44736
rect 29696 44724 29702 44736
rect 29917 44727 29975 44733
rect 29917 44724 29929 44727
rect 29696 44696 29929 44724
rect 29696 44684 29702 44696
rect 29917 44693 29929 44696
rect 29963 44693 29975 44727
rect 29917 44687 29975 44693
rect 1104 44634 30820 44656
rect 1104 44582 10880 44634
rect 10932 44582 10944 44634
rect 10996 44582 11008 44634
rect 11060 44582 11072 44634
rect 11124 44582 11136 44634
rect 11188 44582 20811 44634
rect 20863 44582 20875 44634
rect 20927 44582 20939 44634
rect 20991 44582 21003 44634
rect 21055 44582 21067 44634
rect 21119 44582 30820 44634
rect 1104 44560 30820 44582
rect 2409 44523 2467 44529
rect 2409 44520 2421 44523
rect 1780 44492 2421 44520
rect 1581 44455 1639 44461
rect 1581 44421 1593 44455
rect 1627 44452 1639 44455
rect 1670 44452 1676 44464
rect 1627 44424 1676 44452
rect 1627 44421 1639 44424
rect 1581 44415 1639 44421
rect 1670 44412 1676 44424
rect 1728 44412 1734 44464
rect 1780 44461 1808 44492
rect 2409 44489 2421 44492
rect 2455 44489 2467 44523
rect 2409 44483 2467 44489
rect 2590 44480 2596 44532
rect 2648 44520 2654 44532
rect 12342 44520 12348 44532
rect 2648 44492 7604 44520
rect 2648 44480 2654 44492
rect 1765 44455 1823 44461
rect 1765 44421 1777 44455
rect 1811 44421 1823 44455
rect 1765 44415 1823 44421
rect 2593 44387 2651 44393
rect 2593 44353 2605 44387
rect 2639 44384 2651 44387
rect 2774 44384 2780 44396
rect 2639 44356 2780 44384
rect 2639 44353 2651 44356
rect 2593 44347 2651 44353
rect 2774 44344 2780 44356
rect 2832 44344 2838 44396
rect 7576 44384 7604 44492
rect 10796 44492 12348 44520
rect 10796 44461 10824 44492
rect 12342 44480 12348 44492
rect 12400 44480 12406 44532
rect 12434 44480 12440 44532
rect 12492 44520 12498 44532
rect 13081 44523 13139 44529
rect 13081 44520 13093 44523
rect 12492 44492 13093 44520
rect 12492 44480 12498 44492
rect 13081 44489 13093 44492
rect 13127 44489 13139 44523
rect 13081 44483 13139 44489
rect 14734 44480 14740 44532
rect 14792 44520 14798 44532
rect 15933 44523 15991 44529
rect 15933 44520 15945 44523
rect 14792 44492 15945 44520
rect 14792 44480 14798 44492
rect 15933 44489 15945 44492
rect 15979 44489 15991 44523
rect 15933 44483 15991 44489
rect 16751 44523 16809 44529
rect 16751 44489 16763 44523
rect 16797 44520 16809 44523
rect 17770 44520 17776 44532
rect 16797 44492 17776 44520
rect 16797 44489 16809 44492
rect 16751 44483 16809 44489
rect 17770 44480 17776 44492
rect 17828 44480 17834 44532
rect 19886 44480 19892 44532
rect 19944 44520 19950 44532
rect 20622 44520 20628 44532
rect 19944 44492 20628 44520
rect 19944 44480 19950 44492
rect 20622 44480 20628 44492
rect 20680 44520 20686 44532
rect 20809 44523 20867 44529
rect 20809 44520 20821 44523
rect 20680 44492 20821 44520
rect 20680 44480 20686 44492
rect 20809 44489 20821 44492
rect 20855 44489 20867 44523
rect 20809 44483 20867 44489
rect 23658 44480 23664 44532
rect 23716 44480 23722 44532
rect 24486 44520 24492 44532
rect 24447 44492 24492 44520
rect 24486 44480 24492 44492
rect 24544 44480 24550 44532
rect 27154 44480 27160 44532
rect 27212 44520 27218 44532
rect 27430 44520 27436 44532
rect 27212 44492 27436 44520
rect 27212 44480 27218 44492
rect 27430 44480 27436 44492
rect 27488 44480 27494 44532
rect 29273 44523 29331 44529
rect 29273 44489 29285 44523
rect 29319 44520 29331 44523
rect 30006 44520 30012 44532
rect 29319 44492 30012 44520
rect 29319 44489 29331 44492
rect 29273 44483 29331 44489
rect 30006 44480 30012 44492
rect 30064 44480 30070 44532
rect 10781 44455 10839 44461
rect 10781 44421 10793 44455
rect 10827 44421 10839 44455
rect 10781 44415 10839 44421
rect 10965 44455 11023 44461
rect 10965 44421 10977 44455
rect 11011 44452 11023 44455
rect 11698 44452 11704 44464
rect 11011 44424 11704 44452
rect 11011 44421 11023 44424
rect 10965 44415 11023 44421
rect 11698 44412 11704 44424
rect 11756 44412 11762 44464
rect 12802 44452 12808 44464
rect 12268 44424 12808 44452
rect 11606 44384 11612 44396
rect 7576 44356 11612 44384
rect 11606 44344 11612 44356
rect 11664 44344 11670 44396
rect 12066 44384 12072 44396
rect 12027 44356 12072 44384
rect 12066 44344 12072 44356
rect 12124 44344 12130 44396
rect 12268 44393 12296 44424
rect 12802 44412 12808 44424
rect 12860 44412 12866 44464
rect 12989 44455 13047 44461
rect 12989 44421 13001 44455
rect 13035 44452 13047 44455
rect 13170 44452 13176 44464
rect 13035 44424 13176 44452
rect 13035 44421 13047 44424
rect 12989 44415 13047 44421
rect 13170 44412 13176 44424
rect 13228 44412 13234 44464
rect 14182 44452 14188 44464
rect 14143 44424 14188 44452
rect 14182 44412 14188 44424
rect 14240 44412 14246 44464
rect 15470 44452 15476 44464
rect 14752 44424 15476 44452
rect 12158 44387 12216 44393
rect 12158 44353 12170 44387
rect 12204 44353 12216 44387
rect 12158 44347 12216 44353
rect 12253 44387 12311 44393
rect 12253 44353 12265 44387
rect 12299 44353 12311 44387
rect 12253 44347 12311 44353
rect 12437 44387 12495 44393
rect 12437 44353 12449 44387
rect 12483 44384 12495 44387
rect 12526 44384 12532 44396
rect 12483 44356 12532 44384
rect 12483 44353 12495 44356
rect 12437 44347 12495 44353
rect 11790 44316 11796 44328
rect 11751 44288 11796 44316
rect 11790 44276 11796 44288
rect 11848 44276 11854 44328
rect 12176 44316 12204 44347
rect 12526 44344 12532 44356
rect 12584 44344 12590 44396
rect 14752 44393 14780 44424
rect 15470 44412 15476 44424
rect 15528 44412 15534 44464
rect 15654 44412 15660 44464
rect 15712 44452 15718 44464
rect 15749 44455 15807 44461
rect 15749 44452 15761 44455
rect 15712 44424 15761 44452
rect 15712 44412 15718 44424
rect 15749 44421 15761 44424
rect 15795 44421 15807 44455
rect 15749 44415 15807 44421
rect 16025 44455 16083 44461
rect 16025 44421 16037 44455
rect 16071 44452 16083 44455
rect 16298 44452 16304 44464
rect 16071 44424 16304 44452
rect 16071 44421 16083 44424
rect 16025 44415 16083 44421
rect 14001 44387 14059 44393
rect 14001 44353 14013 44387
rect 14047 44353 14059 44387
rect 14001 44347 14059 44353
rect 14737 44387 14795 44393
rect 14737 44353 14749 44387
rect 14783 44353 14795 44387
rect 14737 44347 14795 44353
rect 14921 44387 14979 44393
rect 14921 44353 14933 44387
rect 14967 44384 14979 44387
rect 16040 44384 16068 44415
rect 16298 44412 16304 44424
rect 16356 44412 16362 44464
rect 17218 44452 17224 44464
rect 17179 44424 17224 44452
rect 17218 44412 17224 44424
rect 17276 44412 17282 44464
rect 17678 44412 17684 44464
rect 17736 44452 17742 44464
rect 19518 44452 19524 44464
rect 17736 44424 18368 44452
rect 19479 44424 19524 44452
rect 17736 44412 17742 44424
rect 14967 44356 16068 44384
rect 16316 44384 16344 44412
rect 18340 44396 18368 44424
rect 19518 44412 19524 44424
rect 19576 44412 19582 44464
rect 21266 44412 21272 44464
rect 21324 44452 21330 44464
rect 21913 44455 21971 44461
rect 21913 44452 21925 44455
rect 21324 44424 21925 44452
rect 21324 44412 21330 44424
rect 21913 44421 21925 44424
rect 21959 44421 21971 44455
rect 21913 44415 21971 44421
rect 23290 44412 23296 44464
rect 23348 44452 23354 44464
rect 23676 44452 23704 44480
rect 24397 44455 24455 44461
rect 24397 44452 24409 44455
rect 23348 44424 23612 44452
rect 23676 44424 24409 44452
rect 23348 44412 23354 44424
rect 17313 44387 17371 44393
rect 17313 44384 17325 44387
rect 16316 44356 17325 44384
rect 14967 44353 14979 44356
rect 14921 44347 14979 44353
rect 17313 44353 17325 44356
rect 17359 44353 17371 44387
rect 17313 44347 17371 44353
rect 12710 44316 12716 44328
rect 12176 44288 12716 44316
rect 12710 44276 12716 44288
rect 12768 44276 12774 44328
rect 14016 44316 14044 44347
rect 18046 44344 18052 44396
rect 18104 44384 18110 44396
rect 18141 44387 18199 44393
rect 18141 44384 18153 44387
rect 18104 44356 18153 44384
rect 18104 44344 18110 44356
rect 18141 44353 18153 44356
rect 18187 44353 18199 44387
rect 18141 44347 18199 44353
rect 18233 44387 18291 44393
rect 18233 44353 18245 44387
rect 18279 44353 18291 44387
rect 18233 44347 18291 44353
rect 17126 44316 17132 44328
rect 14016 44288 15976 44316
rect 17087 44288 17132 44316
rect 1949 44251 2007 44257
rect 1949 44217 1961 44251
rect 1995 44248 2007 44251
rect 1995 44220 2774 44248
rect 1995 44217 2007 44220
rect 1949 44211 2007 44217
rect 2746 44180 2774 44220
rect 12066 44208 12072 44260
rect 12124 44248 12130 44260
rect 13538 44248 13544 44260
rect 12124 44220 13544 44248
rect 12124 44208 12130 44220
rect 13538 44208 13544 44220
rect 13596 44208 13602 44260
rect 15378 44208 15384 44260
rect 15436 44248 15442 44260
rect 15473 44251 15531 44257
rect 15473 44248 15485 44251
rect 15436 44220 15485 44248
rect 15436 44208 15442 44220
rect 15473 44217 15485 44220
rect 15519 44217 15531 44251
rect 15948 44248 15976 44288
rect 17126 44276 17132 44288
rect 17184 44276 17190 44328
rect 17586 44276 17592 44328
rect 17644 44316 17650 44328
rect 18248 44316 18276 44347
rect 18322 44344 18328 44396
rect 18380 44384 18386 44396
rect 18509 44387 18567 44393
rect 18380 44356 18425 44384
rect 18380 44344 18386 44356
rect 18509 44353 18521 44387
rect 18555 44384 18567 44387
rect 18598 44384 18604 44396
rect 18555 44356 18604 44384
rect 18555 44353 18567 44356
rect 18509 44347 18567 44353
rect 18598 44344 18604 44356
rect 18656 44344 18662 44396
rect 22649 44387 22707 44393
rect 22649 44353 22661 44387
rect 22695 44384 22707 44387
rect 22738 44384 22744 44396
rect 22695 44356 22744 44384
rect 22695 44353 22707 44356
rect 22649 44347 22707 44353
rect 22738 44344 22744 44356
rect 22796 44344 22802 44396
rect 23477 44387 23535 44393
rect 23477 44353 23489 44387
rect 23523 44353 23535 44387
rect 23477 44347 23535 44353
rect 17644 44288 18276 44316
rect 17644 44276 17650 44288
rect 19242 44276 19248 44328
rect 19300 44316 19306 44328
rect 19518 44316 19524 44328
rect 19300 44288 19524 44316
rect 19300 44276 19306 44288
rect 19518 44276 19524 44288
rect 19576 44276 19582 44328
rect 16574 44248 16580 44260
rect 15948 44220 16580 44248
rect 15473 44211 15531 44217
rect 16574 44208 16580 44220
rect 16632 44208 16638 44260
rect 23492 44248 23520 44347
rect 23584 44316 23612 44424
rect 24397 44421 24409 44424
rect 24443 44452 24455 44455
rect 24670 44452 24676 44464
rect 24443 44424 24676 44452
rect 24443 44421 24455 44424
rect 24397 44415 24455 44421
rect 24670 44412 24676 44424
rect 24728 44412 24734 44464
rect 27617 44455 27675 44461
rect 27617 44421 27629 44455
rect 27663 44452 27675 44455
rect 28350 44452 28356 44464
rect 27663 44424 28356 44452
rect 27663 44421 27675 44424
rect 27617 44415 27675 44421
rect 28350 44412 28356 44424
rect 28408 44412 28414 44464
rect 23661 44387 23719 44393
rect 23661 44353 23673 44387
rect 23707 44384 23719 44387
rect 23750 44384 23756 44396
rect 23707 44356 23756 44384
rect 23707 44353 23719 44356
rect 23661 44347 23719 44353
rect 23750 44344 23756 44356
rect 23808 44344 23814 44396
rect 25498 44344 25504 44396
rect 25556 44384 25562 44396
rect 25593 44387 25651 44393
rect 25593 44384 25605 44387
rect 25556 44356 25605 44384
rect 25556 44344 25562 44356
rect 25593 44353 25605 44356
rect 25639 44353 25651 44387
rect 25593 44347 25651 44353
rect 26878 44344 26884 44396
rect 26936 44384 26942 44396
rect 27801 44387 27859 44393
rect 27801 44384 27813 44387
rect 26936 44356 27813 44384
rect 26936 44344 26942 44356
rect 27801 44353 27813 44356
rect 27847 44353 27859 44387
rect 27982 44384 27988 44396
rect 27943 44356 27988 44384
rect 27801 44347 27859 44353
rect 27982 44344 27988 44356
rect 28040 44344 28046 44396
rect 28077 44387 28135 44393
rect 28077 44353 28089 44387
rect 28123 44384 28135 44387
rect 28258 44384 28264 44396
rect 28123 44356 28264 44384
rect 28123 44353 28135 44356
rect 28077 44347 28135 44353
rect 28258 44344 28264 44356
rect 28316 44384 28322 44396
rect 28534 44384 28540 44396
rect 28316 44356 28540 44384
rect 28316 44344 28322 44356
rect 28534 44344 28540 44356
rect 28592 44344 28598 44396
rect 28810 44344 28816 44396
rect 28868 44384 28874 44396
rect 29089 44387 29147 44393
rect 29089 44384 29101 44387
rect 28868 44356 29101 44384
rect 28868 44344 28874 44356
rect 29089 44353 29101 44356
rect 29135 44353 29147 44387
rect 29822 44384 29828 44396
rect 29783 44356 29828 44384
rect 29089 44347 29147 44353
rect 29822 44344 29828 44356
rect 29880 44344 29886 44396
rect 23845 44319 23903 44325
rect 23845 44316 23857 44319
rect 23584 44288 23857 44316
rect 23845 44285 23857 44288
rect 23891 44285 23903 44319
rect 23845 44279 23903 44285
rect 25314 44276 25320 44328
rect 25372 44316 25378 44328
rect 25869 44319 25927 44325
rect 25869 44316 25881 44319
rect 25372 44288 25881 44316
rect 25372 44276 25378 44288
rect 25869 44285 25881 44288
rect 25915 44285 25927 44319
rect 25869 44279 25927 44285
rect 24486 44248 24492 44260
rect 23492 44220 24492 44248
rect 24486 44208 24492 44220
rect 24544 44208 24550 44260
rect 30006 44248 30012 44260
rect 29967 44220 30012 44248
rect 30006 44208 30012 44220
rect 30064 44208 30070 44260
rect 12986 44180 12992 44192
rect 2746 44152 12992 44180
rect 12986 44140 12992 44152
rect 13044 44140 13050 44192
rect 17678 44140 17684 44192
rect 17736 44180 17742 44192
rect 17865 44183 17923 44189
rect 17865 44180 17877 44183
rect 17736 44152 17877 44180
rect 17736 44140 17742 44152
rect 17865 44149 17877 44152
rect 17911 44149 17923 44183
rect 17865 44143 17923 44149
rect 18046 44140 18052 44192
rect 18104 44180 18110 44192
rect 18782 44180 18788 44192
rect 18104 44152 18788 44180
rect 18104 44140 18110 44152
rect 18782 44140 18788 44152
rect 18840 44140 18846 44192
rect 20990 44140 20996 44192
rect 21048 44180 21054 44192
rect 22005 44183 22063 44189
rect 22005 44180 22017 44183
rect 21048 44152 22017 44180
rect 21048 44140 21054 44152
rect 22005 44149 22017 44152
rect 22051 44149 22063 44183
rect 22005 44143 22063 44149
rect 22833 44183 22891 44189
rect 22833 44149 22845 44183
rect 22879 44180 22891 44183
rect 23290 44180 23296 44192
rect 22879 44152 23296 44180
rect 22879 44149 22891 44152
rect 22833 44143 22891 44149
rect 23290 44140 23296 44152
rect 23348 44140 23354 44192
rect 1104 44090 30820 44112
rect 1104 44038 5915 44090
rect 5967 44038 5979 44090
rect 6031 44038 6043 44090
rect 6095 44038 6107 44090
rect 6159 44038 6171 44090
rect 6223 44038 15846 44090
rect 15898 44038 15910 44090
rect 15962 44038 15974 44090
rect 16026 44038 16038 44090
rect 16090 44038 16102 44090
rect 16154 44038 25776 44090
rect 25828 44038 25840 44090
rect 25892 44038 25904 44090
rect 25956 44038 25968 44090
rect 26020 44038 26032 44090
rect 26084 44038 30820 44090
rect 1104 44016 30820 44038
rect 2777 43979 2835 43985
rect 2777 43945 2789 43979
rect 2823 43976 2835 43979
rect 12526 43976 12532 43988
rect 2823 43948 12532 43976
rect 2823 43945 2835 43948
rect 2777 43939 2835 43945
rect 12526 43936 12532 43948
rect 12584 43936 12590 43988
rect 13541 43979 13599 43985
rect 13541 43945 13553 43979
rect 13587 43976 13599 43979
rect 13722 43976 13728 43988
rect 13587 43948 13728 43976
rect 13587 43945 13599 43948
rect 13541 43939 13599 43945
rect 13722 43936 13728 43948
rect 13780 43936 13786 43988
rect 15194 43936 15200 43988
rect 15252 43976 15258 43988
rect 15381 43979 15439 43985
rect 15381 43976 15393 43979
rect 15252 43948 15393 43976
rect 15252 43936 15258 43948
rect 15381 43945 15393 43948
rect 15427 43945 15439 43979
rect 15381 43939 15439 43945
rect 16574 43936 16580 43988
rect 16632 43976 16638 43988
rect 17770 43976 17776 43988
rect 16632 43948 17776 43976
rect 16632 43936 16638 43948
rect 17770 43936 17776 43948
rect 17828 43976 17834 43988
rect 17865 43979 17923 43985
rect 17865 43976 17877 43979
rect 17828 43948 17877 43976
rect 17828 43936 17834 43948
rect 17865 43945 17877 43948
rect 17911 43945 17923 43979
rect 17865 43939 17923 43945
rect 19702 43936 19708 43988
rect 19760 43976 19766 43988
rect 22649 43979 22707 43985
rect 22649 43976 22661 43979
rect 19760 43948 22661 43976
rect 19760 43936 19766 43948
rect 22649 43945 22661 43948
rect 22695 43945 22707 43979
rect 22649 43939 22707 43945
rect 23385 43979 23443 43985
rect 23385 43945 23397 43979
rect 23431 43976 23443 43979
rect 24302 43976 24308 43988
rect 23431 43948 24308 43976
rect 23431 43945 23443 43948
rect 23385 43939 23443 43945
rect 24302 43936 24308 43948
rect 24360 43936 24366 43988
rect 26326 43936 26332 43988
rect 26384 43976 26390 43988
rect 26881 43979 26939 43985
rect 26881 43976 26893 43979
rect 26384 43948 26893 43976
rect 26384 43936 26390 43948
rect 26881 43945 26893 43948
rect 26927 43945 26939 43979
rect 26881 43939 26939 43945
rect 9674 43868 9680 43920
rect 9732 43908 9738 43920
rect 10873 43911 10931 43917
rect 10873 43908 10885 43911
rect 9732 43880 10885 43908
rect 9732 43868 9738 43880
rect 10873 43877 10885 43880
rect 10919 43877 10931 43911
rect 10873 43871 10931 43877
rect 12710 43868 12716 43920
rect 12768 43868 12774 43920
rect 12986 43868 12992 43920
rect 13044 43908 13050 43920
rect 14185 43911 14243 43917
rect 14185 43908 14197 43911
rect 13044 43880 14197 43908
rect 13044 43868 13050 43880
rect 14185 43877 14197 43880
rect 14231 43877 14243 43911
rect 14185 43871 14243 43877
rect 19150 43868 19156 43920
rect 19208 43908 19214 43920
rect 19337 43911 19395 43917
rect 19337 43908 19349 43911
rect 19208 43880 19349 43908
rect 19208 43868 19214 43880
rect 19337 43877 19349 43880
rect 19383 43877 19395 43911
rect 19337 43871 19395 43877
rect 19886 43868 19892 43920
rect 19944 43908 19950 43920
rect 20533 43911 20591 43917
rect 20533 43908 20545 43911
rect 19944 43880 20545 43908
rect 19944 43868 19950 43880
rect 20533 43877 20545 43880
rect 20579 43877 20591 43911
rect 20533 43871 20591 43877
rect 23750 43868 23756 43920
rect 23808 43908 23814 43920
rect 23808 43880 23888 43908
rect 23808 43868 23814 43880
rect 10410 43840 10416 43852
rect 9948 43812 10416 43840
rect 1762 43772 1768 43784
rect 1723 43744 1768 43772
rect 1762 43732 1768 43744
rect 1820 43732 1826 43784
rect 9948 43781 9976 43812
rect 10410 43800 10416 43812
rect 10468 43800 10474 43852
rect 11333 43843 11391 43849
rect 11333 43809 11345 43843
rect 11379 43840 11391 43843
rect 12342 43840 12348 43852
rect 11379 43812 12348 43840
rect 11379 43809 11391 43812
rect 11333 43803 11391 43809
rect 12342 43800 12348 43812
rect 12400 43800 12406 43852
rect 12728 43840 12756 43868
rect 14366 43840 14372 43852
rect 12617 43812 14372 43840
rect 9933 43775 9991 43781
rect 9933 43741 9945 43775
rect 9979 43741 9991 43775
rect 9933 43735 9991 43741
rect 10042 43772 10100 43778
rect 10042 43738 10054 43772
rect 10088 43738 10100 43772
rect 10042 43732 10100 43738
rect 1581 43707 1639 43713
rect 1581 43673 1593 43707
rect 1627 43704 1639 43707
rect 1670 43704 1676 43716
rect 1627 43676 1676 43704
rect 1627 43673 1639 43676
rect 1581 43667 1639 43673
rect 1670 43664 1676 43676
rect 1728 43704 1734 43716
rect 2409 43707 2467 43713
rect 2409 43704 2421 43707
rect 1728 43676 2421 43704
rect 1728 43664 1734 43676
rect 2409 43673 2421 43676
rect 2455 43673 2467 43707
rect 2590 43704 2596 43716
rect 2551 43676 2596 43704
rect 2409 43667 2467 43673
rect 2590 43664 2596 43676
rect 2648 43664 2654 43716
rect 9677 43707 9735 43713
rect 9677 43673 9689 43707
rect 9723 43704 9735 43707
rect 9766 43704 9772 43716
rect 9723 43676 9772 43704
rect 9723 43673 9735 43676
rect 9677 43667 9735 43673
rect 9766 43664 9772 43676
rect 9824 43664 9830 43716
rect 10057 43704 10085 43732
rect 10134 43729 10140 43781
rect 10192 43769 10198 43781
rect 10318 43772 10324 43784
rect 10192 43741 10237 43769
rect 10279 43744 10324 43772
rect 10192 43729 10198 43741
rect 10318 43732 10324 43744
rect 10376 43732 10382 43784
rect 12617 43781 12645 43812
rect 14366 43800 14372 43812
rect 14424 43800 14430 43852
rect 14550 43800 14556 43852
rect 14608 43840 14614 43852
rect 14737 43843 14795 43849
rect 14737 43840 14749 43843
rect 14608 43812 14749 43840
rect 14608 43800 14614 43812
rect 14737 43809 14749 43812
rect 14783 43809 14795 43843
rect 14737 43803 14795 43809
rect 15841 43843 15899 43849
rect 15841 43809 15853 43843
rect 15887 43840 15899 43843
rect 17126 43840 17132 43852
rect 15887 43812 17132 43840
rect 15887 43809 15899 43812
rect 15841 43803 15899 43809
rect 17126 43800 17132 43812
rect 17184 43800 17190 43852
rect 19794 43840 19800 43852
rect 19707 43812 19800 43840
rect 19794 43800 19800 43812
rect 19852 43840 19858 43852
rect 20990 43840 20996 43852
rect 19852 43812 20996 43840
rect 19852 43800 19858 43812
rect 20990 43800 20996 43812
rect 21048 43800 21054 43852
rect 23569 43843 23627 43849
rect 23569 43809 23581 43843
rect 23615 43840 23627 43843
rect 23658 43840 23664 43852
rect 23615 43812 23664 43840
rect 23615 43809 23627 43812
rect 23569 43803 23627 43809
rect 23658 43800 23664 43812
rect 23716 43800 23722 43852
rect 23860 43840 23888 43880
rect 24486 43840 24492 43852
rect 23860 43812 24492 43840
rect 12509 43775 12567 43781
rect 12509 43741 12521 43775
rect 12555 43741 12567 43775
rect 12509 43735 12567 43741
rect 12602 43775 12660 43781
rect 12602 43741 12614 43775
rect 12648 43741 12660 43775
rect 12602 43735 12660 43741
rect 12713 43775 12771 43781
rect 12713 43741 12725 43775
rect 12759 43772 12771 43775
rect 12802 43772 12808 43784
rect 12759 43744 12808 43772
rect 12759 43741 12771 43744
rect 12713 43735 12771 43741
rect 9968 43676 10085 43704
rect 11425 43707 11483 43713
rect 9968 43648 9996 43676
rect 11425 43673 11437 43707
rect 11471 43704 11483 43707
rect 11514 43704 11520 43716
rect 11471 43676 11520 43704
rect 11471 43673 11483 43676
rect 11425 43667 11483 43673
rect 11514 43664 11520 43676
rect 11572 43664 11578 43716
rect 12524 43704 12552 43735
rect 12802 43732 12808 43744
rect 12860 43732 12866 43784
rect 12897 43775 12955 43781
rect 12897 43741 12909 43775
rect 12943 43772 12955 43775
rect 13078 43772 13084 43784
rect 12943 43744 13084 43772
rect 12943 43741 12955 43744
rect 12897 43735 12955 43741
rect 13078 43732 13084 43744
rect 13136 43732 13142 43784
rect 13357 43775 13415 43781
rect 13357 43741 13369 43775
rect 13403 43772 13415 43775
rect 14182 43772 14188 43784
rect 13403 43744 14188 43772
rect 13403 43741 13415 43744
rect 13357 43735 13415 43741
rect 14182 43732 14188 43744
rect 14240 43732 14246 43784
rect 15933 43775 15991 43781
rect 15933 43741 15945 43775
rect 15979 43772 15991 43775
rect 16298 43772 16304 43784
rect 15979 43744 16304 43772
rect 15979 43741 15991 43744
rect 15933 43735 15991 43741
rect 16298 43732 16304 43744
rect 16356 43732 16362 43784
rect 16390 43732 16396 43784
rect 16448 43772 16454 43784
rect 19889 43775 19947 43781
rect 16448 43744 19380 43772
rect 16448 43732 16454 43744
rect 14090 43704 14096 43716
rect 12524 43676 14096 43704
rect 14090 43664 14096 43676
rect 14148 43664 14154 43716
rect 14458 43704 14464 43716
rect 14419 43676 14464 43704
rect 14458 43664 14464 43676
rect 14516 43664 14522 43716
rect 14642 43704 14648 43716
rect 14603 43676 14648 43704
rect 14642 43664 14648 43676
rect 14700 43664 14706 43716
rect 15562 43664 15568 43716
rect 15620 43704 15626 43716
rect 15841 43707 15899 43713
rect 15841 43704 15853 43707
rect 15620 43676 15853 43704
rect 15620 43664 15626 43676
rect 15841 43673 15853 43676
rect 15887 43673 15899 43707
rect 15841 43667 15899 43673
rect 16577 43707 16635 43713
rect 16577 43673 16589 43707
rect 16623 43704 16635 43707
rect 19242 43704 19248 43716
rect 16623 43676 19248 43704
rect 16623 43673 16635 43676
rect 16577 43667 16635 43673
rect 19242 43664 19248 43676
rect 19300 43664 19306 43716
rect 19352 43704 19380 43744
rect 19889 43741 19901 43775
rect 19935 43772 19947 43775
rect 19978 43772 19984 43784
rect 19935 43744 19984 43772
rect 19935 43741 19947 43744
rect 19889 43735 19947 43741
rect 19978 43732 19984 43744
rect 20036 43772 20042 43784
rect 21085 43775 21143 43781
rect 21085 43772 21097 43775
rect 20036 43744 21097 43772
rect 20036 43732 20042 43744
rect 21085 43741 21097 43744
rect 21131 43741 21143 43775
rect 22002 43772 22008 43784
rect 21963 43744 22008 43772
rect 21085 43735 21143 43741
rect 22002 43732 22008 43744
rect 22060 43732 22066 43784
rect 22462 43772 22468 43784
rect 22423 43744 22468 43772
rect 22462 43732 22468 43744
rect 22520 43732 22526 43784
rect 23750 43772 23756 43784
rect 23711 43744 23756 43772
rect 23750 43732 23756 43744
rect 23808 43732 23814 43784
rect 23860 43781 23888 43812
rect 24486 43800 24492 43812
rect 24544 43800 24550 43852
rect 24670 43840 24676 43852
rect 24631 43812 24676 43840
rect 24670 43800 24676 43812
rect 24728 43800 24734 43852
rect 28258 43840 28264 43852
rect 28219 43812 28264 43840
rect 28258 43800 28264 43812
rect 28316 43800 28322 43852
rect 23845 43775 23903 43781
rect 23845 43741 23857 43775
rect 23891 43741 23903 43775
rect 23845 43735 23903 43741
rect 24026 43732 24032 43784
rect 24084 43772 24090 43784
rect 24581 43775 24639 43781
rect 24581 43772 24593 43775
rect 24084 43744 24593 43772
rect 24084 43732 24090 43744
rect 24581 43741 24593 43744
rect 24627 43741 24639 43775
rect 24581 43735 24639 43741
rect 24762 43732 24768 43784
rect 24820 43772 24826 43784
rect 25041 43775 25099 43781
rect 25041 43772 25053 43775
rect 24820 43744 25053 43772
rect 24820 43732 24826 43744
rect 25041 43741 25053 43744
rect 25087 43741 25099 43775
rect 25041 43735 25099 43741
rect 26878 43732 26884 43784
rect 26936 43772 26942 43784
rect 27065 43775 27123 43781
rect 27065 43772 27077 43775
rect 26936 43744 27077 43772
rect 26936 43732 26942 43744
rect 27065 43741 27077 43744
rect 27111 43741 27123 43775
rect 27065 43735 27123 43741
rect 27341 43775 27399 43781
rect 27341 43741 27353 43775
rect 27387 43741 27399 43775
rect 27341 43735 27399 43741
rect 27985 43775 28043 43781
rect 27985 43741 27997 43775
rect 28031 43772 28043 43775
rect 28350 43772 28356 43784
rect 28031 43744 28356 43772
rect 28031 43741 28043 43744
rect 27985 43735 28043 43741
rect 27356 43704 27384 43735
rect 28350 43732 28356 43744
rect 28408 43732 28414 43784
rect 29822 43772 29828 43784
rect 29783 43744 29828 43772
rect 29822 43732 29828 43744
rect 29880 43732 29886 43784
rect 28258 43704 28264 43716
rect 19352 43676 24808 43704
rect 27356 43676 28264 43704
rect 1946 43636 1952 43648
rect 1907 43608 1952 43636
rect 1946 43596 1952 43608
rect 2004 43596 2010 43648
rect 9950 43596 9956 43648
rect 10008 43596 10014 43648
rect 11333 43639 11391 43645
rect 11333 43605 11345 43639
rect 11379 43636 11391 43639
rect 12158 43636 12164 43648
rect 11379 43608 12164 43636
rect 11379 43605 11391 43608
rect 11333 43599 11391 43605
rect 12158 43596 12164 43608
rect 12216 43596 12222 43648
rect 12253 43639 12311 43645
rect 12253 43605 12265 43639
rect 12299 43636 12311 43639
rect 13078 43636 13084 43648
rect 12299 43608 13084 43636
rect 12299 43605 12311 43608
rect 12253 43599 12311 43605
rect 13078 43596 13084 43608
rect 13136 43596 13142 43648
rect 19797 43639 19855 43645
rect 19797 43605 19809 43639
rect 19843 43636 19855 43639
rect 20162 43636 20168 43648
rect 19843 43608 20168 43636
rect 19843 43605 19855 43608
rect 19797 43599 19855 43605
rect 20162 43596 20168 43608
rect 20220 43636 20226 43648
rect 20993 43639 21051 43645
rect 20993 43636 21005 43639
rect 20220 43608 21005 43636
rect 20220 43596 20226 43608
rect 20993 43605 21005 43608
rect 21039 43605 21051 43639
rect 20993 43599 21051 43605
rect 21821 43639 21879 43645
rect 21821 43605 21833 43639
rect 21867 43636 21879 43639
rect 22186 43636 22192 43648
rect 21867 43608 22192 43636
rect 21867 43605 21879 43608
rect 21821 43599 21879 43605
rect 22186 43596 22192 43608
rect 22244 43596 22250 43648
rect 23750 43596 23756 43648
rect 23808 43636 23814 43648
rect 24780 43645 24808 43676
rect 28258 43664 28264 43676
rect 28316 43664 28322 43716
rect 24397 43639 24455 43645
rect 24397 43636 24409 43639
rect 23808 43608 24409 43636
rect 23808 43596 23814 43608
rect 24397 43605 24409 43608
rect 24443 43605 24455 43639
rect 24397 43599 24455 43605
rect 24765 43639 24823 43645
rect 24765 43605 24777 43639
rect 24811 43605 24823 43639
rect 24765 43599 24823 43605
rect 24949 43639 25007 43645
rect 24949 43605 24961 43639
rect 24995 43636 25007 43639
rect 25130 43636 25136 43648
rect 24995 43608 25136 43636
rect 24995 43605 25007 43608
rect 24949 43599 25007 43605
rect 25130 43596 25136 43608
rect 25188 43596 25194 43648
rect 26418 43596 26424 43648
rect 26476 43636 26482 43648
rect 27249 43639 27307 43645
rect 27249 43636 27261 43639
rect 26476 43608 27261 43636
rect 26476 43596 26482 43608
rect 27249 43605 27261 43608
rect 27295 43605 27307 43639
rect 30006 43636 30012 43648
rect 29967 43608 30012 43636
rect 27249 43599 27307 43605
rect 30006 43596 30012 43608
rect 30064 43596 30070 43648
rect 1104 43546 30820 43568
rect 1104 43494 10880 43546
rect 10932 43494 10944 43546
rect 10996 43494 11008 43546
rect 11060 43494 11072 43546
rect 11124 43494 11136 43546
rect 11188 43494 20811 43546
rect 20863 43494 20875 43546
rect 20927 43494 20939 43546
rect 20991 43494 21003 43546
rect 21055 43494 21067 43546
rect 21119 43494 30820 43546
rect 1104 43472 30820 43494
rect 2409 43435 2467 43441
rect 2409 43432 2421 43435
rect 1688 43404 2421 43432
rect 1688 43376 1716 43404
rect 2409 43401 2421 43404
rect 2455 43401 2467 43435
rect 9582 43432 9588 43444
rect 9543 43404 9588 43432
rect 2409 43395 2467 43401
rect 9582 43392 9588 43404
rect 9640 43392 9646 43444
rect 9858 43432 9864 43444
rect 9856 43392 9864 43432
rect 9916 43392 9922 43444
rect 9950 43392 9956 43444
rect 10008 43392 10014 43444
rect 18138 43392 18144 43444
rect 18196 43432 18202 43444
rect 18325 43435 18383 43441
rect 18325 43432 18337 43435
rect 18196 43404 18337 43432
rect 18196 43392 18202 43404
rect 18325 43401 18337 43404
rect 18371 43401 18383 43435
rect 18325 43395 18383 43401
rect 19702 43392 19708 43444
rect 19760 43432 19766 43444
rect 20530 43432 20536 43444
rect 19760 43404 20536 43432
rect 19760 43392 19766 43404
rect 20530 43392 20536 43404
rect 20588 43432 20594 43444
rect 20809 43435 20867 43441
rect 20809 43432 20821 43435
rect 20588 43404 20821 43432
rect 20588 43392 20594 43404
rect 20809 43401 20821 43404
rect 20855 43401 20867 43435
rect 20809 43395 20867 43401
rect 23661 43435 23719 43441
rect 23661 43401 23673 43435
rect 23707 43432 23719 43435
rect 24578 43432 24584 43444
rect 23707 43404 24584 43432
rect 23707 43401 23719 43404
rect 23661 43395 23719 43401
rect 24578 43392 24584 43404
rect 24636 43392 24642 43444
rect 1581 43367 1639 43373
rect 1581 43333 1593 43367
rect 1627 43364 1639 43367
rect 1670 43364 1676 43376
rect 1627 43336 1676 43364
rect 1627 43333 1639 43336
rect 1581 43327 1639 43333
rect 1670 43324 1676 43336
rect 1728 43324 1734 43376
rect 1946 43324 1952 43376
rect 2004 43364 2010 43376
rect 9398 43364 9404 43376
rect 2004 43336 9404 43364
rect 2004 43324 2010 43336
rect 9398 43324 9404 43336
rect 9456 43324 9462 43376
rect 1762 43296 1768 43308
rect 1723 43268 1768 43296
rect 1762 43256 1768 43268
rect 1820 43256 1826 43308
rect 2222 43256 2228 43308
rect 2280 43296 2286 43308
rect 2498 43296 2504 43308
rect 2280 43268 2504 43296
rect 2280 43256 2286 43268
rect 2498 43256 2504 43268
rect 2556 43296 2562 43308
rect 9856 43305 9884 43392
rect 9968 43311 9996 43392
rect 12802 43364 12808 43376
rect 11808 43336 12808 43364
rect 9950 43305 10008 43311
rect 2593 43299 2651 43305
rect 2593 43296 2605 43299
rect 2556 43268 2605 43296
rect 2556 43256 2562 43268
rect 2593 43265 2605 43268
rect 2639 43265 2651 43299
rect 2593 43259 2651 43265
rect 9841 43299 9899 43305
rect 9841 43265 9853 43299
rect 9887 43265 9899 43299
rect 9950 43271 9962 43305
rect 9996 43271 10008 43305
rect 9950 43265 10008 43271
rect 9841 43259 9899 43265
rect 10042 43256 10048 43308
rect 10100 43296 10106 43308
rect 10226 43296 10232 43308
rect 10100 43268 10145 43296
rect 10187 43268 10232 43296
rect 10100 43256 10106 43268
rect 10226 43256 10232 43268
rect 10284 43256 10290 43308
rect 11808 43305 11836 43336
rect 12802 43324 12808 43336
rect 12860 43324 12866 43376
rect 14550 43324 14556 43376
rect 14608 43364 14614 43376
rect 15933 43367 15991 43373
rect 15933 43364 15945 43367
rect 14608 43336 15945 43364
rect 14608 43324 14614 43336
rect 15933 43333 15945 43336
rect 15979 43333 15991 43367
rect 15933 43327 15991 43333
rect 19521 43367 19579 43373
rect 19521 43333 19533 43367
rect 19567 43364 19579 43367
rect 19610 43364 19616 43376
rect 19567 43336 19616 43364
rect 19567 43333 19579 43336
rect 19521 43327 19579 43333
rect 19610 43324 19616 43336
rect 19668 43324 19674 43376
rect 22281 43367 22339 43373
rect 22281 43364 22293 43367
rect 21008 43336 22293 43364
rect 11793 43299 11851 43305
rect 11793 43265 11805 43299
rect 11839 43265 11851 43299
rect 13078 43296 13084 43308
rect 13039 43268 13084 43296
rect 11793 43259 11851 43265
rect 13078 43256 13084 43268
rect 13136 43256 13142 43308
rect 15010 43296 15016 43308
rect 14971 43268 15016 43296
rect 15010 43256 15016 43268
rect 15068 43256 15074 43308
rect 15470 43256 15476 43308
rect 15528 43296 15534 43308
rect 15749 43299 15807 43305
rect 15749 43296 15761 43299
rect 15528 43268 15761 43296
rect 15528 43256 15534 43268
rect 15749 43265 15761 43268
rect 15795 43296 15807 43299
rect 16298 43296 16304 43308
rect 15795 43268 16304 43296
rect 15795 43265 15807 43268
rect 15749 43259 15807 43265
rect 16298 43256 16304 43268
rect 16356 43256 16362 43308
rect 17034 43296 17040 43308
rect 16995 43268 17040 43296
rect 17034 43256 17040 43268
rect 17092 43256 17098 43308
rect 11517 43231 11575 43237
rect 11517 43197 11529 43231
rect 11563 43228 11575 43231
rect 12066 43228 12072 43240
rect 11563 43200 12072 43228
rect 11563 43197 11575 43200
rect 11517 43191 11575 43197
rect 12066 43188 12072 43200
rect 12124 43188 12130 43240
rect 12802 43228 12808 43240
rect 12763 43200 12808 43228
rect 12802 43188 12808 43200
rect 12860 43188 12866 43240
rect 13262 43188 13268 43240
rect 13320 43228 13326 43240
rect 13320 43200 17954 43228
rect 13320 43188 13326 43200
rect 1949 43163 2007 43169
rect 1949 43129 1961 43163
rect 1995 43160 2007 43163
rect 10318 43160 10324 43172
rect 1995 43132 10324 43160
rect 1995 43129 2007 43132
rect 1949 43123 2007 43129
rect 10318 43120 10324 43132
rect 10376 43120 10382 43172
rect 14274 43120 14280 43172
rect 14332 43160 14338 43172
rect 15194 43160 15200 43172
rect 14332 43132 15200 43160
rect 14332 43120 14338 43132
rect 15194 43120 15200 43132
rect 15252 43120 15258 43172
rect 17926 43160 17954 43200
rect 20622 43188 20628 43240
rect 20680 43228 20686 43240
rect 21008 43228 21036 43336
rect 22281 43333 22293 43336
rect 22327 43333 22339 43367
rect 22281 43327 22339 43333
rect 23753 43367 23811 43373
rect 23753 43333 23765 43367
rect 23799 43364 23811 43367
rect 25130 43364 25136 43376
rect 23799 43336 25136 43364
rect 23799 43333 23811 43336
rect 23753 43327 23811 43333
rect 25130 43324 25136 43336
rect 25188 43324 25194 43376
rect 29546 43324 29552 43376
rect 29604 43364 29610 43376
rect 29822 43364 29828 43376
rect 29604 43336 29828 43364
rect 29604 43324 29610 43336
rect 29822 43324 29828 43336
rect 29880 43324 29886 43376
rect 30098 43364 30104 43376
rect 30059 43336 30104 43364
rect 30098 43324 30104 43336
rect 30156 43324 30162 43376
rect 23477 43299 23535 43305
rect 23477 43265 23489 43299
rect 23523 43296 23535 43299
rect 23658 43296 23664 43308
rect 23523 43268 23664 43296
rect 23523 43265 23535 43268
rect 23477 43259 23535 43265
rect 23658 43256 23664 43268
rect 23716 43256 23722 43308
rect 23845 43299 23903 43305
rect 23845 43265 23857 43299
rect 23891 43296 23903 43299
rect 24581 43299 24639 43305
rect 24581 43296 24593 43299
rect 23891 43268 24593 43296
rect 23891 43265 23903 43268
rect 23845 43259 23903 43265
rect 24581 43265 24593 43268
rect 24627 43296 24639 43299
rect 24762 43296 24768 43308
rect 24627 43268 24768 43296
rect 24627 43265 24639 43268
rect 24581 43259 24639 43265
rect 24762 43256 24768 43268
rect 24820 43256 24826 43308
rect 25314 43256 25320 43308
rect 25372 43296 25378 43308
rect 25777 43299 25835 43305
rect 25777 43296 25789 43299
rect 25372 43268 25789 43296
rect 25372 43256 25378 43268
rect 25777 43265 25789 43268
rect 25823 43265 25835 43299
rect 25777 43259 25835 43265
rect 27985 43299 28043 43305
rect 27985 43265 27997 43299
rect 28031 43296 28043 43299
rect 28629 43299 28687 43305
rect 28031 43268 28580 43296
rect 28031 43265 28043 43268
rect 27985 43259 28043 43265
rect 20680 43200 21036 43228
rect 23385 43231 23443 43237
rect 20680 43188 20686 43200
rect 23385 43197 23397 43231
rect 23431 43228 23443 43231
rect 23431 43200 23704 43228
rect 23431 43197 23443 43200
rect 23385 43191 23443 43197
rect 23676 43172 23704 43200
rect 24026 43188 24032 43240
rect 24084 43228 24090 43240
rect 24305 43231 24363 43237
rect 24305 43228 24317 43231
rect 24084 43200 24317 43228
rect 24084 43188 24090 43200
rect 24305 43197 24317 43200
rect 24351 43228 24363 43231
rect 24486 43228 24492 43240
rect 24351 43200 24492 43228
rect 24351 43197 24363 43200
rect 24305 43191 24363 43197
rect 24486 43188 24492 43200
rect 24544 43188 24550 43240
rect 25961 43231 26019 43237
rect 25961 43228 25973 43231
rect 24596 43200 25973 43228
rect 24596 43172 24624 43200
rect 25961 43197 25973 43200
rect 26007 43197 26019 43231
rect 25961 43191 26019 43197
rect 17926 43132 23612 43160
rect 14090 43052 14096 43104
rect 14148 43092 14154 43104
rect 14369 43095 14427 43101
rect 14369 43092 14381 43095
rect 14148 43064 14381 43092
rect 14148 43052 14154 43064
rect 14369 43061 14381 43064
rect 14415 43092 14427 43095
rect 16206 43092 16212 43104
rect 14415 43064 16212 43092
rect 14415 43061 14427 43064
rect 14369 43055 14427 43061
rect 16206 43052 16212 43064
rect 16264 43052 16270 43104
rect 21358 43052 21364 43104
rect 21416 43092 21422 43104
rect 22370 43092 22376 43104
rect 21416 43064 22376 43092
rect 21416 43052 21422 43064
rect 22370 43052 22376 43064
rect 22428 43052 22434 43104
rect 23201 43095 23259 43101
rect 23201 43061 23213 43095
rect 23247 43092 23259 43095
rect 23290 43092 23296 43104
rect 23247 43064 23296 43092
rect 23247 43061 23259 43064
rect 23201 43055 23259 43061
rect 23290 43052 23296 43064
rect 23348 43052 23354 43104
rect 23584 43092 23612 43132
rect 23658 43120 23664 43172
rect 23716 43120 23722 43172
rect 24578 43120 24584 43172
rect 24636 43120 24642 43172
rect 25130 43120 25136 43172
rect 25188 43160 25194 43172
rect 25314 43160 25320 43172
rect 25188 43132 25320 43160
rect 25188 43120 25194 43132
rect 25314 43120 25320 43132
rect 25372 43120 25378 43172
rect 28552 43160 28580 43268
rect 28629 43265 28641 43299
rect 28675 43296 28687 43299
rect 29086 43296 29092 43308
rect 28675 43268 28994 43296
rect 29047 43268 29092 43296
rect 28675 43265 28687 43268
rect 28629 43259 28687 43265
rect 28966 43228 28994 43268
rect 29086 43256 29092 43268
rect 29144 43256 29150 43308
rect 29914 43296 29920 43308
rect 29875 43268 29920 43296
rect 29914 43256 29920 43268
rect 29972 43256 29978 43308
rect 30098 43228 30104 43240
rect 28966 43200 30104 43228
rect 30098 43188 30104 43200
rect 30156 43188 30162 43240
rect 28552 43132 29592 43160
rect 29564 43104 29592 43132
rect 24762 43092 24768 43104
rect 23584 43064 24768 43092
rect 24762 43052 24768 43064
rect 24820 43092 24826 43104
rect 26418 43092 26424 43104
rect 24820 43064 26424 43092
rect 24820 43052 24826 43064
rect 26418 43052 26424 43064
rect 26476 43052 26482 43104
rect 27798 43092 27804 43104
rect 27759 43064 27804 43092
rect 27798 43052 27804 43064
rect 27856 43052 27862 43104
rect 27982 43052 27988 43104
rect 28040 43092 28046 43104
rect 28445 43095 28503 43101
rect 28445 43092 28457 43095
rect 28040 43064 28457 43092
rect 28040 43052 28046 43064
rect 28445 43061 28457 43064
rect 28491 43061 28503 43095
rect 29270 43092 29276 43104
rect 29231 43064 29276 43092
rect 28445 43055 28503 43061
rect 29270 43052 29276 43064
rect 29328 43052 29334 43104
rect 29546 43052 29552 43104
rect 29604 43052 29610 43104
rect 1104 43002 30820 43024
rect 1104 42950 5915 43002
rect 5967 42950 5979 43002
rect 6031 42950 6043 43002
rect 6095 42950 6107 43002
rect 6159 42950 6171 43002
rect 6223 42950 15846 43002
rect 15898 42950 15910 43002
rect 15962 42950 15974 43002
rect 16026 42950 16038 43002
rect 16090 42950 16102 43002
rect 16154 42950 25776 43002
rect 25828 42950 25840 43002
rect 25892 42950 25904 43002
rect 25956 42950 25968 43002
rect 26020 42950 26032 43002
rect 26084 42950 30820 43002
rect 1104 42928 30820 42950
rect 1397 42891 1455 42897
rect 1397 42857 1409 42891
rect 1443 42888 1455 42891
rect 1762 42888 1768 42900
rect 1443 42860 1768 42888
rect 1443 42857 1455 42860
rect 1397 42851 1455 42857
rect 1762 42848 1768 42860
rect 1820 42848 1826 42900
rect 2041 42891 2099 42897
rect 2041 42857 2053 42891
rect 2087 42888 2099 42891
rect 2590 42888 2596 42900
rect 2087 42860 2596 42888
rect 2087 42857 2099 42860
rect 2041 42851 2099 42857
rect 2590 42848 2596 42860
rect 2648 42848 2654 42900
rect 12529 42891 12587 42897
rect 12529 42857 12541 42891
rect 12575 42888 12587 42891
rect 12802 42888 12808 42900
rect 12575 42860 12808 42888
rect 12575 42857 12587 42860
rect 12529 42851 12587 42857
rect 12802 42848 12808 42860
rect 12860 42848 12866 42900
rect 23658 42848 23664 42900
rect 23716 42888 23722 42900
rect 23716 42860 24624 42888
rect 23716 42848 23722 42860
rect 13998 42780 14004 42832
rect 14056 42820 14062 42832
rect 24596 42820 24624 42860
rect 24670 42848 24676 42900
rect 24728 42888 24734 42900
rect 27525 42891 27583 42897
rect 24728 42860 24900 42888
rect 24728 42848 24734 42860
rect 24762 42820 24768 42832
rect 14056 42792 16068 42820
rect 14056 42780 14062 42792
rect 9674 42752 9680 42764
rect 9508 42724 9680 42752
rect 1578 42684 1584 42696
rect 1539 42656 1584 42684
rect 1578 42644 1584 42656
rect 1636 42644 1642 42696
rect 2222 42684 2228 42696
rect 2183 42656 2228 42684
rect 2222 42644 2228 42656
rect 2280 42644 2286 42696
rect 9508 42693 9536 42724
rect 9674 42712 9680 42724
rect 9732 42712 9738 42764
rect 11514 42712 11520 42764
rect 11572 42752 11578 42764
rect 13265 42755 13323 42761
rect 13265 42752 13277 42755
rect 11572 42724 13277 42752
rect 11572 42712 11578 42724
rect 13265 42721 13277 42724
rect 13311 42721 13323 42755
rect 13265 42715 13323 42721
rect 14093 42755 14151 42761
rect 14093 42721 14105 42755
rect 14139 42752 14151 42755
rect 15010 42752 15016 42764
rect 14139 42724 15016 42752
rect 14139 42721 14151 42724
rect 14093 42715 14151 42721
rect 15010 42712 15016 42724
rect 15068 42712 15074 42764
rect 15194 42712 15200 42764
rect 15252 42752 15258 42764
rect 15252 42724 15792 42752
rect 15252 42712 15258 42724
rect 9493 42687 9551 42693
rect 9493 42653 9505 42687
rect 9539 42653 9551 42687
rect 10137 42687 10195 42693
rect 10137 42684 10149 42687
rect 9493 42647 9551 42653
rect 9692 42656 10149 42684
rect 9692 42557 9720 42656
rect 10137 42653 10149 42656
rect 10183 42653 10195 42687
rect 10410 42684 10416 42696
rect 10371 42656 10416 42684
rect 10137 42647 10195 42653
rect 10410 42644 10416 42656
rect 10468 42644 10474 42696
rect 12345 42687 12403 42693
rect 12345 42653 12357 42687
rect 12391 42653 12403 42687
rect 14366 42684 14372 42696
rect 14327 42656 14372 42684
rect 12345 42647 12403 42653
rect 11793 42619 11851 42625
rect 11793 42585 11805 42619
rect 11839 42616 11851 42619
rect 11974 42616 11980 42628
rect 11839 42588 11980 42616
rect 11839 42585 11851 42588
rect 11793 42579 11851 42585
rect 11974 42576 11980 42588
rect 12032 42576 12038 42628
rect 9677 42551 9735 42557
rect 9677 42517 9689 42551
rect 9723 42517 9735 42551
rect 12360 42548 12388 42647
rect 14366 42644 14372 42656
rect 14424 42644 14430 42696
rect 15470 42684 15476 42696
rect 14936 42656 15476 42684
rect 13081 42619 13139 42625
rect 13081 42585 13093 42619
rect 13127 42616 13139 42619
rect 14936 42616 14964 42656
rect 15470 42644 15476 42656
rect 15528 42644 15534 42696
rect 15654 42684 15660 42696
rect 15615 42656 15660 42684
rect 15654 42644 15660 42656
rect 15712 42644 15718 42696
rect 15764 42693 15792 42724
rect 16040 42693 16068 42792
rect 24596 42792 24768 42820
rect 17126 42712 17132 42764
rect 17184 42752 17190 42764
rect 19521 42755 19579 42761
rect 19521 42752 19533 42755
rect 17184 42724 19533 42752
rect 17184 42712 17190 42724
rect 19521 42721 19533 42724
rect 19567 42721 19579 42755
rect 21910 42752 21916 42764
rect 21871 42724 21916 42752
rect 19521 42715 19579 42721
rect 21910 42712 21916 42724
rect 21968 42712 21974 42764
rect 23290 42712 23296 42764
rect 23348 42752 23354 42764
rect 24486 42752 24492 42764
rect 23348 42724 24492 42752
rect 23348 42712 23354 42724
rect 24486 42712 24492 42724
rect 24544 42712 24550 42764
rect 24596 42761 24624 42792
rect 24762 42780 24768 42792
rect 24820 42780 24826 42832
rect 24581 42755 24639 42761
rect 24581 42721 24593 42755
rect 24627 42721 24639 42755
rect 24581 42715 24639 42721
rect 15749 42687 15807 42693
rect 15749 42653 15761 42687
rect 15795 42653 15807 42687
rect 15749 42647 15807 42653
rect 15841 42687 15899 42693
rect 15841 42653 15853 42687
rect 15887 42653 15899 42687
rect 15841 42647 15899 42653
rect 16025 42687 16083 42693
rect 16025 42653 16037 42687
rect 16071 42653 16083 42687
rect 16025 42647 16083 42653
rect 13127 42588 14964 42616
rect 13127 42585 13139 42588
rect 13081 42579 13139 42585
rect 15102 42576 15108 42628
rect 15160 42616 15166 42628
rect 15856 42616 15884 42647
rect 18414 42644 18420 42696
rect 18472 42684 18478 42696
rect 19337 42687 19395 42693
rect 19337 42684 19349 42687
rect 18472 42656 19349 42684
rect 18472 42644 18478 42656
rect 19337 42653 19349 42656
rect 19383 42653 19395 42687
rect 19337 42647 19395 42653
rect 20070 42644 20076 42696
rect 20128 42684 20134 42696
rect 20257 42687 20315 42693
rect 20257 42684 20269 42687
rect 20128 42656 20269 42684
rect 20128 42644 20134 42656
rect 20257 42653 20269 42656
rect 20303 42653 20315 42687
rect 20257 42647 20315 42653
rect 22278 42644 22284 42696
rect 22336 42684 22342 42696
rect 22465 42687 22523 42693
rect 22465 42684 22477 42687
rect 22336 42656 22477 42684
rect 22336 42644 22342 42656
rect 22465 42653 22477 42656
rect 22511 42653 22523 42687
rect 22465 42647 22523 42653
rect 24673 42687 24731 42693
rect 24673 42653 24685 42687
rect 24719 42684 24731 42687
rect 24872 42684 24900 42860
rect 27525 42857 27537 42891
rect 27571 42888 27583 42891
rect 28258 42888 28264 42900
rect 27571 42860 28264 42888
rect 27571 42857 27583 42860
rect 27525 42851 27583 42857
rect 28258 42848 28264 42860
rect 28316 42888 28322 42900
rect 28626 42888 28632 42900
rect 28316 42860 28632 42888
rect 28316 42848 28322 42860
rect 28626 42848 28632 42860
rect 28684 42848 28690 42900
rect 29822 42848 29828 42900
rect 29880 42888 29886 42900
rect 29880 42860 31524 42888
rect 29880 42848 29886 42860
rect 25130 42780 25136 42832
rect 25188 42780 25194 42832
rect 27586 42792 30236 42820
rect 25148 42752 25176 42780
rect 25056 42724 25176 42752
rect 25056 42693 25084 42724
rect 25774 42712 25780 42764
rect 25832 42752 25838 42764
rect 27586 42752 27614 42792
rect 28902 42752 28908 42764
rect 25832 42724 27614 42752
rect 28644 42724 28908 42752
rect 25832 42712 25838 42724
rect 24719 42656 24900 42684
rect 25041 42687 25099 42693
rect 24719 42653 24731 42656
rect 24673 42647 24731 42653
rect 25041 42653 25053 42687
rect 25087 42653 25099 42687
rect 25041 42647 25099 42653
rect 25130 42644 25136 42696
rect 25188 42684 25194 42696
rect 25188 42656 26004 42684
rect 25188 42644 25194 42656
rect 15160 42588 15884 42616
rect 16945 42619 17003 42625
rect 15160 42576 15166 42588
rect 16945 42585 16957 42619
rect 16991 42616 17003 42619
rect 18598 42616 18604 42628
rect 16991 42588 18604 42616
rect 16991 42585 17003 42588
rect 16945 42579 17003 42585
rect 18598 42576 18604 42588
rect 18656 42576 18662 42628
rect 24397 42619 24455 42625
rect 24397 42585 24409 42619
rect 24443 42616 24455 42619
rect 25682 42616 25688 42628
rect 24443 42588 25688 42616
rect 24443 42585 24455 42588
rect 24397 42579 24455 42585
rect 25682 42576 25688 42588
rect 25740 42576 25746 42628
rect 25866 42616 25872 42628
rect 25827 42588 25872 42616
rect 25866 42576 25872 42588
rect 25924 42576 25930 42628
rect 25976 42616 26004 42656
rect 26234 42644 26240 42696
rect 26292 42684 26298 42696
rect 26789 42687 26847 42693
rect 26789 42684 26801 42687
rect 26292 42656 26801 42684
rect 26292 42644 26298 42656
rect 26789 42653 26801 42656
rect 26835 42653 26847 42687
rect 26789 42647 26847 42653
rect 28258 42644 28264 42696
rect 28316 42684 28322 42696
rect 28644 42694 28672 42724
rect 28902 42712 28908 42724
rect 28960 42752 28966 42764
rect 28960 42724 29776 42752
rect 28960 42712 28966 42724
rect 28644 42693 28764 42694
rect 29748 42693 29776 42724
rect 28644 42687 28779 42693
rect 28316 42656 28580 42684
rect 28644 42666 28733 42687
rect 28316 42644 28322 42656
rect 26605 42619 26663 42625
rect 26605 42616 26617 42619
rect 25976 42588 26617 42616
rect 26605 42585 26617 42588
rect 26651 42585 26663 42619
rect 26605 42579 26663 42585
rect 27433 42619 27491 42625
rect 27433 42585 27445 42619
rect 27479 42616 27491 42619
rect 28350 42616 28356 42628
rect 27479 42588 28356 42616
rect 27479 42585 27491 42588
rect 27433 42579 27491 42585
rect 12986 42548 12992 42560
rect 12360 42520 12992 42548
rect 9677 42511 9735 42517
rect 12986 42508 12992 42520
rect 13044 42508 13050 42560
rect 15378 42548 15384 42560
rect 15339 42520 15384 42548
rect 15378 42508 15384 42520
rect 15436 42508 15442 42560
rect 16390 42508 16396 42560
rect 16448 42548 16454 42560
rect 18230 42548 18236 42560
rect 16448 42520 18236 42548
rect 16448 42508 16454 42520
rect 18230 42508 18236 42520
rect 18288 42508 18294 42560
rect 18966 42508 18972 42560
rect 19024 42548 19030 42560
rect 22278 42548 22284 42560
rect 19024 42520 22284 42548
rect 19024 42508 19030 42520
rect 22278 42508 22284 42520
rect 22336 42508 22342 42560
rect 22646 42548 22652 42560
rect 22607 42520 22652 42548
rect 22646 42508 22652 42520
rect 22704 42508 22710 42560
rect 24670 42508 24676 42560
rect 24728 42548 24734 42560
rect 24765 42551 24823 42557
rect 24765 42548 24777 42551
rect 24728 42520 24777 42548
rect 24728 42508 24734 42520
rect 24765 42517 24777 42520
rect 24811 42517 24823 42551
rect 24765 42511 24823 42517
rect 24949 42551 25007 42557
rect 24949 42517 24961 42551
rect 24995 42548 25007 42551
rect 25314 42548 25320 42560
rect 24995 42520 25320 42548
rect 24995 42517 25007 42520
rect 24949 42511 25007 42517
rect 25314 42508 25320 42520
rect 25372 42508 25378 42560
rect 25958 42548 25964 42560
rect 25919 42520 25964 42548
rect 25958 42508 25964 42520
rect 26016 42508 26022 42560
rect 26050 42508 26056 42560
rect 26108 42548 26114 42560
rect 27448 42548 27476 42579
rect 28350 42576 28356 42588
rect 28408 42576 28414 42628
rect 28552 42616 28580 42656
rect 28721 42653 28733 42666
rect 28767 42653 28779 42687
rect 28721 42647 28779 42653
rect 28997 42687 29055 42693
rect 28997 42653 29009 42687
rect 29043 42653 29055 42687
rect 28997 42647 29055 42653
rect 29733 42687 29791 42693
rect 29733 42653 29745 42687
rect 29779 42653 29791 42687
rect 29733 42647 29791 42653
rect 30009 42687 30067 42693
rect 30009 42653 30021 42687
rect 30055 42653 30067 42687
rect 30009 42647 30067 42653
rect 29012 42616 29040 42647
rect 30024 42616 30052 42647
rect 28552 42588 30052 42616
rect 29748 42560 29776 42588
rect 26108 42520 27476 42548
rect 28537 42551 28595 42557
rect 26108 42508 26114 42520
rect 28537 42517 28549 42551
rect 28583 42548 28595 42551
rect 28810 42548 28816 42560
rect 28583 42520 28816 42548
rect 28583 42517 28595 42520
rect 28537 42511 28595 42517
rect 28810 42508 28816 42520
rect 28868 42508 28874 42560
rect 28905 42551 28963 42557
rect 28905 42517 28917 42551
rect 28951 42548 28963 42551
rect 28994 42548 29000 42560
rect 28951 42520 29000 42548
rect 28951 42517 28963 42520
rect 28905 42511 28963 42517
rect 28994 42508 29000 42520
rect 29052 42508 29058 42560
rect 29549 42551 29607 42557
rect 29549 42517 29561 42551
rect 29595 42548 29607 42551
rect 29638 42548 29644 42560
rect 29595 42520 29644 42548
rect 29595 42517 29607 42520
rect 29549 42511 29607 42517
rect 29638 42508 29644 42520
rect 29696 42508 29702 42560
rect 29730 42508 29736 42560
rect 29788 42508 29794 42560
rect 29917 42551 29975 42557
rect 29917 42517 29929 42551
rect 29963 42548 29975 42551
rect 30208 42548 30236 42792
rect 29963 42520 30236 42548
rect 29963 42517 29975 42520
rect 29917 42511 29975 42517
rect 1104 42458 30820 42480
rect 1104 42406 10880 42458
rect 10932 42406 10944 42458
rect 10996 42406 11008 42458
rect 11060 42406 11072 42458
rect 11124 42406 11136 42458
rect 11188 42406 20811 42458
rect 20863 42406 20875 42458
rect 20927 42406 20939 42458
rect 20991 42406 21003 42458
rect 21055 42406 21067 42458
rect 21119 42406 30820 42458
rect 1104 42384 30820 42406
rect 1397 42347 1455 42353
rect 1397 42313 1409 42347
rect 1443 42344 1455 42347
rect 9677 42347 9735 42353
rect 1443 42316 2774 42344
rect 1443 42313 1455 42316
rect 1397 42307 1455 42313
rect 2746 42276 2774 42316
rect 9677 42313 9689 42347
rect 9723 42344 9735 42347
rect 10410 42344 10416 42356
rect 9723 42316 10416 42344
rect 9723 42313 9735 42316
rect 9677 42307 9735 42313
rect 10410 42304 10416 42316
rect 10468 42304 10474 42356
rect 11882 42304 11888 42356
rect 11940 42344 11946 42356
rect 12161 42347 12219 42353
rect 12161 42344 12173 42347
rect 11940 42316 12173 42344
rect 11940 42304 11946 42316
rect 12161 42313 12173 42316
rect 12207 42313 12219 42347
rect 12161 42307 12219 42313
rect 14553 42347 14611 42353
rect 14553 42313 14565 42347
rect 14599 42344 14611 42347
rect 14642 42344 14648 42356
rect 14599 42316 14648 42344
rect 14599 42313 14611 42316
rect 14553 42307 14611 42313
rect 14642 42304 14648 42316
rect 14700 42304 14706 42356
rect 15102 42304 15108 42356
rect 15160 42344 15166 42356
rect 15381 42347 15439 42353
rect 15381 42344 15393 42347
rect 15160 42316 15393 42344
rect 15160 42304 15166 42316
rect 15381 42313 15393 42316
rect 15427 42313 15439 42347
rect 15381 42307 15439 42313
rect 16117 42347 16175 42353
rect 16117 42313 16129 42347
rect 16163 42344 16175 42347
rect 17034 42344 17040 42356
rect 16163 42316 17040 42344
rect 16163 42313 16175 42316
rect 16117 42307 16175 42313
rect 17034 42304 17040 42316
rect 17092 42304 17098 42356
rect 19242 42304 19248 42356
rect 19300 42344 19306 42356
rect 20073 42347 20131 42353
rect 20073 42344 20085 42347
rect 19300 42316 20085 42344
rect 19300 42304 19306 42316
rect 20073 42313 20085 42316
rect 20119 42313 20131 42347
rect 20073 42307 20131 42313
rect 21358 42304 21364 42356
rect 21416 42344 21422 42356
rect 23290 42344 23296 42356
rect 21416 42316 23296 42344
rect 21416 42304 21422 42316
rect 23290 42304 23296 42316
rect 23348 42344 23354 42356
rect 23477 42347 23535 42353
rect 23477 42344 23489 42347
rect 23348 42316 23489 42344
rect 23348 42304 23354 42316
rect 23477 42313 23489 42316
rect 23523 42313 23535 42347
rect 23477 42307 23535 42313
rect 25774 42304 25780 42356
rect 25832 42344 25838 42356
rect 27183 42347 27241 42353
rect 25832 42316 27108 42344
rect 25832 42304 25838 42316
rect 8573 42279 8631 42285
rect 8573 42276 8585 42279
rect 2746 42248 8585 42276
rect 8573 42245 8585 42248
rect 8619 42245 8631 42279
rect 8573 42239 8631 42245
rect 8757 42279 8815 42285
rect 8757 42245 8769 42279
rect 8803 42276 8815 42279
rect 13541 42279 13599 42285
rect 8803 42248 10272 42276
rect 8803 42245 8815 42248
rect 8757 42239 8815 42245
rect 10244 42220 10272 42248
rect 13541 42245 13553 42279
rect 13587 42276 13599 42279
rect 14369 42279 14427 42285
rect 14369 42276 14381 42279
rect 13587 42248 14381 42276
rect 13587 42245 13599 42248
rect 13541 42239 13599 42245
rect 14369 42245 14381 42248
rect 14415 42276 14427 42279
rect 14458 42276 14464 42288
rect 14415 42248 14464 42276
rect 14415 42245 14427 42248
rect 14369 42239 14427 42245
rect 14458 42236 14464 42248
rect 14516 42236 14522 42288
rect 15746 42276 15752 42288
rect 15212 42248 15752 42276
rect 1578 42208 1584 42220
rect 1539 42180 1584 42208
rect 1578 42168 1584 42180
rect 1636 42168 1642 42220
rect 8386 42208 8392 42220
rect 8347 42180 8392 42208
rect 8386 42168 8392 42180
rect 8444 42168 8450 42220
rect 9933 42211 9991 42217
rect 9933 42208 9945 42211
rect 9856 42180 9945 42208
rect 9856 42004 9884 42180
rect 9933 42177 9945 42180
rect 9979 42177 9991 42211
rect 9933 42171 9991 42177
rect 10026 42211 10084 42217
rect 10026 42177 10038 42211
rect 10072 42177 10084 42211
rect 10026 42171 10084 42177
rect 10137 42211 10195 42217
rect 10137 42177 10149 42211
rect 10183 42177 10195 42211
rect 10137 42171 10195 42177
rect 10041 42140 10069 42171
rect 9959 42112 10069 42140
rect 9959 42084 9987 42112
rect 9950 42032 9956 42084
rect 10008 42032 10014 42084
rect 10042 42032 10048 42084
rect 10100 42072 10106 42084
rect 10152 42072 10180 42171
rect 10226 42168 10232 42220
rect 10284 42168 10290 42220
rect 10321 42211 10379 42217
rect 10321 42177 10333 42211
rect 10367 42177 10379 42211
rect 10321 42171 10379 42177
rect 11977 42211 12035 42217
rect 11977 42177 11989 42211
rect 12023 42208 12035 42211
rect 13357 42211 13415 42217
rect 12023 42180 12434 42208
rect 12023 42177 12035 42180
rect 11977 42171 12035 42177
rect 10336 42084 10364 42171
rect 12406 42140 12434 42180
rect 13357 42177 13369 42211
rect 13403 42208 13415 42211
rect 15212 42208 15240 42248
rect 15746 42236 15752 42248
rect 15804 42236 15810 42288
rect 16761 42279 16819 42285
rect 16761 42245 16773 42279
rect 16807 42276 16819 42279
rect 16942 42276 16948 42288
rect 16807 42248 16948 42276
rect 16807 42245 16819 42248
rect 16761 42239 16819 42245
rect 16942 42236 16948 42248
rect 17000 42236 17006 42288
rect 22094 42276 22100 42288
rect 19260 42248 20116 42276
rect 13403 42180 15240 42208
rect 15289 42211 15347 42217
rect 13403 42177 13415 42180
rect 13357 42171 13415 42177
rect 15289 42177 15301 42211
rect 15335 42177 15347 42211
rect 15289 42171 15347 42177
rect 15933 42211 15991 42217
rect 15933 42177 15945 42211
rect 15979 42208 15991 42211
rect 16666 42208 16672 42220
rect 15979 42180 16672 42208
rect 15979 42177 15991 42180
rect 15933 42171 15991 42177
rect 14274 42140 14280 42152
rect 12406 42112 14280 42140
rect 14274 42100 14280 42112
rect 14332 42100 14338 42152
rect 14550 42100 14556 42152
rect 14608 42140 14614 42152
rect 14645 42143 14703 42149
rect 14645 42140 14657 42143
rect 14608 42112 14657 42140
rect 14608 42100 14614 42112
rect 14645 42109 14657 42112
rect 14691 42109 14703 42143
rect 14645 42103 14703 42109
rect 15304 42140 15332 42171
rect 16666 42168 16672 42180
rect 16724 42168 16730 42220
rect 17678 42217 17684 42220
rect 17672 42208 17684 42217
rect 17639 42180 17684 42208
rect 17672 42171 17684 42180
rect 17678 42168 17684 42171
rect 17736 42168 17742 42220
rect 19260 42217 19288 42248
rect 20088 42220 20116 42248
rect 20456 42248 22100 42276
rect 19245 42211 19303 42217
rect 19245 42177 19257 42211
rect 19291 42177 19303 42211
rect 19245 42171 19303 42177
rect 19337 42211 19395 42217
rect 19337 42177 19349 42211
rect 19383 42208 19395 42211
rect 19889 42211 19947 42217
rect 19889 42208 19901 42211
rect 19383 42180 19901 42208
rect 19383 42177 19395 42180
rect 19337 42171 19395 42177
rect 19889 42177 19901 42180
rect 19935 42177 19947 42211
rect 19889 42171 19947 42177
rect 20070 42168 20076 42220
rect 20128 42168 20134 42220
rect 20456 42208 20484 42248
rect 22094 42236 22100 42248
rect 22152 42236 22158 42288
rect 22186 42236 22192 42288
rect 22244 42276 22250 42288
rect 22342 42279 22400 42285
rect 22342 42276 22354 42279
rect 22244 42248 22354 42276
rect 22244 42236 22250 42248
rect 22342 42245 22354 42248
rect 22388 42245 22400 42279
rect 26234 42276 26240 42288
rect 22342 42239 22400 42245
rect 24136 42248 26240 42276
rect 20180 42180 20484 42208
rect 20533 42211 20591 42217
rect 16850 42140 16856 42152
rect 15304 42112 16856 42140
rect 10100 42044 10180 42072
rect 10100 42032 10106 42044
rect 10318 42032 10324 42084
rect 10376 42032 10382 42084
rect 12066 42032 12072 42084
rect 12124 42072 12130 42084
rect 15304 42072 15332 42112
rect 16850 42100 16856 42112
rect 16908 42100 16914 42152
rect 17402 42140 17408 42152
rect 17363 42112 17408 42140
rect 17402 42100 17408 42112
rect 17460 42100 17466 42152
rect 18874 42100 18880 42152
rect 18932 42140 18938 42152
rect 20180 42140 20208 42180
rect 20533 42177 20545 42211
rect 20579 42208 20591 42211
rect 20622 42208 20628 42220
rect 20579 42180 20628 42208
rect 20579 42177 20591 42180
rect 20533 42171 20591 42177
rect 20622 42168 20628 42180
rect 20680 42168 20686 42220
rect 24136 42208 24164 42248
rect 26234 42236 26240 42248
rect 26292 42236 26298 42288
rect 26418 42236 26424 42288
rect 26476 42276 26482 42288
rect 26973 42279 27031 42285
rect 26973 42276 26985 42279
rect 26476 42248 26985 42276
rect 26476 42236 26482 42248
rect 26973 42245 26985 42248
rect 27019 42245 27031 42279
rect 27080 42276 27108 42316
rect 27183 42313 27195 42347
rect 27229 42344 27241 42347
rect 27982 42344 27988 42356
rect 27229 42316 27988 42344
rect 27229 42313 27241 42316
rect 27183 42307 27241 42313
rect 27724 42288 27752 42316
rect 27982 42304 27988 42316
rect 28040 42304 28046 42356
rect 29638 42304 29644 42356
rect 29696 42304 29702 42356
rect 29730 42304 29736 42356
rect 29788 42344 29794 42356
rect 30098 42344 30104 42356
rect 29788 42316 30104 42344
rect 29788 42304 29794 42316
rect 30098 42304 30104 42316
rect 30156 42304 30162 42356
rect 31386 42344 31392 42356
rect 30392 42316 31392 42344
rect 27430 42276 27436 42288
rect 27080 42248 27436 42276
rect 26973 42239 27031 42245
rect 27430 42236 27436 42248
rect 27488 42236 27494 42288
rect 27706 42236 27712 42288
rect 27764 42236 27770 42288
rect 28350 42276 28356 42288
rect 28184 42248 28356 42276
rect 20732 42180 24164 42208
rect 24857 42211 24915 42217
rect 20732 42140 20760 42180
rect 24857 42177 24869 42211
rect 24903 42208 24915 42211
rect 25406 42208 25412 42220
rect 24903 42180 25412 42208
rect 24903 42177 24915 42180
rect 24857 42171 24915 42177
rect 25406 42168 25412 42180
rect 25464 42168 25470 42220
rect 26053 42211 26111 42217
rect 26053 42177 26065 42211
rect 26099 42208 26111 42211
rect 26510 42208 26516 42220
rect 26099 42180 26516 42208
rect 26099 42177 26111 42180
rect 26053 42171 26111 42177
rect 26510 42168 26516 42180
rect 26568 42168 26574 42220
rect 27798 42208 27804 42220
rect 27172 42180 27804 42208
rect 18932 42112 20208 42140
rect 20272 42112 20760 42140
rect 22097 42143 22155 42149
rect 18932 42100 18938 42112
rect 12124 42044 15332 42072
rect 16945 42075 17003 42081
rect 12124 42032 12130 42044
rect 16945 42041 16957 42075
rect 16991 42072 17003 42075
rect 17126 42072 17132 42084
rect 16991 42044 17132 42072
rect 16991 42041 17003 42044
rect 16945 42035 17003 42041
rect 17126 42032 17132 42044
rect 17184 42032 17190 42084
rect 18782 42072 18788 42084
rect 18695 42044 18788 42072
rect 18782 42032 18788 42044
rect 18840 42072 18846 42084
rect 20272 42072 20300 42112
rect 22097 42109 22109 42143
rect 22143 42109 22155 42143
rect 25774 42140 25780 42152
rect 22097 42103 22155 42109
rect 23124 42112 25780 42140
rect 18840 42044 20300 42072
rect 20717 42075 20775 42081
rect 18840 42032 18846 42044
rect 20717 42041 20729 42075
rect 20763 42072 20775 42075
rect 22112 42072 22140 42103
rect 20763 42044 22140 42072
rect 20763 42041 20775 42044
rect 20717 42035 20775 42041
rect 11974 42004 11980 42016
rect 9856 41976 11980 42004
rect 11974 41964 11980 41976
rect 12032 41964 12038 42016
rect 14090 42004 14096 42016
rect 14051 41976 14096 42004
rect 14090 41964 14096 41976
rect 14148 41964 14154 42016
rect 16666 41964 16672 42016
rect 16724 42004 16730 42016
rect 18506 42004 18512 42016
rect 16724 41976 18512 42004
rect 16724 41964 16730 41976
rect 18506 41964 18512 41976
rect 18564 41964 18570 42016
rect 19518 41964 19524 42016
rect 19576 42004 19582 42016
rect 20254 42004 20260 42016
rect 19576 41976 20260 42004
rect 19576 41964 19582 41976
rect 20254 41964 20260 41976
rect 20312 41964 20318 42016
rect 21450 41964 21456 42016
rect 21508 42004 21514 42016
rect 23124 42004 23152 42112
rect 25774 42100 25780 42112
rect 25832 42100 25838 42152
rect 24762 42032 24768 42084
rect 24820 42072 24826 42084
rect 25958 42072 25964 42084
rect 24820 42044 25964 42072
rect 24820 42032 24826 42044
rect 25958 42032 25964 42044
rect 26016 42032 26022 42084
rect 26050 42032 26056 42084
rect 26108 42032 26114 42084
rect 26237 42075 26295 42081
rect 26237 42041 26249 42075
rect 26283 42072 26295 42075
rect 26326 42072 26332 42084
rect 26283 42044 26332 42072
rect 26283 42041 26295 42044
rect 26237 42035 26295 42041
rect 26326 42032 26332 42044
rect 26384 42072 26390 42084
rect 26694 42072 26700 42084
rect 26384 42044 26700 42072
rect 26384 42032 26390 42044
rect 26694 42032 26700 42044
rect 26752 42032 26758 42084
rect 27172 42072 27200 42180
rect 27798 42168 27804 42180
rect 27856 42168 27862 42220
rect 28184 42217 28212 42248
rect 28350 42236 28356 42248
rect 28408 42276 28414 42288
rect 28902 42276 28908 42288
rect 28408 42248 28908 42276
rect 28408 42236 28414 42248
rect 28902 42236 28908 42248
rect 28960 42236 28966 42288
rect 29656 42276 29684 42304
rect 29656 42248 30144 42276
rect 28169 42211 28227 42217
rect 28169 42177 28181 42211
rect 28215 42177 28227 42211
rect 28169 42171 28227 42177
rect 28258 42168 28264 42220
rect 28316 42208 28322 42220
rect 28445 42211 28503 42217
rect 28445 42208 28457 42211
rect 28316 42180 28457 42208
rect 28316 42168 28322 42180
rect 28445 42177 28457 42180
rect 28491 42177 28503 42211
rect 28445 42171 28503 42177
rect 28534 42168 28540 42220
rect 28592 42208 28598 42220
rect 29733 42211 29791 42217
rect 29733 42208 29745 42211
rect 28592 42180 29745 42208
rect 28592 42168 28598 42180
rect 29733 42177 29745 42180
rect 29779 42177 29791 42211
rect 29733 42171 29791 42177
rect 29825 42211 29883 42217
rect 29825 42177 29837 42211
rect 29871 42177 29883 42211
rect 29825 42171 29883 42177
rect 27430 42100 27436 42152
rect 27488 42140 27494 42152
rect 29840 42140 29868 42171
rect 29914 42168 29920 42220
rect 29972 42208 29978 42220
rect 30116 42217 30144 42248
rect 30101 42211 30159 42217
rect 29972 42180 30017 42208
rect 29972 42168 29978 42180
rect 30101 42177 30113 42211
rect 30147 42177 30159 42211
rect 30101 42171 30159 42177
rect 30392 42140 30420 42316
rect 31386 42304 31392 42316
rect 31444 42304 31450 42356
rect 30650 42236 30656 42288
rect 30708 42276 30714 42288
rect 31496 42276 31524 42860
rect 30708 42248 31340 42276
rect 30708 42236 30714 42248
rect 30466 42168 30472 42220
rect 30524 42168 30530 42220
rect 27488 42112 29592 42140
rect 29840 42112 30420 42140
rect 27488 42100 27494 42112
rect 27172 42044 27580 42072
rect 21508 41976 23152 42004
rect 21508 41964 21514 41976
rect 24670 41964 24676 42016
rect 24728 42004 24734 42016
rect 24949 42007 25007 42013
rect 24949 42004 24961 42007
rect 24728 41976 24961 42004
rect 24728 41964 24734 41976
rect 24949 41973 24961 41976
rect 24995 41973 25007 42007
rect 24949 41967 25007 41973
rect 25314 41964 25320 42016
rect 25372 42004 25378 42016
rect 26068 42004 26096 42032
rect 27172 42013 27200 42044
rect 25372 41976 26096 42004
rect 27157 42007 27215 42013
rect 25372 41964 25378 41976
rect 27157 41973 27169 42007
rect 27203 41973 27215 42007
rect 27157 41967 27215 41973
rect 27341 42007 27399 42013
rect 27341 41973 27353 42007
rect 27387 42004 27399 42007
rect 27430 42004 27436 42016
rect 27387 41976 27436 42004
rect 27387 41973 27399 41976
rect 27341 41967 27399 41973
rect 27430 41964 27436 41976
rect 27488 41964 27494 42016
rect 27552 42004 27580 42044
rect 27614 42032 27620 42084
rect 27672 42072 27678 42084
rect 28350 42072 28356 42084
rect 27672 42044 28356 42072
rect 27672 42032 27678 42044
rect 28350 42032 28356 42044
rect 28408 42072 28414 42084
rect 29086 42072 29092 42084
rect 28408 42044 29092 42072
rect 28408 42032 28414 42044
rect 29086 42032 29092 42044
rect 29144 42032 29150 42084
rect 27982 42004 27988 42016
rect 27552 41976 27988 42004
rect 27982 41964 27988 41976
rect 28040 41964 28046 42016
rect 29454 42004 29460 42016
rect 29415 41976 29460 42004
rect 29454 41964 29460 41976
rect 29512 41964 29518 42016
rect 29564 42004 29592 42112
rect 29638 42032 29644 42084
rect 29696 42072 29702 42084
rect 29914 42072 29920 42084
rect 29696 42044 29920 42072
rect 29696 42032 29702 42044
rect 29914 42032 29920 42044
rect 29972 42032 29978 42084
rect 30484 42072 30512 42168
rect 30484 42044 30880 42072
rect 30006 42004 30012 42016
rect 29564 41976 30012 42004
rect 30006 41964 30012 41976
rect 30064 41964 30070 42016
rect 1104 41914 30820 41936
rect 1104 41862 5915 41914
rect 5967 41862 5979 41914
rect 6031 41862 6043 41914
rect 6095 41862 6107 41914
rect 6159 41862 6171 41914
rect 6223 41862 15846 41914
rect 15898 41862 15910 41914
rect 15962 41862 15974 41914
rect 16026 41862 16038 41914
rect 16090 41862 16102 41914
rect 16154 41862 25776 41914
rect 25828 41862 25840 41914
rect 25892 41862 25904 41914
rect 25956 41862 25968 41914
rect 26020 41862 26032 41914
rect 26084 41862 30820 41914
rect 1104 41840 30820 41862
rect 9309 41803 9367 41809
rect 9309 41769 9321 41803
rect 9355 41800 9367 41803
rect 10318 41800 10324 41812
rect 9355 41772 10324 41800
rect 9355 41769 9367 41772
rect 9309 41763 9367 41769
rect 10318 41760 10324 41772
rect 10376 41760 10382 41812
rect 12894 41760 12900 41812
rect 12952 41800 12958 41812
rect 12989 41803 13047 41809
rect 12989 41800 13001 41803
rect 12952 41772 13001 41800
rect 12952 41760 12958 41772
rect 12989 41769 13001 41772
rect 13035 41769 13047 41803
rect 12989 41763 13047 41769
rect 15654 41760 15660 41812
rect 15712 41800 15718 41812
rect 15712 41772 16160 41800
rect 15712 41760 15718 41772
rect 16132 41741 16160 41772
rect 17218 41760 17224 41812
rect 17276 41800 17282 41812
rect 17681 41803 17739 41809
rect 17681 41800 17693 41803
rect 17276 41772 17693 41800
rect 17276 41760 17282 41772
rect 17681 41769 17693 41772
rect 17727 41769 17739 41803
rect 19429 41803 19487 41809
rect 17681 41763 17739 41769
rect 17972 41772 18644 41800
rect 14277 41735 14335 41741
rect 14277 41701 14289 41735
rect 14323 41701 14335 41735
rect 14277 41695 14335 41701
rect 16117 41735 16175 41741
rect 16117 41701 16129 41735
rect 16163 41732 16175 41735
rect 17972 41732 18000 41772
rect 18506 41732 18512 41744
rect 16163 41704 18000 41732
rect 18467 41704 18512 41732
rect 16163 41701 16175 41704
rect 16117 41695 16175 41701
rect 10413 41667 10471 41673
rect 10413 41633 10425 41667
rect 10459 41664 10471 41667
rect 12066 41664 12072 41676
rect 10459 41636 12072 41664
rect 10459 41633 10471 41636
rect 10413 41627 10471 41633
rect 12066 41624 12072 41636
rect 12124 41624 12130 41676
rect 14292 41664 14320 41695
rect 18506 41692 18512 41704
rect 18564 41692 18570 41744
rect 18616 41732 18644 41772
rect 19429 41769 19441 41803
rect 19475 41800 19487 41803
rect 20622 41800 20628 41812
rect 19475 41772 20628 41800
rect 19475 41769 19487 41772
rect 19429 41763 19487 41769
rect 20622 41760 20628 41772
rect 20680 41760 20686 41812
rect 21818 41800 21824 41812
rect 21779 41772 21824 41800
rect 21818 41760 21824 41772
rect 21876 41760 21882 41812
rect 22002 41760 22008 41812
rect 22060 41800 22066 41812
rect 26789 41803 26847 41809
rect 22060 41772 25636 41800
rect 22060 41760 22066 41772
rect 22094 41732 22100 41744
rect 18616 41704 22100 41732
rect 22094 41692 22100 41704
rect 22152 41692 22158 41744
rect 22186 41692 22192 41744
rect 22244 41732 22250 41744
rect 24673 41735 24731 41741
rect 24673 41732 24685 41735
rect 22244 41704 24685 41732
rect 22244 41692 22250 41704
rect 24673 41701 24685 41704
rect 24719 41732 24731 41735
rect 24719 41704 25544 41732
rect 24719 41701 24731 41704
rect 24673 41695 24731 41701
rect 14737 41667 14795 41673
rect 14737 41664 14749 41667
rect 14292 41636 14749 41664
rect 14737 41633 14749 41636
rect 14783 41633 14795 41667
rect 14737 41627 14795 41633
rect 17770 41624 17776 41676
rect 17828 41664 17834 41676
rect 17828 41636 18368 41664
rect 17828 41624 17834 41636
rect 1578 41596 1584 41608
rect 1539 41568 1584 41596
rect 1578 41556 1584 41568
rect 1636 41556 1642 41608
rect 8386 41556 8392 41608
rect 8444 41596 8450 41608
rect 8941 41599 8999 41605
rect 8941 41596 8953 41599
rect 8444 41568 8953 41596
rect 8444 41556 8450 41568
rect 8941 41565 8953 41568
rect 8987 41565 8999 41599
rect 8941 41559 8999 41565
rect 10042 41556 10048 41608
rect 10100 41596 10106 41608
rect 10689 41599 10747 41605
rect 10689 41596 10701 41599
rect 10100 41568 10701 41596
rect 10100 41556 10106 41568
rect 10689 41565 10701 41568
rect 10735 41565 10747 41599
rect 14090 41596 14096 41608
rect 14051 41568 14096 41596
rect 10689 41559 10747 41565
rect 14090 41556 14096 41568
rect 14148 41556 14154 41608
rect 15004 41599 15062 41605
rect 15004 41565 15016 41599
rect 15050 41596 15062 41599
rect 15378 41596 15384 41608
rect 15050 41568 15384 41596
rect 15050 41565 15062 41568
rect 15004 41559 15062 41565
rect 15378 41556 15384 41568
rect 15436 41556 15442 41608
rect 16853 41599 16911 41605
rect 16853 41565 16865 41599
rect 16899 41596 16911 41599
rect 17954 41596 17960 41608
rect 16899 41568 17960 41596
rect 16899 41565 16911 41568
rect 16853 41559 16911 41565
rect 17954 41556 17960 41568
rect 18012 41556 18018 41608
rect 18340 41605 18368 41636
rect 19334 41624 19340 41676
rect 19392 41664 19398 41676
rect 19981 41667 20039 41673
rect 19981 41664 19993 41667
rect 19392 41636 19993 41664
rect 19392 41624 19398 41636
rect 19981 41633 19993 41636
rect 20027 41664 20039 41667
rect 20162 41664 20168 41676
rect 20027 41636 20168 41664
rect 20027 41633 20039 41636
rect 19981 41627 20039 41633
rect 20162 41624 20168 41636
rect 20220 41624 20226 41676
rect 22281 41667 22339 41673
rect 22281 41633 22293 41667
rect 22327 41664 22339 41667
rect 23661 41667 23719 41673
rect 23661 41664 23673 41667
rect 22327 41636 23673 41664
rect 22327 41633 22339 41636
rect 22281 41627 22339 41633
rect 23661 41633 23673 41636
rect 23707 41633 23719 41667
rect 23661 41627 23719 41633
rect 25314 41624 25320 41676
rect 25372 41664 25378 41676
rect 25516 41673 25544 41704
rect 25608 41673 25636 41772
rect 26789 41769 26801 41803
rect 26835 41800 26847 41803
rect 27982 41800 27988 41812
rect 26835 41772 27988 41800
rect 26835 41769 26847 41772
rect 26789 41763 26847 41769
rect 27982 41760 27988 41772
rect 28040 41760 28046 41812
rect 28810 41760 28816 41812
rect 28868 41760 28874 41812
rect 29822 41760 29828 41812
rect 29880 41800 29886 41812
rect 29880 41772 30144 41800
rect 29880 41760 29886 41772
rect 25958 41692 25964 41744
rect 26016 41732 26022 41744
rect 26418 41732 26424 41744
rect 26016 41704 26424 41732
rect 26016 41692 26022 41704
rect 26418 41692 26424 41704
rect 26476 41692 26482 41744
rect 26973 41735 27031 41741
rect 26973 41701 26985 41735
rect 27019 41701 27031 41735
rect 26973 41695 27031 41701
rect 27433 41735 27491 41741
rect 27433 41701 27445 41735
rect 27479 41732 27491 41735
rect 28828 41732 28856 41760
rect 30116 41732 30144 41772
rect 30558 41760 30564 41812
rect 30616 41800 30622 41812
rect 30852 41800 30880 42044
rect 30616 41772 30880 41800
rect 30616 41760 30622 41772
rect 27479 41704 28488 41732
rect 28828 41704 29132 41732
rect 30116 41704 30604 41732
rect 27479 41701 27491 41704
rect 27433 41695 27491 41701
rect 25409 41667 25467 41673
rect 25409 41664 25421 41667
rect 25372 41636 25421 41664
rect 25372 41624 25378 41636
rect 25409 41633 25421 41636
rect 25455 41633 25467 41667
rect 25409 41627 25467 41633
rect 25501 41667 25559 41673
rect 25501 41633 25513 41667
rect 25547 41633 25559 41667
rect 25501 41627 25559 41633
rect 25593 41667 25651 41673
rect 25593 41633 25605 41667
rect 25639 41633 25651 41667
rect 25593 41627 25651 41633
rect 25682 41624 25688 41676
rect 25740 41664 25746 41676
rect 26988 41664 27016 41695
rect 25740 41636 25785 41664
rect 25884 41636 27016 41664
rect 25740 41624 25746 41636
rect 18325 41599 18383 41605
rect 18325 41565 18337 41599
rect 18371 41565 18383 41599
rect 18325 41559 18383 41565
rect 19886 41556 19892 41608
rect 19944 41596 19950 41608
rect 20625 41599 20683 41605
rect 20625 41596 20637 41599
rect 19944 41568 20637 41596
rect 19944 41556 19950 41568
rect 20625 41565 20637 41568
rect 20671 41565 20683 41599
rect 20625 41559 20683 41565
rect 20714 41556 20720 41608
rect 20772 41596 20778 41608
rect 22925 41599 22983 41605
rect 22925 41596 22937 41599
rect 20772 41568 22937 41596
rect 20772 41556 20778 41568
rect 9125 41531 9183 41537
rect 9125 41497 9137 41531
rect 9171 41497 9183 41531
rect 9125 41491 9183 41497
rect 11701 41531 11759 41537
rect 11701 41497 11713 41531
rect 11747 41528 11759 41531
rect 12342 41528 12348 41540
rect 11747 41500 12348 41528
rect 11747 41497 11759 41500
rect 11701 41491 11759 41497
rect 1397 41463 1455 41469
rect 1397 41429 1409 41463
rect 1443 41460 1455 41463
rect 9140 41460 9168 41491
rect 12342 41488 12348 41500
rect 12400 41488 12406 41540
rect 17589 41531 17647 41537
rect 17589 41497 17601 41531
rect 17635 41528 17647 41531
rect 18230 41528 18236 41540
rect 17635 41500 18236 41528
rect 17635 41497 17647 41500
rect 17589 41491 17647 41497
rect 18230 41488 18236 41500
rect 18288 41488 18294 41540
rect 19702 41528 19708 41540
rect 19663 41500 19708 41528
rect 19702 41488 19708 41500
rect 19760 41488 19766 41540
rect 20070 41488 20076 41540
rect 20128 41528 20134 41540
rect 20824 41528 20852 41568
rect 22925 41565 22937 41568
rect 22971 41565 22983 41599
rect 23566 41596 23572 41608
rect 23527 41568 23572 41596
rect 22925 41559 22983 41565
rect 23566 41556 23572 41568
rect 23624 41556 23630 41608
rect 24489 41599 24547 41605
rect 24489 41565 24501 41599
rect 24535 41596 24547 41599
rect 24762 41596 24768 41608
rect 24535 41568 24768 41596
rect 24535 41565 24547 41568
rect 24489 41559 24547 41565
rect 24762 41556 24768 41568
rect 24820 41556 24826 41608
rect 25884 41596 25912 41636
rect 24872 41568 25912 41596
rect 20128 41500 20852 41528
rect 22373 41531 22431 41537
rect 20128 41488 20134 41500
rect 22373 41497 22385 41531
rect 22419 41528 22431 41531
rect 24026 41528 24032 41540
rect 22419 41500 24032 41528
rect 22419 41497 22431 41500
rect 22373 41491 22431 41497
rect 24026 41488 24032 41500
rect 24084 41488 24090 41540
rect 24302 41488 24308 41540
rect 24360 41528 24366 41540
rect 24872 41528 24900 41568
rect 27522 41556 27528 41608
rect 27580 41596 27586 41608
rect 27617 41599 27675 41605
rect 27617 41596 27629 41599
rect 27580 41568 27629 41596
rect 27580 41556 27586 41568
rect 27617 41565 27629 41568
rect 27663 41565 27675 41599
rect 27617 41559 27675 41565
rect 27893 41599 27951 41605
rect 27893 41565 27905 41599
rect 27939 41596 27951 41599
rect 28166 41596 28172 41608
rect 27939 41568 28172 41596
rect 27939 41565 27951 41568
rect 27893 41559 27951 41565
rect 28166 41556 28172 41568
rect 28224 41556 28230 41608
rect 24360 41500 24900 41528
rect 24360 41488 24366 41500
rect 25130 41488 25136 41540
rect 25188 41528 25194 41540
rect 25188 41500 25452 41528
rect 25188 41488 25194 41500
rect 1443 41432 9168 41460
rect 16945 41463 17003 41469
rect 1443 41429 1455 41432
rect 1397 41423 1455 41429
rect 16945 41429 16957 41463
rect 16991 41460 17003 41463
rect 18138 41460 18144 41472
rect 16991 41432 18144 41460
rect 16991 41429 17003 41432
rect 16945 41423 17003 41429
rect 18138 41420 18144 41432
rect 18196 41420 18202 41472
rect 19518 41420 19524 41472
rect 19576 41460 19582 41472
rect 19889 41463 19947 41469
rect 19889 41460 19901 41463
rect 19576 41432 19901 41460
rect 19576 41420 19582 41432
rect 19889 41429 19901 41432
rect 19935 41429 19947 41463
rect 19889 41423 19947 41429
rect 20714 41420 20720 41472
rect 20772 41460 20778 41472
rect 20809 41463 20867 41469
rect 20809 41460 20821 41463
rect 20772 41432 20821 41460
rect 20772 41420 20778 41432
rect 20809 41429 20821 41432
rect 20855 41429 20867 41463
rect 20809 41423 20867 41429
rect 22281 41463 22339 41469
rect 22281 41429 22293 41463
rect 22327 41460 22339 41463
rect 23017 41463 23075 41469
rect 23017 41460 23029 41463
rect 22327 41432 23029 41460
rect 22327 41429 22339 41432
rect 22281 41423 22339 41429
rect 23017 41429 23029 41432
rect 23063 41429 23075 41463
rect 23017 41423 23075 41429
rect 24854 41420 24860 41472
rect 24912 41460 24918 41472
rect 25225 41463 25283 41469
rect 25225 41460 25237 41463
rect 24912 41432 25237 41460
rect 24912 41420 24918 41432
rect 25225 41429 25237 41432
rect 25271 41429 25283 41463
rect 25424 41460 25452 41500
rect 25498 41488 25504 41540
rect 25556 41528 25562 41540
rect 26050 41528 26056 41540
rect 25556 41500 26056 41528
rect 25556 41488 25562 41500
rect 26050 41488 26056 41500
rect 26108 41488 26114 41540
rect 26789 41531 26847 41537
rect 26789 41497 26801 41531
rect 26835 41528 26847 41531
rect 27706 41528 27712 41540
rect 26835 41500 27712 41528
rect 26835 41497 26847 41500
rect 26789 41491 26847 41497
rect 27706 41488 27712 41500
rect 27764 41488 27770 41540
rect 27801 41531 27859 41537
rect 27801 41497 27813 41531
rect 27847 41528 27859 41531
rect 27847 41500 27936 41528
rect 27847 41497 27859 41500
rect 27801 41491 27859 41497
rect 25774 41460 25780 41472
rect 25424 41432 25780 41460
rect 25225 41423 25283 41429
rect 25774 41420 25780 41432
rect 25832 41420 25838 41472
rect 26510 41420 26516 41472
rect 26568 41460 26574 41472
rect 27908 41460 27936 41500
rect 26568 41432 27936 41460
rect 26568 41420 26574 41432
rect 27982 41420 27988 41472
rect 28040 41460 28046 41472
rect 28353 41463 28411 41469
rect 28353 41460 28365 41463
rect 28040 41432 28365 41460
rect 28040 41420 28046 41432
rect 28353 41429 28365 41432
rect 28399 41429 28411 41463
rect 28460 41460 28488 41704
rect 28534 41556 28540 41608
rect 28592 41596 28598 41608
rect 28629 41599 28687 41605
rect 28629 41596 28641 41599
rect 28592 41568 28641 41596
rect 28592 41556 28598 41568
rect 28629 41565 28641 41568
rect 28675 41565 28687 41599
rect 28721 41593 28779 41599
rect 28721 41586 28733 41593
rect 28767 41586 28779 41593
rect 28629 41559 28687 41565
rect 28718 41534 28724 41586
rect 28776 41534 28782 41586
rect 28810 41556 28816 41608
rect 28868 41593 28874 41608
rect 29009 41599 29067 41605
rect 28868 41565 28910 41593
rect 29009 41565 29021 41599
rect 29055 41596 29067 41599
rect 29104 41596 29132 41704
rect 29178 41624 29184 41676
rect 29236 41664 29242 41676
rect 29236 41636 29776 41664
rect 29236 41624 29242 41636
rect 29748 41605 29776 41636
rect 29055 41568 29132 41596
rect 29733 41599 29791 41605
rect 29055 41565 29067 41568
rect 28868 41556 28874 41565
rect 29009 41559 29067 41565
rect 29733 41565 29745 41599
rect 29779 41565 29791 41599
rect 29914 41596 29920 41608
rect 29875 41568 29920 41596
rect 29733 41559 29791 41565
rect 29914 41556 29920 41568
rect 29972 41556 29978 41608
rect 30009 41599 30067 41605
rect 30009 41565 30021 41599
rect 30055 41596 30067 41599
rect 30098 41596 30104 41608
rect 30055 41568 30104 41596
rect 30055 41565 30067 41568
rect 30009 41559 30067 41565
rect 30098 41556 30104 41568
rect 30156 41556 30162 41608
rect 30576 41528 30604 41704
rect 31110 41528 31116 41540
rect 29012 41500 30144 41528
rect 29012 41460 29040 41500
rect 30116 41472 30144 41500
rect 30392 41500 30604 41528
rect 30852 41500 31116 41528
rect 28460 41432 29040 41460
rect 28353 41423 28411 41429
rect 29086 41420 29092 41472
rect 29144 41460 29150 41472
rect 29549 41463 29607 41469
rect 29549 41460 29561 41463
rect 29144 41432 29561 41460
rect 29144 41420 29150 41432
rect 29549 41429 29561 41432
rect 29595 41429 29607 41463
rect 29549 41423 29607 41429
rect 30098 41420 30104 41472
rect 30156 41420 30162 41472
rect 30282 41420 30288 41472
rect 30340 41460 30346 41472
rect 30392 41460 30420 41500
rect 30852 41472 30880 41500
rect 31110 41488 31116 41500
rect 31168 41488 31174 41540
rect 31312 41528 31340 42248
rect 31404 42248 31524 42276
rect 31404 41812 31432 42248
rect 31386 41760 31392 41812
rect 31444 41760 31450 41812
rect 31220 41500 31340 41528
rect 30340 41432 30420 41460
rect 30340 41420 30346 41432
rect 30466 41420 30472 41472
rect 30524 41460 30530 41472
rect 30650 41460 30656 41472
rect 30524 41432 30656 41460
rect 30524 41420 30530 41432
rect 30650 41420 30656 41432
rect 30708 41420 30714 41472
rect 30834 41420 30840 41472
rect 30892 41420 30898 41472
rect 1104 41370 30820 41392
rect 1104 41318 10880 41370
rect 10932 41318 10944 41370
rect 10996 41318 11008 41370
rect 11060 41318 11072 41370
rect 11124 41318 11136 41370
rect 11188 41318 20811 41370
rect 20863 41318 20875 41370
rect 20927 41318 20939 41370
rect 20991 41318 21003 41370
rect 21055 41318 21067 41370
rect 21119 41318 30820 41370
rect 31110 41352 31116 41404
rect 31168 41392 31174 41404
rect 31220 41392 31248 41500
rect 31168 41364 31248 41392
rect 31168 41352 31174 41364
rect 1104 41296 30820 41318
rect 15286 41216 15292 41268
rect 15344 41256 15350 41268
rect 15381 41259 15439 41265
rect 15381 41256 15393 41259
rect 15344 41228 15393 41256
rect 15344 41216 15350 41228
rect 15381 41225 15393 41228
rect 15427 41225 15439 41259
rect 15381 41219 15439 41225
rect 17586 41216 17592 41268
rect 17644 41216 17650 41268
rect 18598 41256 18604 41268
rect 18559 41228 18604 41256
rect 18598 41216 18604 41228
rect 18656 41216 18662 41268
rect 19245 41259 19303 41265
rect 19245 41225 19257 41259
rect 19291 41256 19303 41259
rect 19978 41256 19984 41268
rect 19291 41228 19984 41256
rect 19291 41225 19303 41228
rect 19245 41219 19303 41225
rect 19978 41216 19984 41228
rect 20036 41256 20042 41268
rect 20349 41259 20407 41265
rect 20349 41256 20361 41259
rect 20036 41228 20361 41256
rect 20036 41216 20042 41228
rect 20349 41225 20361 41228
rect 20395 41225 20407 41259
rect 21177 41259 21235 41265
rect 21177 41256 21189 41259
rect 20349 41219 20407 41225
rect 20456 41228 21189 41256
rect 1854 41148 1860 41200
rect 1912 41188 1918 41200
rect 15933 41191 15991 41197
rect 1912 41160 15332 41188
rect 1912 41148 1918 41160
rect 1578 41120 1584 41132
rect 1539 41092 1584 41120
rect 1578 41080 1584 41092
rect 1636 41080 1642 41132
rect 15197 41123 15255 41129
rect 15197 41089 15209 41123
rect 15243 41089 15255 41123
rect 15304 41120 15332 41160
rect 15933 41157 15945 41191
rect 15979 41188 15991 41191
rect 16390 41188 16396 41200
rect 15979 41160 16396 41188
rect 15979 41157 15991 41160
rect 15933 41151 15991 41157
rect 16390 41148 16396 41160
rect 16448 41148 16454 41200
rect 17604 41188 17632 41216
rect 18322 41188 18328 41200
rect 17604 41160 17721 41188
rect 17693 41132 17721 41160
rect 17880 41160 18328 41188
rect 16666 41120 16672 41132
rect 15304 41092 16252 41120
rect 16627 41092 16672 41120
rect 15197 41083 15255 41089
rect 15212 41052 15240 41083
rect 15746 41052 15752 41064
rect 15212 41024 15752 41052
rect 15746 41012 15752 41024
rect 15804 41052 15810 41064
rect 16117 41055 16175 41061
rect 16117 41052 16129 41055
rect 15804 41024 16129 41052
rect 15804 41012 15810 41024
rect 16117 41021 16129 41024
rect 16163 41021 16175 41055
rect 16224 41052 16252 41092
rect 16666 41080 16672 41092
rect 16724 41080 16730 41132
rect 17494 41080 17500 41132
rect 17552 41120 17558 41132
rect 17589 41123 17647 41129
rect 17589 41120 17601 41123
rect 17552 41092 17601 41120
rect 17552 41080 17558 41092
rect 17589 41089 17601 41092
rect 17635 41089 17647 41123
rect 17589 41083 17647 41089
rect 17678 41126 17736 41132
rect 17678 41092 17690 41126
rect 17724 41092 17736 41126
rect 17678 41086 17736 41092
rect 17794 41123 17852 41129
rect 17794 41089 17806 41123
rect 17840 41120 17852 41123
rect 17880 41120 17908 41160
rect 18322 41148 18328 41160
rect 18380 41148 18386 41200
rect 19153 41191 19211 41197
rect 19153 41157 19165 41191
rect 19199 41188 19211 41191
rect 19610 41188 19616 41200
rect 19199 41160 19616 41188
rect 19199 41157 19211 41160
rect 19153 41151 19211 41157
rect 19610 41148 19616 41160
rect 19668 41148 19674 41200
rect 19702 41148 19708 41200
rect 19760 41188 19766 41200
rect 20165 41191 20223 41197
rect 20165 41188 20177 41191
rect 19760 41160 20177 41188
rect 19760 41148 19766 41160
rect 20165 41157 20177 41160
rect 20211 41188 20223 41191
rect 20456 41188 20484 41228
rect 21177 41225 21189 41228
rect 21223 41225 21235 41259
rect 21177 41219 21235 41225
rect 21910 41216 21916 41268
rect 21968 41216 21974 41268
rect 22002 41216 22008 41268
rect 22060 41256 22066 41268
rect 22462 41256 22468 41268
rect 22060 41228 22468 41256
rect 22060 41216 22066 41228
rect 22462 41216 22468 41228
rect 22520 41216 22526 41268
rect 23106 41256 23112 41268
rect 22572 41228 23112 41256
rect 20211 41160 20484 41188
rect 21085 41191 21143 41197
rect 20211 41157 20223 41160
rect 20165 41151 20223 41157
rect 21085 41157 21097 41191
rect 21131 41188 21143 41191
rect 21928 41188 21956 41216
rect 21131 41160 21956 41188
rect 21131 41157 21143 41160
rect 21085 41151 21143 41157
rect 22278 41148 22284 41200
rect 22336 41188 22342 41200
rect 22572 41188 22600 41228
rect 23106 41216 23112 41228
rect 23164 41216 23170 41268
rect 25406 41216 25412 41268
rect 25464 41216 25470 41268
rect 25774 41256 25780 41268
rect 25735 41228 25780 41256
rect 25774 41216 25780 41228
rect 25832 41216 25838 41268
rect 26234 41216 26240 41268
rect 26292 41256 26298 41268
rect 27706 41256 27712 41268
rect 26292 41228 27712 41256
rect 26292 41216 26298 41228
rect 27706 41216 27712 41228
rect 27764 41216 27770 41268
rect 27890 41216 27896 41268
rect 27948 41256 27954 41268
rect 28074 41256 28080 41268
rect 27948 41228 28080 41256
rect 27948 41216 27954 41228
rect 28074 41216 28080 41228
rect 28132 41216 28138 41268
rect 28718 41256 28724 41268
rect 28625 41228 28724 41256
rect 25225 41191 25283 41197
rect 22336 41160 22600 41188
rect 24596 41160 25184 41188
rect 22336 41148 22342 41160
rect 17840 41092 17908 41120
rect 17957 41123 18015 41129
rect 17840 41089 17852 41092
rect 17794 41083 17852 41089
rect 17957 41089 17969 41123
rect 18003 41089 18015 41123
rect 17957 41083 18015 41089
rect 18417 41123 18475 41129
rect 18417 41089 18429 41123
rect 18463 41120 18475 41123
rect 19334 41120 19340 41132
rect 18463 41092 19340 41120
rect 18463 41089 18475 41092
rect 18417 41083 18475 41089
rect 17972 41052 18000 41083
rect 19334 41080 19340 41092
rect 19392 41080 19398 41132
rect 21358 41080 21364 41132
rect 21416 41120 21422 41132
rect 21634 41120 21640 41132
rect 21416 41092 21640 41120
rect 21416 41080 21422 41092
rect 21634 41080 21640 41092
rect 21692 41080 21698 41132
rect 22462 41120 22468 41132
rect 22423 41092 22468 41120
rect 22462 41080 22468 41092
rect 22520 41080 22526 41132
rect 22738 41080 22744 41132
rect 22796 41120 22802 41132
rect 23109 41123 23167 41129
rect 23109 41120 23121 41123
rect 22796 41092 23121 41120
rect 22796 41080 22802 41092
rect 23109 41089 23121 41092
rect 23155 41089 23167 41123
rect 23109 41083 23167 41089
rect 23198 41080 23204 41132
rect 23256 41120 23262 41132
rect 23293 41123 23351 41129
rect 23293 41120 23305 41123
rect 23256 41092 23305 41120
rect 23256 41080 23262 41092
rect 23293 41089 23305 41092
rect 23339 41120 23351 41123
rect 23382 41120 23388 41132
rect 23339 41092 23388 41120
rect 23339 41089 23351 41092
rect 23293 41083 23351 41089
rect 23382 41080 23388 41092
rect 23440 41080 23446 41132
rect 16224 41024 18000 41052
rect 16117 41015 16175 41021
rect 20162 41012 20168 41064
rect 20220 41052 20226 41064
rect 20438 41052 20444 41064
rect 20220 41024 20444 41052
rect 20220 41012 20226 41024
rect 20438 41012 20444 41024
rect 20496 41012 20502 41064
rect 17494 40944 17500 40996
rect 17552 40984 17558 40996
rect 18690 40984 18696 40996
rect 17552 40956 18696 40984
rect 17552 40944 17558 40956
rect 18690 40944 18696 40956
rect 18748 40984 18754 40996
rect 19886 40984 19892 40996
rect 18748 40956 19334 40984
rect 19847 40956 19892 40984
rect 18748 40944 18754 40956
rect 1397 40919 1455 40925
rect 1397 40885 1409 40919
rect 1443 40916 1455 40919
rect 8202 40916 8208 40928
rect 1443 40888 8208 40916
rect 1443 40885 1455 40888
rect 1397 40879 1455 40885
rect 8202 40876 8208 40888
rect 8260 40876 8266 40928
rect 16853 40919 16911 40925
rect 16853 40885 16865 40919
rect 16899 40916 16911 40919
rect 17034 40916 17040 40928
rect 16899 40888 17040 40916
rect 16899 40885 16911 40888
rect 16853 40879 16911 40885
rect 17034 40876 17040 40888
rect 17092 40876 17098 40928
rect 17313 40919 17371 40925
rect 17313 40885 17325 40919
rect 17359 40916 17371 40919
rect 17586 40916 17592 40928
rect 17359 40888 17592 40916
rect 17359 40885 17371 40888
rect 17313 40879 17371 40885
rect 17586 40876 17592 40888
rect 17644 40876 17650 40928
rect 19306 40916 19334 40956
rect 19886 40944 19892 40956
rect 19944 40944 19950 40996
rect 21174 40944 21180 40996
rect 21232 40984 21238 40996
rect 21726 40984 21732 40996
rect 21232 40956 21732 40984
rect 21232 40944 21238 40956
rect 21726 40944 21732 40956
rect 21784 40984 21790 40996
rect 22002 40984 22008 40996
rect 21784 40956 22008 40984
rect 21784 40944 21790 40956
rect 22002 40944 22008 40956
rect 22060 40944 22066 40996
rect 23566 40984 23572 40996
rect 22572 40956 23572 40984
rect 21266 40916 21272 40928
rect 19306 40888 21272 40916
rect 21266 40876 21272 40888
rect 21324 40876 21330 40928
rect 21542 40876 21548 40928
rect 21600 40916 21606 40928
rect 22572 40925 22600 40956
rect 23566 40944 23572 40956
rect 23624 40944 23630 40996
rect 24596 40984 24624 41160
rect 25156 41129 25184 41160
rect 25225 41157 25237 41191
rect 25271 41188 25283 41191
rect 25424 41188 25452 41216
rect 28166 41188 28172 41200
rect 25271 41160 25452 41188
rect 27816 41160 28172 41188
rect 25271 41157 25283 41160
rect 25225 41151 25283 41157
rect 25125 41123 25184 41129
rect 25125 41089 25137 41123
rect 25171 41092 25184 41123
rect 25961 41123 26019 41129
rect 25961 41120 25973 41123
rect 25332 41092 25973 41120
rect 25171 41089 25183 41092
rect 25125 41083 25183 41089
rect 24762 41012 24768 41064
rect 24820 41052 24826 41064
rect 25332 41052 25360 41092
rect 25961 41089 25973 41092
rect 26007 41089 26019 41123
rect 25961 41083 26019 41089
rect 27525 41123 27583 41129
rect 27525 41089 27537 41123
rect 27571 41120 27583 41123
rect 27614 41120 27620 41132
rect 27571 41092 27620 41120
rect 27571 41089 27583 41092
rect 27525 41083 27583 41089
rect 27614 41080 27620 41092
rect 27672 41080 27678 41132
rect 27816 41129 27844 41160
rect 28166 41148 28172 41160
rect 28224 41148 28230 41200
rect 28258 41148 28264 41200
rect 28316 41148 28322 41200
rect 27801 41123 27859 41129
rect 27801 41089 27813 41123
rect 27847 41089 27859 41123
rect 28276 41120 28304 41148
rect 28625 41135 28653 41228
rect 28718 41216 28724 41228
rect 28776 41216 28782 41268
rect 28902 41216 28908 41268
rect 28960 41256 28966 41268
rect 31846 41256 31852 41268
rect 28960 41228 29684 41256
rect 28960 41216 28966 41228
rect 29656 41188 29684 41228
rect 29840 41228 31852 41256
rect 28736 41160 29052 41188
rect 29656 41160 29730 41188
rect 28610 41129 28668 41135
rect 28736 41129 28764 41160
rect 28491 41123 28549 41129
rect 28491 41120 28503 41123
rect 28276 41092 28503 41120
rect 27801 41083 27859 41089
rect 28491 41089 28503 41092
rect 28537 41089 28549 41123
rect 28610 41095 28622 41129
rect 28656 41095 28668 41129
rect 28610 41089 28668 41095
rect 28710 41123 28768 41129
rect 28710 41089 28722 41123
rect 28756 41089 28768 41123
rect 28917 41123 28975 41129
rect 28917 41110 28929 41123
rect 28491 41083 28549 41089
rect 28710 41083 28768 41089
rect 28828 41089 28929 41110
rect 28963 41089 28975 41123
rect 28828 41083 28975 41089
rect 28828 41082 28948 41083
rect 24820 41024 25360 41052
rect 26237 41055 26295 41061
rect 24820 41012 24826 41024
rect 26237 41021 26249 41055
rect 26283 41052 26295 41055
rect 26418 41052 26424 41064
rect 26283 41024 26424 41052
rect 26283 41021 26295 41024
rect 26237 41015 26295 41021
rect 26418 41012 26424 41024
rect 26476 41012 26482 41064
rect 27341 41055 27399 41061
rect 27341 41021 27353 41055
rect 27387 41052 27399 41055
rect 28828 41052 28856 41082
rect 27387 41024 28856 41052
rect 27387 41021 27399 41024
rect 27341 41015 27399 41021
rect 24670 40984 24676 40996
rect 24596 40956 24676 40984
rect 24670 40944 24676 40956
rect 24728 40944 24734 40996
rect 25130 40944 25136 40996
rect 25188 40984 25194 40996
rect 26145 40987 26203 40993
rect 26145 40984 26157 40987
rect 25188 40956 26157 40984
rect 25188 40944 25194 40956
rect 26145 40953 26157 40956
rect 26191 40984 26203 40987
rect 27430 40984 27436 40996
rect 26191 40956 27436 40984
rect 26191 40953 26203 40956
rect 26145 40947 26203 40953
rect 27430 40944 27436 40956
rect 27488 40944 27494 40996
rect 22557 40919 22615 40925
rect 22557 40916 22569 40919
rect 21600 40888 22569 40916
rect 21600 40876 21606 40888
rect 22557 40885 22569 40888
rect 22603 40885 22615 40919
rect 22557 40879 22615 40885
rect 22922 40876 22928 40928
rect 22980 40916 22986 40928
rect 23109 40919 23167 40925
rect 23109 40916 23121 40919
rect 22980 40888 23121 40916
rect 22980 40876 22986 40888
rect 23109 40885 23121 40888
rect 23155 40885 23167 40919
rect 23109 40879 23167 40885
rect 23290 40876 23296 40928
rect 23348 40916 23354 40928
rect 27522 40916 27528 40928
rect 23348 40888 27528 40916
rect 23348 40876 23354 40888
rect 27522 40876 27528 40888
rect 27580 40876 27586 40928
rect 28166 40876 28172 40928
rect 28224 40916 28230 40928
rect 28261 40919 28319 40925
rect 28261 40916 28273 40919
rect 28224 40888 28273 40916
rect 28224 40876 28230 40888
rect 28261 40885 28273 40888
rect 28307 40885 28319 40919
rect 28261 40879 28319 40885
rect 28810 40876 28816 40928
rect 28868 40916 28874 40928
rect 29024 40916 29052 41160
rect 29702 41129 29730 41160
rect 29840 41132 29868 41228
rect 31846 41216 31852 41228
rect 31904 41216 31910 41268
rect 29687 41123 29745 41129
rect 29687 41089 29699 41123
rect 29733 41089 29745 41123
rect 29687 41083 29745 41089
rect 29822 41126 29880 41132
rect 29822 41092 29834 41126
rect 29868 41092 29880 41126
rect 29822 41086 29880 41092
rect 29914 41080 29920 41132
rect 29972 41129 29978 41132
rect 29972 41120 29980 41129
rect 30098 41120 30104 41132
rect 29972 41092 30017 41120
rect 30059 41092 30104 41120
rect 29972 41083 29980 41092
rect 29972 41080 29978 41083
rect 30098 41080 30104 41092
rect 30156 41080 30162 41132
rect 28868 40888 29052 40916
rect 29457 40919 29515 40925
rect 28868 40876 28874 40888
rect 29457 40885 29469 40919
rect 29503 40916 29515 40919
rect 29822 40916 29828 40928
rect 29503 40888 29828 40916
rect 29503 40885 29515 40888
rect 29457 40879 29515 40885
rect 29822 40876 29828 40888
rect 29880 40876 29886 40928
rect 1104 40826 30820 40848
rect 1104 40774 5915 40826
rect 5967 40774 5979 40826
rect 6031 40774 6043 40826
rect 6095 40774 6107 40826
rect 6159 40774 6171 40826
rect 6223 40774 15846 40826
rect 15898 40774 15910 40826
rect 15962 40774 15974 40826
rect 16026 40774 16038 40826
rect 16090 40774 16102 40826
rect 16154 40774 25776 40826
rect 25828 40774 25840 40826
rect 25892 40774 25904 40826
rect 25956 40774 25968 40826
rect 26020 40774 26032 40826
rect 26084 40774 30820 40826
rect 1104 40752 30820 40774
rect 8662 40672 8668 40724
rect 8720 40712 8726 40724
rect 10134 40712 10140 40724
rect 8720 40684 10140 40712
rect 8720 40672 8726 40684
rect 10134 40672 10140 40684
rect 10192 40672 10198 40724
rect 17221 40715 17279 40721
rect 17221 40681 17233 40715
rect 17267 40712 17279 40715
rect 17402 40712 17408 40724
rect 17267 40684 17408 40712
rect 17267 40681 17279 40684
rect 17221 40675 17279 40681
rect 17402 40672 17408 40684
rect 17460 40672 17466 40724
rect 17862 40712 17868 40724
rect 17823 40684 17868 40712
rect 17862 40672 17868 40684
rect 17920 40672 17926 40724
rect 19334 40712 19340 40724
rect 19295 40684 19340 40712
rect 19334 40672 19340 40684
rect 19392 40672 19398 40724
rect 23474 40672 23480 40724
rect 23532 40712 23538 40724
rect 23532 40684 28580 40712
rect 23532 40672 23538 40684
rect 9858 40604 9864 40656
rect 9916 40644 9922 40656
rect 9916 40616 9987 40644
rect 9916 40604 9922 40616
rect 8386 40576 8392 40588
rect 8036 40548 8392 40576
rect 8036 40517 8064 40548
rect 8386 40536 8392 40548
rect 8444 40536 8450 40588
rect 8021 40511 8079 40517
rect 8021 40477 8033 40511
rect 8067 40477 8079 40511
rect 8202 40508 8208 40520
rect 8163 40480 8208 40508
rect 8021 40471 8079 40477
rect 8202 40468 8208 40480
rect 8260 40468 8266 40520
rect 9959 40517 9987 40616
rect 16942 40604 16948 40656
rect 17000 40644 17006 40656
rect 17310 40644 17316 40656
rect 17000 40616 17316 40644
rect 17000 40604 17006 40616
rect 17310 40604 17316 40616
rect 17368 40604 17374 40656
rect 21361 40647 21419 40653
rect 21361 40644 21373 40647
rect 19996 40616 21373 40644
rect 10134 40536 10140 40588
rect 10192 40576 10198 40588
rect 10192 40548 10272 40576
rect 10192 40536 10198 40548
rect 9841 40511 9899 40517
rect 9841 40477 9853 40511
rect 9887 40477 9899 40511
rect 9841 40471 9899 40477
rect 9934 40511 9992 40517
rect 9934 40477 9946 40511
rect 9980 40477 9992 40511
rect 9934 40471 9992 40477
rect 8389 40443 8447 40449
rect 8389 40409 8401 40443
rect 8435 40440 8447 40443
rect 9856 40440 9884 40471
rect 10042 40468 10048 40520
rect 10100 40508 10106 40520
rect 10244 40517 10272 40548
rect 10318 40536 10324 40588
rect 10376 40576 10382 40588
rect 11238 40576 11244 40588
rect 10376 40548 11244 40576
rect 10376 40536 10382 40548
rect 11238 40536 11244 40548
rect 11296 40576 11302 40588
rect 19886 40576 19892 40588
rect 11296 40548 19892 40576
rect 11296 40536 11302 40548
rect 19886 40536 19892 40548
rect 19944 40536 19950 40588
rect 10229 40511 10287 40517
rect 10100 40480 10145 40508
rect 10100 40468 10106 40480
rect 10229 40477 10241 40511
rect 10275 40477 10287 40511
rect 15746 40508 15752 40520
rect 15707 40480 15752 40508
rect 10229 40471 10287 40477
rect 15746 40468 15752 40480
rect 15804 40508 15810 40520
rect 16393 40511 16451 40517
rect 16393 40508 16405 40511
rect 15804 40480 16405 40508
rect 15804 40468 15810 40480
rect 16393 40477 16405 40480
rect 16439 40477 16451 40511
rect 16393 40471 16451 40477
rect 16942 40468 16948 40520
rect 17000 40508 17006 40520
rect 17037 40511 17095 40517
rect 17037 40508 17049 40511
rect 17000 40480 17049 40508
rect 17000 40468 17006 40480
rect 17037 40477 17049 40480
rect 17083 40477 17095 40511
rect 17037 40471 17095 40477
rect 17681 40511 17739 40517
rect 17681 40477 17693 40511
rect 17727 40508 17739 40511
rect 18046 40508 18052 40520
rect 17727 40480 18052 40508
rect 17727 40477 17739 40480
rect 17681 40471 17739 40477
rect 18046 40468 18052 40480
rect 18104 40468 18110 40520
rect 19245 40511 19303 40517
rect 19245 40508 19257 40511
rect 18432 40480 19257 40508
rect 11330 40440 11336 40452
rect 8435 40412 9812 40440
rect 9856 40412 11336 40440
rect 8435 40409 8447 40412
rect 8389 40403 8447 40409
rect 9585 40375 9643 40381
rect 9585 40341 9597 40375
rect 9631 40372 9643 40375
rect 9674 40372 9680 40384
rect 9631 40344 9680 40372
rect 9631 40341 9643 40344
rect 9585 40335 9643 40341
rect 9674 40332 9680 40344
rect 9732 40332 9738 40384
rect 9784 40372 9812 40412
rect 11330 40400 11336 40412
rect 11388 40400 11394 40452
rect 10134 40372 10140 40384
rect 9784 40344 10140 40372
rect 10134 40332 10140 40344
rect 10192 40332 10198 40384
rect 13998 40332 14004 40384
rect 14056 40372 14062 40384
rect 15933 40375 15991 40381
rect 15933 40372 15945 40375
rect 14056 40344 15945 40372
rect 14056 40332 14062 40344
rect 15933 40341 15945 40344
rect 15979 40341 15991 40375
rect 15933 40335 15991 40341
rect 16577 40375 16635 40381
rect 16577 40341 16589 40375
rect 16623 40372 16635 40375
rect 16850 40372 16856 40384
rect 16623 40344 16856 40372
rect 16623 40341 16635 40344
rect 16577 40335 16635 40341
rect 16850 40332 16856 40344
rect 16908 40332 16914 40384
rect 17954 40332 17960 40384
rect 18012 40372 18018 40384
rect 18432 40372 18460 40480
rect 19245 40477 19257 40480
rect 19291 40477 19303 40511
rect 19245 40471 19303 40477
rect 18509 40443 18567 40449
rect 18509 40409 18521 40443
rect 18555 40440 18567 40443
rect 19996 40440 20024 40616
rect 21361 40613 21373 40616
rect 21407 40644 21419 40647
rect 22462 40644 22468 40656
rect 21407 40616 22468 40644
rect 21407 40613 21419 40616
rect 21361 40607 21419 40613
rect 22462 40604 22468 40616
rect 22520 40604 22526 40656
rect 25317 40647 25375 40653
rect 25317 40613 25329 40647
rect 25363 40644 25375 40647
rect 27798 40644 27804 40656
rect 25363 40616 27804 40644
rect 25363 40613 25375 40616
rect 25317 40607 25375 40613
rect 27798 40604 27804 40616
rect 27856 40604 27862 40656
rect 22925 40579 22983 40585
rect 22925 40545 22937 40579
rect 22971 40576 22983 40579
rect 23474 40576 23480 40588
rect 22971 40548 23480 40576
rect 22971 40545 22983 40548
rect 22925 40539 22983 40545
rect 23474 40536 23480 40548
rect 23532 40536 23538 40588
rect 25774 40536 25780 40588
rect 25832 40576 25838 40588
rect 28261 40579 28319 40585
rect 25832 40548 27016 40576
rect 25832 40536 25838 40548
rect 20073 40511 20131 40517
rect 20073 40477 20085 40511
rect 20119 40508 20131 40511
rect 22094 40508 22100 40520
rect 20119 40480 22100 40508
rect 20119 40477 20131 40480
rect 20073 40471 20131 40477
rect 22094 40468 22100 40480
rect 22152 40468 22158 40520
rect 22278 40468 22284 40520
rect 22336 40508 22342 40520
rect 22462 40508 22468 40520
rect 22336 40480 22468 40508
rect 22336 40468 22342 40480
rect 22462 40468 22468 40480
rect 22520 40508 22526 40520
rect 23109 40511 23167 40517
rect 23109 40508 23121 40511
rect 22520 40480 23121 40508
rect 22520 40468 22526 40480
rect 23109 40477 23121 40480
rect 23155 40477 23167 40511
rect 23566 40508 23572 40520
rect 23527 40480 23572 40508
rect 23109 40471 23167 40477
rect 23566 40468 23572 40480
rect 23624 40468 23630 40520
rect 23845 40511 23903 40517
rect 23845 40477 23857 40511
rect 23891 40508 23903 40511
rect 24302 40508 24308 40520
rect 23891 40480 24308 40508
rect 23891 40477 23903 40480
rect 23845 40471 23903 40477
rect 24302 40468 24308 40480
rect 24360 40468 24366 40520
rect 25133 40511 25191 40517
rect 25133 40477 25145 40511
rect 25179 40508 25191 40511
rect 25179 40480 26924 40508
rect 25179 40477 25191 40480
rect 25133 40471 25191 40477
rect 25866 40440 25872 40452
rect 18555 40412 20024 40440
rect 20088 40412 23060 40440
rect 25827 40412 25872 40440
rect 18555 40409 18567 40412
rect 18509 40403 18567 40409
rect 18601 40375 18659 40381
rect 18601 40372 18613 40375
rect 18012 40344 18613 40372
rect 18012 40332 18018 40344
rect 18601 40341 18613 40344
rect 18647 40341 18659 40375
rect 18601 40335 18659 40341
rect 19610 40332 19616 40384
rect 19668 40372 19674 40384
rect 20088 40372 20116 40412
rect 19668 40344 20116 40372
rect 23032 40372 23060 40412
rect 25866 40400 25872 40412
rect 25924 40400 25930 40452
rect 26050 40440 26056 40452
rect 26011 40412 26056 40440
rect 26050 40400 26056 40412
rect 26108 40400 26114 40452
rect 26896 40449 26924 40480
rect 26237 40443 26295 40449
rect 26237 40440 26249 40443
rect 26160 40412 26249 40440
rect 26160 40372 26188 40412
rect 26237 40409 26249 40412
rect 26283 40409 26295 40443
rect 26237 40403 26295 40409
rect 26881 40443 26939 40449
rect 26881 40409 26893 40443
rect 26927 40409 26939 40443
rect 26988 40440 27016 40548
rect 27172 40548 28212 40576
rect 27172 40517 27200 40548
rect 27157 40511 27215 40517
rect 27157 40477 27169 40511
rect 27203 40477 27215 40511
rect 27157 40471 27215 40477
rect 27249 40511 27307 40517
rect 27249 40477 27261 40511
rect 27295 40477 27307 40511
rect 27249 40471 27307 40477
rect 27341 40511 27399 40517
rect 27341 40477 27353 40511
rect 27387 40477 27399 40511
rect 27341 40471 27399 40477
rect 27264 40440 27292 40471
rect 26988 40412 27292 40440
rect 26881 40403 26939 40409
rect 23032 40344 26188 40372
rect 19668 40332 19674 40344
rect 26326 40332 26332 40384
rect 26384 40372 26390 40384
rect 27356 40372 27384 40471
rect 27522 40468 27528 40520
rect 27580 40517 27586 40520
rect 27580 40511 27595 40517
rect 27583 40477 27595 40511
rect 27985 40511 28043 40517
rect 27985 40508 27997 40511
rect 27580 40471 27595 40477
rect 27724 40480 27997 40508
rect 27580 40468 27586 40471
rect 26384 40344 27384 40372
rect 26384 40332 26390 40344
rect 27430 40332 27436 40384
rect 27488 40372 27494 40384
rect 27724 40372 27752 40480
rect 27985 40477 27997 40480
rect 28031 40477 28043 40511
rect 27985 40471 28043 40477
rect 28184 40440 28212 40548
rect 28261 40545 28273 40579
rect 28307 40576 28319 40579
rect 28350 40576 28356 40588
rect 28307 40548 28356 40576
rect 28307 40545 28319 40548
rect 28261 40539 28319 40545
rect 28350 40536 28356 40548
rect 28408 40536 28414 40588
rect 28552 40576 28580 40684
rect 30101 40579 30159 40585
rect 30101 40576 30113 40579
rect 28552 40548 30113 40576
rect 30101 40545 30113 40548
rect 30147 40545 30159 40579
rect 30101 40539 30159 40545
rect 29914 40508 29920 40520
rect 29875 40480 29920 40508
rect 29914 40468 29920 40480
rect 29972 40468 29978 40520
rect 28350 40440 28356 40452
rect 28184 40412 28356 40440
rect 28350 40400 28356 40412
rect 28408 40440 28414 40452
rect 28994 40440 29000 40452
rect 28408 40412 29000 40440
rect 28408 40400 28414 40412
rect 28994 40400 29000 40412
rect 29052 40400 29058 40452
rect 27488 40344 27752 40372
rect 27488 40332 27494 40344
rect 1104 40282 30820 40304
rect 1104 40230 10880 40282
rect 10932 40230 10944 40282
rect 10996 40230 11008 40282
rect 11060 40230 11072 40282
rect 11124 40230 11136 40282
rect 11188 40230 20811 40282
rect 20863 40230 20875 40282
rect 20927 40230 20939 40282
rect 20991 40230 21003 40282
rect 21055 40230 21067 40282
rect 21119 40230 30820 40282
rect 1104 40208 30820 40230
rect 1397 40171 1455 40177
rect 1397 40137 1409 40171
rect 1443 40168 1455 40171
rect 8662 40168 8668 40180
rect 1443 40140 2774 40168
rect 8623 40140 8668 40168
rect 1443 40137 1455 40140
rect 1397 40131 1455 40137
rect 2746 40100 2774 40140
rect 8662 40128 8668 40140
rect 8720 40128 8726 40180
rect 10318 40168 10324 40180
rect 9959 40140 10324 40168
rect 8481 40103 8539 40109
rect 8481 40100 8493 40103
rect 2746 40072 8493 40100
rect 8481 40069 8493 40072
rect 8527 40069 8539 40103
rect 9959 40100 9987 40140
rect 10318 40128 10324 40140
rect 10376 40128 10382 40180
rect 19978 40168 19984 40180
rect 19939 40140 19984 40168
rect 19978 40128 19984 40140
rect 20036 40128 20042 40180
rect 21091 40171 21149 40177
rect 21091 40137 21103 40171
rect 21137 40168 21149 40171
rect 22738 40168 22744 40180
rect 21137 40140 22140 40168
rect 22699 40140 22744 40168
rect 21137 40137 21149 40140
rect 21091 40131 21149 40137
rect 8481 40063 8539 40069
rect 9876 40072 9987 40100
rect 1578 40032 1584 40044
rect 1539 40004 1584 40032
rect 1578 39992 1584 40004
rect 1636 39992 1642 40044
rect 8297 40035 8355 40041
rect 8297 40001 8309 40035
rect 8343 40032 8355 40035
rect 8386 40032 8392 40044
rect 8343 40004 8392 40032
rect 8343 40001 8355 40004
rect 8297 39995 8355 40001
rect 8386 39992 8392 40004
rect 8444 39992 8450 40044
rect 9876 40041 9904 40072
rect 10134 40060 10140 40112
rect 10192 40060 10198 40112
rect 11977 40103 12035 40109
rect 11977 40069 11989 40103
rect 12023 40100 12035 40103
rect 12894 40100 12900 40112
rect 12023 40072 12900 40100
rect 12023 40069 12035 40072
rect 11977 40063 12035 40069
rect 12894 40060 12900 40072
rect 12952 40060 12958 40112
rect 15746 40060 15752 40112
rect 15804 40100 15810 40112
rect 15933 40103 15991 40109
rect 15933 40100 15945 40103
rect 15804 40072 15945 40100
rect 15804 40060 15810 40072
rect 15933 40069 15945 40072
rect 15979 40069 15991 40103
rect 17034 40100 17040 40112
rect 16995 40072 17040 40100
rect 15933 40063 15991 40069
rect 17034 40060 17040 40072
rect 17092 40060 17098 40112
rect 19702 40060 19708 40112
rect 19760 40100 19766 40112
rect 19797 40103 19855 40109
rect 19797 40100 19809 40103
rect 19760 40072 19809 40100
rect 19760 40060 19766 40072
rect 19797 40069 19809 40072
rect 19843 40069 19855 40103
rect 19797 40063 19855 40069
rect 20073 40103 20131 40109
rect 20073 40069 20085 40103
rect 20119 40100 20131 40103
rect 20438 40100 20444 40112
rect 20119 40072 20444 40100
rect 20119 40069 20131 40072
rect 20073 40063 20131 40069
rect 20438 40060 20444 40072
rect 20496 40060 20502 40112
rect 20993 40103 21051 40109
rect 20993 40069 21005 40103
rect 21039 40100 21051 40103
rect 21450 40100 21456 40112
rect 21039 40072 21456 40100
rect 21039 40069 21051 40072
rect 20993 40063 21051 40069
rect 21450 40060 21456 40072
rect 21508 40060 21514 40112
rect 21634 40100 21640 40112
rect 21560 40072 21640 40100
rect 9841 40035 9904 40041
rect 9841 40001 9853 40035
rect 9887 40004 9904 40035
rect 9934 40035 9992 40041
rect 9887 40001 9899 40004
rect 9841 39995 9899 40001
rect 9934 40001 9946 40035
rect 9980 40001 9992 40035
rect 10045 40035 10103 40041
rect 10045 40032 10057 40035
rect 9934 39995 9992 40001
rect 10041 40001 10057 40032
rect 10091 40001 10103 40035
rect 10152 40032 10180 40060
rect 10229 40035 10287 40041
rect 10229 40032 10241 40035
rect 10152 40004 10241 40032
rect 10041 39995 10103 40001
rect 10229 40001 10241 40004
rect 10275 40001 10287 40035
rect 21174 40032 21180 40044
rect 21135 40004 21180 40032
rect 10229 39995 10287 40001
rect 9858 39856 9864 39908
rect 9916 39896 9922 39908
rect 9959 39896 9987 39995
rect 10041 39964 10069 39995
rect 21174 39992 21180 40004
rect 21232 39992 21238 40044
rect 21269 40035 21327 40041
rect 21269 40001 21281 40035
rect 21315 40032 21327 40035
rect 21560 40032 21588 40072
rect 21634 40060 21640 40072
rect 21692 40060 21698 40112
rect 22112 40041 22140 40140
rect 22738 40128 22744 40140
rect 22796 40128 22802 40180
rect 23198 40168 23204 40180
rect 23159 40140 23204 40168
rect 23198 40128 23204 40140
rect 23256 40128 23262 40180
rect 26050 40128 26056 40180
rect 26108 40168 26114 40180
rect 26234 40168 26240 40180
rect 26108 40140 26240 40168
rect 26108 40128 26114 40140
rect 26234 40128 26240 40140
rect 26292 40128 26298 40180
rect 27249 40171 27307 40177
rect 27249 40137 27261 40171
rect 27295 40168 27307 40171
rect 27522 40168 27528 40180
rect 27295 40140 27528 40168
rect 27295 40137 27307 40140
rect 27249 40131 27307 40137
rect 27522 40128 27528 40140
rect 27580 40128 27586 40180
rect 27614 40128 27620 40180
rect 27672 40168 27678 40180
rect 27672 40140 27717 40168
rect 27672 40128 27678 40140
rect 22646 40060 22652 40112
rect 22704 40100 22710 40112
rect 24121 40103 24179 40109
rect 24121 40100 24133 40103
rect 22704 40072 24133 40100
rect 22704 40060 22710 40072
rect 24121 40069 24133 40072
rect 24167 40069 24179 40103
rect 28166 40100 28172 40112
rect 24121 40063 24179 40069
rect 26160 40072 28172 40100
rect 21315 40004 21588 40032
rect 22097 40035 22155 40041
rect 21315 40001 21327 40004
rect 21269 39995 21327 40001
rect 22097 40001 22109 40035
rect 22143 40001 22155 40035
rect 22097 39995 22155 40001
rect 22462 39992 22468 40044
rect 22520 40032 22526 40044
rect 22738 40032 22744 40044
rect 22520 40004 22744 40032
rect 22520 39992 22526 40004
rect 22738 39992 22744 40004
rect 22796 39992 22802 40044
rect 23385 40035 23443 40041
rect 23385 40001 23397 40035
rect 23431 40032 23443 40035
rect 23566 40032 23572 40044
rect 23431 40004 23572 40032
rect 23431 40001 23443 40004
rect 23385 39995 23443 40001
rect 23566 39992 23572 40004
rect 23624 40032 23630 40044
rect 24302 40032 24308 40044
rect 23624 40004 23888 40032
rect 24263 40004 24308 40032
rect 23624 39992 23630 40004
rect 10134 39964 10140 39976
rect 10041 39936 10140 39964
rect 10134 39924 10140 39936
rect 10192 39924 10198 39976
rect 23290 39924 23296 39976
rect 23348 39964 23354 39976
rect 23474 39964 23480 39976
rect 23348 39936 23480 39964
rect 23348 39924 23354 39936
rect 23474 39924 23480 39936
rect 23532 39964 23538 39976
rect 23661 39967 23719 39973
rect 23661 39964 23673 39967
rect 23532 39936 23673 39964
rect 23532 39924 23538 39936
rect 23661 39933 23673 39936
rect 23707 39933 23719 39967
rect 23860 39964 23888 40004
rect 24302 39992 24308 40004
rect 24360 39992 24366 40044
rect 26160 40041 26188 40072
rect 28166 40060 28172 40072
rect 28224 40060 28230 40112
rect 28534 40100 28540 40112
rect 28276 40072 28540 40100
rect 26145 40035 26203 40041
rect 26145 40001 26157 40035
rect 26191 40001 26203 40035
rect 27430 40032 27436 40044
rect 27391 40004 27436 40032
rect 26145 39995 26203 40001
rect 27430 39992 27436 40004
rect 27488 39992 27494 40044
rect 27709 40035 27767 40041
rect 27709 40001 27721 40035
rect 27755 40032 27767 40035
rect 28276 40032 28304 40072
rect 28534 40060 28540 40072
rect 28592 40100 28598 40112
rect 28810 40100 28816 40112
rect 28592 40072 28816 40100
rect 28592 40060 28598 40072
rect 28810 40060 28816 40072
rect 28868 40060 28874 40112
rect 27755 40004 28304 40032
rect 27755 40001 27767 40004
rect 27709 39995 27767 40001
rect 28350 39992 28356 40044
rect 28408 40032 28414 40044
rect 28445 40035 28503 40041
rect 28445 40032 28457 40035
rect 28408 40004 28457 40032
rect 28408 39992 28414 40004
rect 28445 40001 28457 40004
rect 28491 40001 28503 40035
rect 28445 39995 28503 40001
rect 29825 40035 29883 40041
rect 29825 40001 29837 40035
rect 29871 40001 29883 40035
rect 29825 39995 29883 40001
rect 24489 39967 24547 39973
rect 24489 39964 24501 39967
rect 23860 39936 24501 39964
rect 23661 39927 23719 39933
rect 24489 39933 24501 39936
rect 24535 39933 24547 39967
rect 28166 39964 28172 39976
rect 28127 39936 28172 39964
rect 24489 39927 24547 39933
rect 28166 39924 28172 39936
rect 28224 39924 28230 39976
rect 10594 39896 10600 39908
rect 9916 39868 10600 39896
rect 9916 39856 9922 39868
rect 10594 39856 10600 39868
rect 10652 39856 10658 39908
rect 18230 39856 18236 39908
rect 18288 39896 18294 39908
rect 18325 39899 18383 39905
rect 18325 39896 18337 39899
rect 18288 39868 18337 39896
rect 18288 39856 18294 39868
rect 18325 39865 18337 39868
rect 18371 39865 18383 39899
rect 18325 39859 18383 39865
rect 21450 39856 21456 39908
rect 21508 39896 21514 39908
rect 22094 39896 22100 39908
rect 21508 39868 22100 39896
rect 21508 39856 21514 39868
rect 22094 39856 22100 39868
rect 22152 39856 22158 39908
rect 24762 39896 24768 39908
rect 23400 39868 24768 39896
rect 9585 39831 9643 39837
rect 9585 39797 9597 39831
rect 9631 39828 9643 39831
rect 9950 39828 9956 39840
rect 9631 39800 9956 39828
rect 9631 39797 9643 39800
rect 9585 39791 9643 39797
rect 9950 39788 9956 39800
rect 10008 39788 10014 39840
rect 11514 39788 11520 39840
rect 11572 39828 11578 39840
rect 12069 39831 12127 39837
rect 12069 39828 12081 39831
rect 11572 39800 12081 39828
rect 11572 39788 11578 39800
rect 12069 39797 12081 39800
rect 12115 39828 12127 39831
rect 12158 39828 12164 39840
rect 12115 39800 12164 39828
rect 12115 39797 12127 39800
rect 12069 39791 12127 39797
rect 12158 39788 12164 39800
rect 12216 39788 12222 39840
rect 16025 39831 16083 39837
rect 16025 39797 16037 39831
rect 16071 39828 16083 39831
rect 16574 39828 16580 39840
rect 16071 39800 16580 39828
rect 16071 39797 16083 39800
rect 16025 39791 16083 39797
rect 16574 39788 16580 39800
rect 16632 39788 16638 39840
rect 19521 39831 19579 39837
rect 19521 39797 19533 39831
rect 19567 39828 19579 39831
rect 19610 39828 19616 39840
rect 19567 39800 19616 39828
rect 19567 39797 19579 39800
rect 19521 39791 19579 39797
rect 19610 39788 19616 39800
rect 19668 39788 19674 39840
rect 21818 39788 21824 39840
rect 21876 39828 21882 39840
rect 23400 39828 23428 39868
rect 24762 39856 24768 39868
rect 24820 39856 24826 39908
rect 26329 39899 26387 39905
rect 26329 39865 26341 39899
rect 26375 39896 26387 39899
rect 27614 39896 27620 39908
rect 26375 39868 27620 39896
rect 26375 39865 26387 39868
rect 26329 39859 26387 39865
rect 27614 39856 27620 39868
rect 27672 39856 27678 39908
rect 21876 39800 23428 39828
rect 21876 39788 21882 39800
rect 23474 39788 23480 39840
rect 23532 39828 23538 39840
rect 23569 39831 23627 39837
rect 23569 39828 23581 39831
rect 23532 39800 23581 39828
rect 23532 39788 23538 39800
rect 23569 39797 23581 39800
rect 23615 39828 23627 39831
rect 24578 39828 24584 39840
rect 23615 39800 24584 39828
rect 23615 39797 23627 39800
rect 23569 39791 23627 39797
rect 24578 39788 24584 39800
rect 24636 39788 24642 39840
rect 24670 39788 24676 39840
rect 24728 39828 24734 39840
rect 25130 39828 25136 39840
rect 24728 39800 25136 39828
rect 24728 39788 24734 39800
rect 25130 39788 25136 39800
rect 25188 39788 25194 39840
rect 27522 39788 27528 39840
rect 27580 39828 27586 39840
rect 29840 39828 29868 39995
rect 29914 39856 29920 39908
rect 29972 39896 29978 39908
rect 30190 39896 30196 39908
rect 29972 39868 30196 39896
rect 29972 39856 29978 39868
rect 30190 39856 30196 39868
rect 30248 39856 30254 39908
rect 30006 39828 30012 39840
rect 27580 39800 29868 39828
rect 29967 39800 30012 39828
rect 27580 39788 27586 39800
rect 30006 39788 30012 39800
rect 30064 39788 30070 39840
rect 1104 39738 30820 39760
rect 1104 39686 5915 39738
rect 5967 39686 5979 39738
rect 6031 39686 6043 39738
rect 6095 39686 6107 39738
rect 6159 39686 6171 39738
rect 6223 39686 15846 39738
rect 15898 39686 15910 39738
rect 15962 39686 15974 39738
rect 16026 39686 16038 39738
rect 16090 39686 16102 39738
rect 16154 39686 25776 39738
rect 25828 39686 25840 39738
rect 25892 39686 25904 39738
rect 25956 39686 25968 39738
rect 26020 39686 26032 39738
rect 26084 39686 30820 39738
rect 1104 39664 30820 39686
rect 11882 39584 11888 39636
rect 11940 39624 11946 39636
rect 12989 39627 13047 39633
rect 12989 39624 13001 39627
rect 11940 39596 13001 39624
rect 11940 39584 11946 39596
rect 12989 39593 13001 39596
rect 13035 39624 13047 39627
rect 13906 39624 13912 39636
rect 13035 39596 13912 39624
rect 13035 39593 13047 39596
rect 12989 39587 13047 39593
rect 13906 39584 13912 39596
rect 13964 39584 13970 39636
rect 14274 39624 14280 39636
rect 14235 39596 14280 39624
rect 14274 39584 14280 39596
rect 14332 39584 14338 39636
rect 16209 39627 16267 39633
rect 16209 39593 16221 39627
rect 16255 39624 16267 39627
rect 16942 39624 16948 39636
rect 16255 39596 16948 39624
rect 16255 39593 16267 39596
rect 16209 39587 16267 39593
rect 16942 39584 16948 39596
rect 17000 39584 17006 39636
rect 18690 39624 18696 39636
rect 17052 39596 18276 39624
rect 18651 39596 18696 39624
rect 13538 39516 13544 39568
rect 13596 39556 13602 39568
rect 17052 39556 17080 39596
rect 13596 39528 17080 39556
rect 18248 39556 18276 39596
rect 18690 39584 18696 39596
rect 18748 39584 18754 39636
rect 19306 39596 22094 39624
rect 19306 39556 19334 39596
rect 18248 39528 19334 39556
rect 13596 39516 13602 39528
rect 10594 39488 10600 39500
rect 10555 39460 10600 39488
rect 10594 39448 10600 39460
rect 10652 39448 10658 39500
rect 16574 39488 16580 39500
rect 16535 39460 16580 39488
rect 16574 39448 16580 39460
rect 16632 39448 16638 39500
rect 20714 39448 20720 39500
rect 20772 39488 20778 39500
rect 20901 39491 20959 39497
rect 20901 39488 20913 39491
rect 20772 39460 20913 39488
rect 20772 39448 20778 39460
rect 20901 39457 20913 39460
rect 20947 39457 20959 39491
rect 22066 39488 22094 39596
rect 23198 39584 23204 39636
rect 23256 39624 23262 39636
rect 23385 39627 23443 39633
rect 23385 39624 23397 39627
rect 23256 39596 23397 39624
rect 23256 39584 23262 39596
rect 23385 39593 23397 39596
rect 23431 39593 23443 39627
rect 23385 39587 23443 39593
rect 26602 39584 26608 39636
rect 26660 39624 26666 39636
rect 26973 39627 27031 39633
rect 26973 39624 26985 39627
rect 26660 39596 26985 39624
rect 26660 39584 26666 39596
rect 26973 39593 26985 39596
rect 27019 39593 27031 39627
rect 26973 39587 27031 39593
rect 28258 39584 28264 39636
rect 28316 39624 28322 39636
rect 28902 39624 28908 39636
rect 28316 39596 28908 39624
rect 28316 39584 28322 39596
rect 28902 39584 28908 39596
rect 28960 39584 28966 39636
rect 24486 39516 24492 39568
rect 24544 39556 24550 39568
rect 24544 39528 24900 39556
rect 24544 39516 24550 39528
rect 24872 39497 24900 39528
rect 24765 39491 24823 39497
rect 24765 39488 24777 39491
rect 22066 39460 24777 39488
rect 20901 39451 20959 39457
rect 24765 39457 24777 39460
rect 24811 39457 24823 39491
rect 24765 39451 24823 39457
rect 24857 39491 24915 39497
rect 24857 39457 24869 39491
rect 24903 39457 24915 39491
rect 24857 39451 24915 39457
rect 1578 39420 1584 39432
rect 1539 39392 1584 39420
rect 1578 39380 1584 39392
rect 1636 39380 1642 39432
rect 10321 39423 10379 39429
rect 10321 39389 10333 39423
rect 10367 39420 10379 39423
rect 11422 39420 11428 39432
rect 10367 39392 11428 39420
rect 10367 39389 10379 39392
rect 10321 39383 10379 39389
rect 11422 39380 11428 39392
rect 11480 39380 11486 39432
rect 11606 39420 11612 39432
rect 11567 39392 11612 39420
rect 11606 39380 11612 39392
rect 11664 39380 11670 39432
rect 15010 39380 15016 39432
rect 15068 39420 15074 39432
rect 17586 39429 17592 39432
rect 17313 39423 17371 39429
rect 15068 39392 15332 39420
rect 15068 39380 15074 39392
rect 11698 39312 11704 39364
rect 11756 39352 11762 39364
rect 11854 39355 11912 39361
rect 11854 39352 11866 39355
rect 11756 39324 11866 39352
rect 11756 39312 11762 39324
rect 11854 39321 11866 39324
rect 11900 39321 11912 39355
rect 14182 39352 14188 39364
rect 14143 39324 14188 39352
rect 11854 39315 11912 39321
rect 14182 39312 14188 39324
rect 14240 39312 14246 39364
rect 15304 39361 15332 39392
rect 17313 39389 17325 39423
rect 17359 39420 17371 39423
rect 17359 39392 17540 39420
rect 17359 39389 17371 39392
rect 17313 39383 17371 39389
rect 15105 39355 15163 39361
rect 15105 39321 15117 39355
rect 15151 39321 15163 39355
rect 15105 39315 15163 39321
rect 15289 39355 15347 39361
rect 15289 39321 15301 39355
rect 15335 39352 15347 39355
rect 15378 39352 15384 39364
rect 15335 39324 15384 39352
rect 15335 39321 15347 39324
rect 15289 39315 15347 39321
rect 1397 39287 1455 39293
rect 1397 39253 1409 39287
rect 1443 39284 1455 39287
rect 8570 39284 8576 39296
rect 1443 39256 8576 39284
rect 1443 39253 1455 39256
rect 1397 39247 1455 39253
rect 8570 39244 8576 39256
rect 8628 39244 8634 39296
rect 10042 39244 10048 39296
rect 10100 39284 10106 39296
rect 12158 39284 12164 39296
rect 10100 39256 12164 39284
rect 10100 39244 10106 39256
rect 12158 39244 12164 39256
rect 12216 39244 12222 39296
rect 12710 39244 12716 39296
rect 12768 39284 12774 39296
rect 15120 39284 15148 39315
rect 15378 39312 15384 39324
rect 15436 39312 15442 39364
rect 16761 39355 16819 39361
rect 16761 39321 16773 39355
rect 16807 39352 16819 39355
rect 17402 39352 17408 39364
rect 16807 39324 17408 39352
rect 16807 39321 16819 39324
rect 16761 39315 16819 39321
rect 17402 39312 17408 39324
rect 17460 39312 17466 39364
rect 15654 39284 15660 39296
rect 12768 39256 15660 39284
rect 12768 39244 12774 39256
rect 15654 39244 15660 39256
rect 15712 39244 15718 39296
rect 16669 39287 16727 39293
rect 16669 39253 16681 39287
rect 16715 39284 16727 39287
rect 17218 39284 17224 39296
rect 16715 39256 17224 39284
rect 16715 39253 16727 39256
rect 16669 39247 16727 39253
rect 17218 39244 17224 39256
rect 17276 39244 17282 39296
rect 17512 39284 17540 39392
rect 17580 39383 17592 39429
rect 17644 39420 17650 39432
rect 21168 39423 21226 39429
rect 17644 39392 17680 39420
rect 17586 39380 17592 39383
rect 17644 39380 17650 39392
rect 21168 39389 21180 39423
rect 21214 39420 21226 39423
rect 22922 39420 22928 39432
rect 21214 39392 22928 39420
rect 21214 39389 21226 39392
rect 21168 39383 21226 39389
rect 22922 39380 22928 39392
rect 22980 39380 22986 39432
rect 23290 39420 23296 39432
rect 23251 39392 23296 39420
rect 23290 39380 23296 39392
rect 23348 39380 23354 39432
rect 24578 39420 24584 39432
rect 24539 39392 24584 39420
rect 24578 39380 24584 39392
rect 24636 39380 24642 39432
rect 24673 39423 24731 39429
rect 24673 39389 24685 39423
rect 24719 39389 24731 39423
rect 24673 39383 24731 39389
rect 18690 39312 18696 39364
rect 18748 39352 18754 39364
rect 19705 39355 19763 39361
rect 19705 39352 19717 39355
rect 18748 39324 19717 39352
rect 18748 39312 18754 39324
rect 19705 39321 19717 39324
rect 19751 39321 19763 39355
rect 19705 39315 19763 39321
rect 22646 39312 22652 39364
rect 22704 39352 22710 39364
rect 23109 39355 23167 39361
rect 23109 39352 23121 39355
rect 22704 39324 23121 39352
rect 22704 39312 22710 39324
rect 23109 39321 23121 39324
rect 23155 39321 23167 39355
rect 24688 39352 24716 39383
rect 26234 39380 26240 39432
rect 26292 39420 26298 39432
rect 26789 39423 26847 39429
rect 26789 39420 26801 39423
rect 26292 39392 26801 39420
rect 26292 39380 26298 39392
rect 26789 39389 26801 39392
rect 26835 39389 26847 39423
rect 27982 39420 27988 39432
rect 27943 39392 27988 39420
rect 26789 39383 26847 39389
rect 27982 39380 27988 39392
rect 28040 39380 28046 39432
rect 28721 39423 28779 39429
rect 28721 39389 28733 39423
rect 28767 39420 28779 39423
rect 29454 39420 29460 39432
rect 28767 39392 29460 39420
rect 28767 39389 28779 39392
rect 28721 39383 28779 39389
rect 29454 39380 29460 39392
rect 29512 39380 29518 39432
rect 29825 39423 29883 39429
rect 29825 39389 29837 39423
rect 29871 39389 29883 39423
rect 29825 39383 29883 39389
rect 24762 39352 24768 39364
rect 24688 39324 24768 39352
rect 23109 39315 23167 39321
rect 24762 39312 24768 39324
rect 24820 39312 24826 39364
rect 25866 39312 25872 39364
rect 25924 39352 25930 39364
rect 29840 39352 29868 39383
rect 25924 39324 29868 39352
rect 25924 39312 25930 39324
rect 17862 39284 17868 39296
rect 17512 39256 17868 39284
rect 17862 39244 17868 39256
rect 17920 39244 17926 39296
rect 18414 39244 18420 39296
rect 18472 39284 18478 39296
rect 19797 39287 19855 39293
rect 19797 39284 19809 39287
rect 18472 39256 19809 39284
rect 18472 39244 18478 39256
rect 19797 39253 19809 39256
rect 19843 39284 19855 39287
rect 20162 39284 20168 39296
rect 19843 39256 20168 39284
rect 19843 39253 19855 39256
rect 19797 39247 19855 39253
rect 20162 39244 20168 39256
rect 20220 39244 20226 39296
rect 22278 39284 22284 39296
rect 22239 39256 22284 39284
rect 22278 39244 22284 39256
rect 22336 39244 22342 39296
rect 24397 39287 24455 39293
rect 24397 39253 24409 39287
rect 24443 39284 24455 39287
rect 24670 39284 24676 39296
rect 24443 39256 24676 39284
rect 24443 39253 24455 39256
rect 24397 39247 24455 39253
rect 24670 39244 24676 39256
rect 24728 39244 24734 39296
rect 28166 39284 28172 39296
rect 28127 39256 28172 39284
rect 28166 39244 28172 39256
rect 28224 39244 28230 39296
rect 28902 39284 28908 39296
rect 28863 39256 28908 39284
rect 28902 39244 28908 39256
rect 28960 39244 28966 39296
rect 29178 39244 29184 39296
rect 29236 39284 29242 39296
rect 29638 39284 29644 39296
rect 29236 39256 29644 39284
rect 29236 39244 29242 39256
rect 29638 39244 29644 39256
rect 29696 39244 29702 39296
rect 30009 39287 30067 39293
rect 30009 39253 30021 39287
rect 30055 39284 30067 39287
rect 30098 39284 30104 39296
rect 30055 39256 30104 39284
rect 30055 39253 30067 39256
rect 30009 39247 30067 39253
rect 30098 39244 30104 39256
rect 30156 39244 30162 39296
rect 1104 39194 30820 39216
rect 1104 39142 10880 39194
rect 10932 39142 10944 39194
rect 10996 39142 11008 39194
rect 11060 39142 11072 39194
rect 11124 39142 11136 39194
rect 11188 39142 20811 39194
rect 20863 39142 20875 39194
rect 20927 39142 20939 39194
rect 20991 39142 21003 39194
rect 21055 39142 21067 39194
rect 21119 39142 30820 39194
rect 1104 39120 30820 39142
rect 11517 39083 11575 39089
rect 11517 39049 11529 39083
rect 11563 39080 11575 39083
rect 11698 39080 11704 39092
rect 11563 39052 11704 39080
rect 11563 39049 11575 39052
rect 11517 39043 11575 39049
rect 11698 39040 11704 39052
rect 11756 39040 11762 39092
rect 11882 39040 11888 39092
rect 11940 39040 11946 39092
rect 12805 39083 12863 39089
rect 12805 39049 12817 39083
rect 12851 39080 12863 39083
rect 17218 39080 17224 39092
rect 12851 39052 14381 39080
rect 17179 39052 17224 39080
rect 12851 39049 12863 39052
rect 12805 39043 12863 39049
rect 8386 39012 8392 39024
rect 8347 38984 8392 39012
rect 8386 38972 8392 38984
rect 8444 38972 8450 39024
rect 8570 39012 8576 39024
rect 8531 38984 8576 39012
rect 8570 38972 8576 38984
rect 8628 38972 8634 39024
rect 11900 39012 11928 39040
rect 12526 39012 12532 39024
rect 11808 38984 11928 39012
rect 12084 38984 12532 39012
rect 1578 38944 1584 38956
rect 1539 38916 1584 38944
rect 1578 38904 1584 38916
rect 1636 38904 1642 38956
rect 11808 38953 11836 38984
rect 11773 38947 11836 38953
rect 11773 38913 11785 38947
rect 11819 38916 11836 38947
rect 11882 38947 11940 38953
rect 11819 38913 11831 38916
rect 11773 38907 11831 38913
rect 11882 38913 11894 38947
rect 11928 38913 11940 38947
rect 11882 38907 11940 38913
rect 11998 38947 12056 38953
rect 11998 38913 12010 38947
rect 12044 38944 12056 38947
rect 12084 38944 12112 38984
rect 12526 38972 12532 38984
rect 12584 39012 12590 39024
rect 14353 39021 14381 39052
rect 17218 39040 17224 39052
rect 17276 39080 17282 39092
rect 18506 39080 18512 39092
rect 17276 39052 18512 39080
rect 17276 39040 17282 39052
rect 18506 39040 18512 39052
rect 18564 39040 18570 39092
rect 18785 39083 18843 39089
rect 18785 39049 18797 39083
rect 18831 39049 18843 39083
rect 22646 39080 22652 39092
rect 18785 39043 18843 39049
rect 20916 39052 22652 39080
rect 14338 39015 14396 39021
rect 12584 38984 13400 39012
rect 12584 38972 12590 38984
rect 12044 38916 12112 38944
rect 12044 38913 12056 38916
rect 11998 38907 12056 38913
rect 11900 38876 11928 38907
rect 12158 38904 12164 38956
rect 12216 38944 12222 38956
rect 12216 38916 12261 38944
rect 12216 38904 12222 38916
rect 12986 38904 12992 38956
rect 13044 38928 13050 38956
rect 13081 38947 13139 38953
rect 13081 38928 13093 38947
rect 13044 38913 13093 38928
rect 13127 38913 13139 38947
rect 13044 38907 13139 38913
rect 13170 38947 13228 38953
rect 13170 38913 13182 38947
rect 13216 38913 13228 38947
rect 13170 38907 13228 38913
rect 13265 38947 13323 38953
rect 13372 38947 13400 38984
rect 14338 38981 14350 39015
rect 14384 38981 14396 39015
rect 14338 38975 14396 38981
rect 16574 38972 16580 39024
rect 16632 39012 16638 39024
rect 17037 39015 17095 39021
rect 17037 39012 17049 39015
rect 16632 38984 17049 39012
rect 16632 38972 16638 38984
rect 17037 38981 17049 38984
rect 17083 38981 17095 39015
rect 17037 38975 17095 38981
rect 17862 38972 17868 39024
rect 17920 39012 17926 39024
rect 18800 39012 18828 39043
rect 19518 39012 19524 39024
rect 17920 38984 18828 39012
rect 19479 38984 19524 39012
rect 17920 38972 17926 38984
rect 19518 38972 19524 38984
rect 19576 38972 19582 39024
rect 20806 39012 20812 39024
rect 20767 38984 20812 39012
rect 20806 38972 20812 38984
rect 20864 38972 20870 39024
rect 20916 39021 20944 39052
rect 22646 39040 22652 39052
rect 22704 39040 22710 39092
rect 23566 39040 23572 39092
rect 23624 39080 23630 39092
rect 24762 39080 24768 39092
rect 23624 39052 24768 39080
rect 23624 39040 23630 39052
rect 24762 39040 24768 39052
rect 24820 39080 24826 39092
rect 24857 39083 24915 39089
rect 24857 39080 24869 39083
rect 24820 39052 24869 39080
rect 24820 39040 24826 39052
rect 24857 39049 24869 39052
rect 24903 39049 24915 39083
rect 24857 39043 24915 39049
rect 24949 39083 25007 39089
rect 24949 39049 24961 39083
rect 24995 39080 25007 39083
rect 25958 39080 25964 39092
rect 24995 39052 25964 39080
rect 24995 39049 25007 39052
rect 24949 39043 25007 39049
rect 20901 39015 20959 39021
rect 20901 38981 20913 39015
rect 20947 38981 20959 39015
rect 20901 38975 20959 38981
rect 23014 38972 23020 39024
rect 23072 39012 23078 39024
rect 24964 39012 24992 39043
rect 25958 39040 25964 39052
rect 26016 39040 26022 39092
rect 26050 39040 26056 39092
rect 26108 39080 26114 39092
rect 27157 39083 27215 39089
rect 27157 39080 27169 39083
rect 26108 39052 27169 39080
rect 26108 39040 26114 39052
rect 27157 39049 27169 39052
rect 27203 39049 27215 39083
rect 27157 39043 27215 39049
rect 28350 39040 28356 39092
rect 28408 39080 28414 39092
rect 28626 39080 28632 39092
rect 28408 39052 28632 39080
rect 28408 39040 28414 39052
rect 28626 39040 28632 39052
rect 28684 39040 28690 39092
rect 23072 38984 24992 39012
rect 23072 38972 23078 38984
rect 28994 38972 29000 39024
rect 29052 39012 29058 39024
rect 29730 39012 29736 39024
rect 29052 38984 29736 39012
rect 29052 38972 29058 38984
rect 29730 38972 29736 38984
rect 29788 38972 29794 39024
rect 13265 38913 13277 38947
rect 13311 38919 13400 38947
rect 13461 38947 13519 38953
rect 13311 38913 13323 38919
rect 13265 38907 13323 38913
rect 13461 38913 13473 38947
rect 13507 38913 13519 38947
rect 13461 38907 13519 38913
rect 13044 38904 13124 38907
rect 13009 38900 13124 38904
rect 11900 38848 12204 38876
rect 12176 38820 12204 38848
rect 1397 38811 1455 38817
rect 1397 38777 1409 38811
rect 1443 38808 1455 38811
rect 9030 38808 9036 38820
rect 1443 38780 9036 38808
rect 1443 38777 1455 38780
rect 1397 38771 1455 38777
rect 9030 38768 9036 38780
rect 9088 38768 9094 38820
rect 12158 38768 12164 38820
rect 12216 38808 12222 38820
rect 13188 38808 13216 38907
rect 13464 38820 13492 38907
rect 16298 38904 16304 38956
rect 16356 38944 16362 38956
rect 17957 38947 18015 38953
rect 17957 38944 17969 38947
rect 16356 38916 17969 38944
rect 16356 38904 16362 38916
rect 17957 38913 17969 38916
rect 18003 38944 18015 38947
rect 18414 38944 18420 38956
rect 18003 38916 18420 38944
rect 18003 38913 18015 38916
rect 17957 38907 18015 38913
rect 18414 38904 18420 38916
rect 18472 38904 18478 38956
rect 18601 38947 18659 38953
rect 18601 38913 18613 38947
rect 18647 38913 18659 38947
rect 18601 38907 18659 38913
rect 19337 38947 19395 38953
rect 19337 38913 19349 38947
rect 19383 38944 19395 38947
rect 20070 38944 20076 38956
rect 19383 38916 20076 38944
rect 19383 38913 19395 38916
rect 19337 38907 19395 38913
rect 14090 38876 14096 38888
rect 14051 38848 14096 38876
rect 14090 38836 14096 38848
rect 14148 38836 14154 38888
rect 17313 38879 17371 38885
rect 17313 38845 17325 38879
rect 17359 38876 17371 38879
rect 17402 38876 17408 38888
rect 17359 38848 17408 38876
rect 17359 38845 17371 38848
rect 17313 38839 17371 38845
rect 17402 38836 17408 38848
rect 17460 38836 17466 38888
rect 12216 38780 13216 38808
rect 12216 38768 12222 38780
rect 13446 38768 13452 38820
rect 13504 38768 13510 38820
rect 16761 38811 16819 38817
rect 16761 38777 16773 38811
rect 16807 38808 16819 38811
rect 18616 38808 18644 38907
rect 20070 38904 20076 38916
rect 20128 38904 20134 38956
rect 20162 38904 20168 38956
rect 20220 38944 20226 38956
rect 22281 38947 22339 38953
rect 20220 38916 22232 38944
rect 20220 38904 20226 38916
rect 20809 38879 20867 38885
rect 20809 38845 20821 38879
rect 20855 38845 20867 38879
rect 22204 38876 22232 38916
rect 22281 38913 22293 38947
rect 22327 38944 22339 38947
rect 22327 38916 24532 38944
rect 22327 38913 22339 38916
rect 22281 38907 22339 38913
rect 23017 38879 23075 38885
rect 23017 38876 23029 38879
rect 22204 38848 23029 38876
rect 20809 38839 20867 38845
rect 23017 38845 23029 38848
rect 23063 38845 23075 38879
rect 23017 38839 23075 38845
rect 23293 38879 23351 38885
rect 23293 38845 23305 38879
rect 23339 38876 23351 38879
rect 23566 38876 23572 38888
rect 23339 38848 23572 38876
rect 23339 38845 23351 38848
rect 23293 38839 23351 38845
rect 16807 38780 18644 38808
rect 20824 38808 20852 38839
rect 23566 38836 23572 38848
rect 23624 38836 23630 38888
rect 24504 38876 24532 38916
rect 24578 38904 24584 38956
rect 24636 38944 24642 38956
rect 24765 38947 24823 38953
rect 24765 38944 24777 38947
rect 24636 38916 24777 38944
rect 24636 38904 24642 38916
rect 24765 38913 24777 38916
rect 24811 38913 24823 38947
rect 24765 38907 24823 38913
rect 24946 38904 24952 38956
rect 25004 38944 25010 38956
rect 25133 38947 25191 38953
rect 25133 38944 25145 38947
rect 25004 38916 25145 38944
rect 25004 38904 25010 38916
rect 25133 38913 25145 38916
rect 25179 38913 25191 38947
rect 25133 38907 25191 38913
rect 25222 38904 25228 38956
rect 25280 38944 25286 38956
rect 26973 38947 27031 38953
rect 26973 38944 26985 38947
rect 25280 38916 26985 38944
rect 25280 38904 25286 38916
rect 26973 38913 26985 38916
rect 27019 38913 27031 38947
rect 26973 38907 27031 38913
rect 27522 38904 27528 38956
rect 27580 38944 27586 38956
rect 28353 38947 28411 38953
rect 28353 38944 28365 38947
rect 27580 38916 28365 38944
rect 27580 38904 27586 38916
rect 28353 38913 28365 38916
rect 28399 38913 28411 38947
rect 28353 38907 28411 38913
rect 29089 38947 29147 38953
rect 29089 38913 29101 38947
rect 29135 38913 29147 38947
rect 29822 38944 29828 38956
rect 29783 38916 29828 38944
rect 29089 38907 29147 38913
rect 25240 38876 25268 38904
rect 24504 38848 25268 38876
rect 25866 38836 25872 38888
rect 25924 38876 25930 38888
rect 29104 38876 29132 38907
rect 29822 38904 29828 38916
rect 29880 38904 29886 38956
rect 25924 38848 29132 38876
rect 25924 38836 25930 38848
rect 21082 38808 21088 38820
rect 20824 38780 21088 38808
rect 16807 38777 16819 38780
rect 16761 38771 16819 38777
rect 21082 38768 21088 38780
rect 21140 38768 21146 38820
rect 22922 38768 22928 38820
rect 22980 38808 22986 38820
rect 23658 38808 23664 38820
rect 22980 38780 23664 38808
rect 22980 38768 22986 38780
rect 23658 38768 23664 38780
rect 23716 38768 23722 38820
rect 24581 38811 24639 38817
rect 24581 38777 24593 38811
rect 24627 38777 24639 38811
rect 24581 38771 24639 38777
rect 8757 38743 8815 38749
rect 8757 38709 8769 38743
rect 8803 38740 8815 38743
rect 11790 38740 11796 38752
rect 8803 38712 11796 38740
rect 8803 38709 8815 38712
rect 8757 38703 8815 38709
rect 11790 38700 11796 38712
rect 11848 38700 11854 38752
rect 12986 38700 12992 38752
rect 13044 38740 13050 38752
rect 15473 38743 15531 38749
rect 15473 38740 15485 38743
rect 13044 38712 15485 38740
rect 13044 38700 13050 38712
rect 15473 38709 15485 38712
rect 15519 38740 15531 38743
rect 15562 38740 15568 38752
rect 15519 38712 15568 38740
rect 15519 38709 15531 38712
rect 15473 38703 15531 38709
rect 15562 38700 15568 38712
rect 15620 38700 15626 38752
rect 17402 38700 17408 38752
rect 17460 38740 17466 38752
rect 18049 38743 18107 38749
rect 18049 38740 18061 38743
rect 17460 38712 18061 38740
rect 17460 38700 17466 38712
rect 18049 38709 18061 38712
rect 18095 38709 18107 38743
rect 18049 38703 18107 38709
rect 19334 38700 19340 38752
rect 19392 38740 19398 38752
rect 20349 38743 20407 38749
rect 20349 38740 20361 38743
rect 19392 38712 20361 38740
rect 19392 38700 19398 38712
rect 20349 38709 20361 38712
rect 20395 38709 20407 38743
rect 20349 38703 20407 38709
rect 22465 38743 22523 38749
rect 22465 38709 22477 38743
rect 22511 38740 22523 38743
rect 22738 38740 22744 38752
rect 22511 38712 22744 38740
rect 22511 38709 22523 38712
rect 22465 38703 22523 38709
rect 22738 38700 22744 38712
rect 22796 38700 22802 38752
rect 23842 38700 23848 38752
rect 23900 38740 23906 38752
rect 24596 38740 24624 38771
rect 24946 38768 24952 38820
rect 25004 38808 25010 38820
rect 26050 38808 26056 38820
rect 25004 38780 26056 38808
rect 25004 38768 25010 38780
rect 26050 38768 26056 38780
rect 26108 38768 26114 38820
rect 23900 38712 24624 38740
rect 28537 38743 28595 38749
rect 23900 38700 23906 38712
rect 28537 38709 28549 38743
rect 28583 38740 28595 38743
rect 28626 38740 28632 38752
rect 28583 38712 28632 38740
rect 28583 38709 28595 38712
rect 28537 38703 28595 38709
rect 28626 38700 28632 38712
rect 28684 38700 28690 38752
rect 29273 38743 29331 38749
rect 29273 38709 29285 38743
rect 29319 38740 29331 38743
rect 29362 38740 29368 38752
rect 29319 38712 29368 38740
rect 29319 38709 29331 38712
rect 29273 38703 29331 38709
rect 29362 38700 29368 38712
rect 29420 38700 29426 38752
rect 29914 38700 29920 38752
rect 29972 38740 29978 38752
rect 30009 38743 30067 38749
rect 30009 38740 30021 38743
rect 29972 38712 30021 38740
rect 29972 38700 29978 38712
rect 30009 38709 30021 38712
rect 30055 38709 30067 38743
rect 30009 38703 30067 38709
rect 1104 38650 30820 38672
rect 1104 38598 5915 38650
rect 5967 38598 5979 38650
rect 6031 38598 6043 38650
rect 6095 38598 6107 38650
rect 6159 38598 6171 38650
rect 6223 38598 15846 38650
rect 15898 38598 15910 38650
rect 15962 38598 15974 38650
rect 16026 38598 16038 38650
rect 16090 38598 16102 38650
rect 16154 38598 25776 38650
rect 25828 38598 25840 38650
rect 25892 38598 25904 38650
rect 25956 38598 25968 38650
rect 26020 38598 26032 38650
rect 26084 38598 30820 38650
rect 1104 38576 30820 38598
rect 11057 38539 11115 38545
rect 11057 38505 11069 38539
rect 11103 38536 11115 38539
rect 11238 38536 11244 38548
rect 11103 38508 11244 38536
rect 11103 38505 11115 38508
rect 11057 38499 11115 38505
rect 11238 38496 11244 38508
rect 11296 38496 11302 38548
rect 17221 38539 17279 38545
rect 17221 38505 17233 38539
rect 17267 38536 17279 38539
rect 17678 38536 17684 38548
rect 17267 38508 17684 38536
rect 17267 38505 17279 38508
rect 17221 38499 17279 38505
rect 17678 38496 17684 38508
rect 17736 38496 17742 38548
rect 18046 38536 18052 38548
rect 18007 38508 18052 38536
rect 18046 38496 18052 38508
rect 18104 38496 18110 38548
rect 20441 38539 20499 38545
rect 20441 38505 20453 38539
rect 20487 38536 20499 38539
rect 20806 38536 20812 38548
rect 20487 38508 20812 38536
rect 20487 38505 20499 38508
rect 20441 38499 20499 38505
rect 20806 38496 20812 38508
rect 20864 38496 20870 38548
rect 21082 38536 21088 38548
rect 21043 38508 21088 38536
rect 21082 38496 21088 38508
rect 21140 38496 21146 38548
rect 22922 38496 22928 38548
rect 22980 38536 22986 38548
rect 25222 38536 25228 38548
rect 22980 38508 23888 38536
rect 22980 38496 22986 38508
rect 16482 38428 16488 38480
rect 16540 38468 16546 38480
rect 22186 38468 22192 38480
rect 16540 38440 22192 38468
rect 16540 38428 16546 38440
rect 22186 38428 22192 38440
rect 22244 38428 22250 38480
rect 11422 38360 11428 38412
rect 11480 38400 11486 38412
rect 11793 38403 11851 38409
rect 11793 38400 11805 38403
rect 11480 38372 11805 38400
rect 11480 38360 11486 38372
rect 11793 38369 11805 38372
rect 11839 38400 11851 38403
rect 12618 38400 12624 38412
rect 11839 38372 12624 38400
rect 11839 38369 11851 38372
rect 11793 38363 11851 38369
rect 12618 38360 12624 38372
rect 12676 38360 12682 38412
rect 16206 38360 16212 38412
rect 16264 38400 16270 38412
rect 22922 38400 22928 38412
rect 16264 38372 22928 38400
rect 16264 38360 16270 38372
rect 22922 38360 22928 38372
rect 22980 38360 22986 38412
rect 1578 38332 1584 38344
rect 1539 38304 1584 38332
rect 1578 38292 1584 38304
rect 1636 38292 1642 38344
rect 9677 38335 9735 38341
rect 9677 38301 9689 38335
rect 9723 38332 9735 38335
rect 9766 38332 9772 38344
rect 9723 38304 9772 38332
rect 9723 38301 9735 38304
rect 9677 38295 9735 38301
rect 9766 38292 9772 38304
rect 9824 38292 9830 38344
rect 9950 38341 9956 38344
rect 9944 38332 9956 38341
rect 9911 38304 9956 38332
rect 9944 38295 9956 38304
rect 9950 38292 9956 38295
rect 10008 38292 10014 38344
rect 12069 38335 12127 38341
rect 12069 38301 12081 38335
rect 12115 38332 12127 38335
rect 12158 38332 12164 38344
rect 12115 38304 12164 38332
rect 12115 38301 12127 38304
rect 12069 38295 12127 38301
rect 12158 38292 12164 38304
rect 12216 38292 12222 38344
rect 14090 38332 14096 38344
rect 14051 38304 14096 38332
rect 14090 38292 14096 38304
rect 14148 38292 14154 38344
rect 17954 38332 17960 38344
rect 14200 38304 17264 38332
rect 17915 38304 17960 38332
rect 12986 38224 12992 38276
rect 13044 38264 13050 38276
rect 14200 38264 14228 38304
rect 13044 38236 14228 38264
rect 14360 38267 14418 38273
rect 13044 38224 13050 38236
rect 14360 38233 14372 38267
rect 14406 38264 14418 38267
rect 16666 38264 16672 38276
rect 14406 38236 16672 38264
rect 14406 38233 14418 38236
rect 14360 38227 14418 38233
rect 16666 38224 16672 38236
rect 16724 38224 16730 38276
rect 17129 38267 17187 38273
rect 17129 38233 17141 38267
rect 17175 38233 17187 38267
rect 17236 38264 17264 38304
rect 17954 38292 17960 38304
rect 18012 38292 18018 38344
rect 19245 38335 19303 38341
rect 19245 38301 19257 38335
rect 19291 38332 19303 38335
rect 19334 38332 19340 38344
rect 19291 38304 19340 38332
rect 19291 38301 19303 38304
rect 19245 38295 19303 38301
rect 19334 38292 19340 38304
rect 19392 38292 19398 38344
rect 19978 38292 19984 38344
rect 20036 38332 20042 38344
rect 20349 38335 20407 38341
rect 20349 38332 20361 38335
rect 20036 38304 20361 38332
rect 20036 38292 20042 38304
rect 20349 38301 20361 38304
rect 20395 38301 20407 38335
rect 20349 38295 20407 38301
rect 20993 38335 21051 38341
rect 20993 38301 21005 38335
rect 21039 38332 21051 38335
rect 21542 38332 21548 38344
rect 21039 38304 21548 38332
rect 21039 38301 21051 38304
rect 20993 38295 21051 38301
rect 21542 38292 21548 38304
rect 21600 38292 21606 38344
rect 23032 38264 23060 38508
rect 23566 38428 23572 38480
rect 23624 38428 23630 38480
rect 23658 38428 23664 38480
rect 23716 38428 23722 38480
rect 23382 38360 23388 38412
rect 23440 38400 23446 38412
rect 23478 38403 23536 38409
rect 23478 38400 23490 38403
rect 23440 38372 23490 38400
rect 23440 38360 23446 38372
rect 23478 38369 23490 38372
rect 23524 38369 23536 38403
rect 23478 38363 23536 38369
rect 23584 38341 23612 38428
rect 23676 38400 23704 38428
rect 23753 38403 23811 38409
rect 23753 38400 23765 38403
rect 23676 38372 23765 38400
rect 23753 38369 23765 38372
rect 23799 38369 23811 38403
rect 23753 38363 23811 38369
rect 23569 38335 23627 38341
rect 23569 38301 23581 38335
rect 23615 38301 23627 38335
rect 23569 38295 23627 38301
rect 23661 38335 23719 38341
rect 23661 38301 23673 38335
rect 23707 38332 23719 38335
rect 23860 38332 23888 38508
rect 25056 38508 25228 38536
rect 24026 38360 24032 38412
rect 24084 38400 24090 38412
rect 24673 38403 24731 38409
rect 24084 38372 24532 38400
rect 24084 38360 24090 38372
rect 23707 38304 23888 38332
rect 24397 38335 24455 38341
rect 23707 38301 23719 38304
rect 23661 38295 23719 38301
rect 24397 38301 24409 38335
rect 24443 38301 24455 38335
rect 24504 38332 24532 38372
rect 24673 38369 24685 38403
rect 24719 38400 24731 38403
rect 25056 38400 25084 38508
rect 25222 38496 25228 38508
rect 25280 38496 25286 38548
rect 25498 38496 25504 38548
rect 25556 38536 25562 38548
rect 25556 38508 26096 38536
rect 25556 38496 25562 38508
rect 25516 38440 26004 38468
rect 24719 38372 25084 38400
rect 24719 38369 24731 38372
rect 24673 38363 24731 38369
rect 25222 38360 25228 38412
rect 25280 38400 25286 38412
rect 25516 38400 25544 38440
rect 25866 38400 25872 38412
rect 25280 38372 25544 38400
rect 25608 38372 25872 38400
rect 25280 38360 25286 38372
rect 25608 38332 25636 38372
rect 25866 38360 25872 38372
rect 25924 38360 25930 38412
rect 25976 38409 26004 38440
rect 25961 38403 26019 38409
rect 25961 38369 25973 38403
rect 26007 38369 26019 38403
rect 25961 38363 26019 38369
rect 24504 38304 25636 38332
rect 25685 38335 25743 38341
rect 24397 38295 24455 38301
rect 25685 38301 25697 38335
rect 25731 38334 25743 38335
rect 25774 38334 25780 38344
rect 25731 38306 25780 38334
rect 25731 38301 25743 38306
rect 25685 38295 25743 38301
rect 17236 38236 23060 38264
rect 17129 38227 17187 38233
rect 1397 38199 1455 38205
rect 1397 38165 1409 38199
rect 1443 38196 1455 38199
rect 9858 38196 9864 38208
rect 1443 38168 9864 38196
rect 1443 38165 1455 38168
rect 1397 38159 1455 38165
rect 9858 38156 9864 38168
rect 9916 38156 9922 38208
rect 15470 38196 15476 38208
rect 15431 38168 15476 38196
rect 15470 38156 15476 38168
rect 15528 38156 15534 38208
rect 15654 38156 15660 38208
rect 15712 38196 15718 38208
rect 17144 38196 17172 38227
rect 15712 38168 17172 38196
rect 15712 38156 15718 38168
rect 18874 38156 18880 38208
rect 18932 38196 18938 38208
rect 19429 38199 19487 38205
rect 19429 38196 19441 38199
rect 18932 38168 19441 38196
rect 18932 38156 18938 38168
rect 19429 38165 19441 38168
rect 19475 38165 19487 38199
rect 19429 38159 19487 38165
rect 23293 38199 23351 38205
rect 23293 38165 23305 38199
rect 23339 38196 23351 38199
rect 23842 38196 23848 38208
rect 23339 38168 23848 38196
rect 23339 38165 23351 38168
rect 23293 38159 23351 38165
rect 23842 38156 23848 38168
rect 23900 38156 23906 38208
rect 24118 38156 24124 38208
rect 24176 38196 24182 38208
rect 24412 38196 24440 38295
rect 25774 38292 25780 38306
rect 25832 38292 25838 38344
rect 26068 38332 26096 38508
rect 28902 38496 28908 38548
rect 28960 38536 28966 38548
rect 30374 38536 30380 38548
rect 28960 38508 30380 38536
rect 28960 38496 28966 38508
rect 30374 38496 30380 38508
rect 30432 38496 30438 38548
rect 28166 38428 28172 38480
rect 28224 38468 28230 38480
rect 29822 38468 29828 38480
rect 28224 38440 29828 38468
rect 28224 38428 28230 38440
rect 29822 38428 29828 38440
rect 29880 38428 29886 38480
rect 25976 38304 26096 38332
rect 25498 38224 25504 38276
rect 25556 38264 25562 38276
rect 25976 38264 26004 38304
rect 26602 38292 26608 38344
rect 26660 38332 26666 38344
rect 27341 38335 27399 38341
rect 27341 38332 27353 38335
rect 26660 38304 27353 38332
rect 26660 38292 26666 38304
rect 27341 38301 27353 38304
rect 27387 38301 27399 38335
rect 27341 38295 27399 38301
rect 29178 38292 29184 38344
rect 29236 38332 29242 38344
rect 29825 38335 29883 38341
rect 29825 38332 29837 38335
rect 29236 38304 29837 38332
rect 29236 38292 29242 38304
rect 29825 38301 29837 38304
rect 29871 38301 29883 38335
rect 29825 38295 29883 38301
rect 30190 38292 30196 38344
rect 30248 38332 30254 38344
rect 30374 38332 30380 38344
rect 30248 38304 30380 38332
rect 30248 38292 30254 38304
rect 30374 38292 30380 38304
rect 30432 38292 30438 38344
rect 25556 38236 26004 38264
rect 25556 38224 25562 38236
rect 26050 38224 26056 38276
rect 26108 38264 26114 38276
rect 26234 38264 26240 38276
rect 26108 38236 26240 38264
rect 26108 38224 26114 38236
rect 26234 38224 26240 38236
rect 26292 38264 26298 38276
rect 28169 38267 28227 38273
rect 28169 38264 28181 38267
rect 26292 38236 28181 38264
rect 26292 38224 26298 38236
rect 28169 38233 28181 38236
rect 28215 38233 28227 38267
rect 28169 38227 28227 38233
rect 24176 38168 24440 38196
rect 24176 38156 24182 38168
rect 26602 38156 26608 38208
rect 26660 38196 26666 38208
rect 27525 38199 27583 38205
rect 27525 38196 27537 38199
rect 26660 38168 27537 38196
rect 26660 38156 26666 38168
rect 27525 38165 27537 38168
rect 27571 38165 27583 38199
rect 28258 38196 28264 38208
rect 28219 38168 28264 38196
rect 27525 38159 27583 38165
rect 28258 38156 28264 38168
rect 28316 38156 28322 38208
rect 30009 38199 30067 38205
rect 30009 38165 30021 38199
rect 30055 38196 30067 38199
rect 30190 38196 30196 38208
rect 30055 38168 30196 38196
rect 30055 38165 30067 38168
rect 30009 38159 30067 38165
rect 30190 38156 30196 38168
rect 30248 38156 30254 38208
rect 1104 38106 30820 38128
rect 1104 38054 10880 38106
rect 10932 38054 10944 38106
rect 10996 38054 11008 38106
rect 11060 38054 11072 38106
rect 11124 38054 11136 38106
rect 11188 38054 20811 38106
rect 20863 38054 20875 38106
rect 20927 38054 20939 38106
rect 20991 38054 21003 38106
rect 21055 38054 21067 38106
rect 21119 38054 30820 38106
rect 1104 38032 30820 38054
rect 8113 37995 8171 38001
rect 8113 37961 8125 37995
rect 8159 37992 8171 37995
rect 8386 37992 8392 38004
rect 8159 37964 8392 37992
rect 8159 37961 8171 37964
rect 8113 37955 8171 37961
rect 8386 37952 8392 37964
rect 8444 37952 8450 38004
rect 9217 37995 9275 38001
rect 9217 37961 9229 37995
rect 9263 37992 9275 37995
rect 10042 37992 10048 38004
rect 9263 37964 10048 37992
rect 9263 37961 9275 37964
rect 9217 37955 9275 37961
rect 10042 37952 10048 37964
rect 10100 37952 10106 38004
rect 10965 37995 11023 38001
rect 10965 37961 10977 37995
rect 11011 37992 11023 37995
rect 11606 37992 11612 38004
rect 11011 37964 11612 37992
rect 11011 37961 11023 37964
rect 10965 37955 11023 37961
rect 11606 37952 11612 37964
rect 11664 37952 11670 38004
rect 12710 37952 12716 38004
rect 12768 37992 12774 38004
rect 12986 37992 12992 38004
rect 12768 37964 12992 37992
rect 12768 37952 12774 37964
rect 12986 37952 12992 37964
rect 13044 37952 13050 38004
rect 14182 37952 14188 38004
rect 14240 37992 14246 38004
rect 14550 37992 14556 38004
rect 14240 37964 14556 37992
rect 14240 37952 14246 37964
rect 14550 37952 14556 37964
rect 14608 37992 14614 38004
rect 15289 37995 15347 38001
rect 15289 37992 15301 37995
rect 14608 37964 15301 37992
rect 14608 37952 14614 37964
rect 15289 37961 15301 37964
rect 15335 37961 15347 37995
rect 16666 37992 16672 38004
rect 16627 37964 16672 37992
rect 15289 37955 15347 37961
rect 16666 37952 16672 37964
rect 16724 37952 16730 38004
rect 18506 37952 18512 38004
rect 18564 37992 18570 38004
rect 18693 37995 18751 38001
rect 18693 37992 18705 37995
rect 18564 37964 18705 37992
rect 18564 37952 18570 37964
rect 18693 37961 18705 37964
rect 18739 37961 18751 37995
rect 18693 37955 18751 37961
rect 22646 37952 22652 38004
rect 22704 37992 22710 38004
rect 23661 37995 23719 38001
rect 23661 37992 23673 37995
rect 22704 37964 23673 37992
rect 22704 37952 22710 37964
rect 23661 37961 23673 37964
rect 23707 37961 23719 37995
rect 25222 37992 25228 38004
rect 23661 37955 23719 37961
rect 24780 37964 25228 37992
rect 9030 37924 9036 37936
rect 8991 37896 9036 37924
rect 9030 37884 9036 37896
rect 9088 37884 9094 37936
rect 9858 37924 9864 37936
rect 9819 37896 9864 37924
rect 9858 37884 9864 37896
rect 9916 37884 9922 37936
rect 12158 37884 12164 37936
rect 12216 37924 12222 37936
rect 13998 37924 14004 37936
rect 12216 37896 13860 37924
rect 13959 37896 14004 37924
rect 12216 37884 12222 37896
rect 1394 37816 1400 37868
rect 1452 37856 1458 37868
rect 1581 37859 1639 37865
rect 1581 37856 1593 37859
rect 1452 37828 1593 37856
rect 1452 37816 1458 37828
rect 1581 37825 1593 37828
rect 1627 37825 1639 37859
rect 8294 37856 8300 37868
rect 8255 37828 8300 37856
rect 1581 37819 1639 37825
rect 8294 37816 8300 37828
rect 8352 37816 8358 37868
rect 8849 37859 8907 37865
rect 8849 37825 8861 37859
rect 8895 37856 8907 37859
rect 9582 37856 9588 37868
rect 8895 37828 9588 37856
rect 8895 37825 8907 37828
rect 8849 37819 8907 37825
rect 9582 37816 9588 37828
rect 9640 37856 9646 37868
rect 9677 37859 9735 37865
rect 9677 37856 9689 37859
rect 9640 37828 9689 37856
rect 9640 37816 9646 37828
rect 9677 37825 9689 37828
rect 9723 37825 9735 37859
rect 9677 37819 9735 37825
rect 10781 37859 10839 37865
rect 10781 37825 10793 37859
rect 10827 37856 10839 37859
rect 11422 37856 11428 37868
rect 10827 37828 11428 37856
rect 10827 37825 10839 37828
rect 10781 37819 10839 37825
rect 11422 37816 11428 37828
rect 11480 37816 11486 37868
rect 11876 37859 11934 37865
rect 11876 37825 11888 37859
rect 11922 37856 11934 37859
rect 12434 37856 12440 37868
rect 11922 37828 12440 37856
rect 11922 37825 11934 37828
rect 11876 37819 11934 37825
rect 12434 37816 12440 37828
rect 12492 37816 12498 37868
rect 11606 37788 11612 37800
rect 11567 37760 11612 37788
rect 11606 37748 11612 37760
rect 11664 37748 11670 37800
rect 13832 37788 13860 37896
rect 13998 37884 14004 37896
rect 14056 37884 14062 37936
rect 15470 37884 15476 37936
rect 15528 37924 15534 37936
rect 15528 37896 17908 37924
rect 15528 37884 15534 37896
rect 16960 37865 16988 37896
rect 16945 37859 17003 37865
rect 16945 37825 16957 37859
rect 16991 37825 17003 37859
rect 16945 37819 17003 37825
rect 17037 37859 17095 37865
rect 17037 37825 17049 37859
rect 17083 37825 17095 37859
rect 17037 37819 17095 37825
rect 17129 37859 17187 37865
rect 17129 37825 17141 37859
rect 17175 37825 17187 37859
rect 17310 37856 17316 37868
rect 17271 37828 17316 37856
rect 17129 37819 17187 37825
rect 17052 37788 17080 37819
rect 13832 37760 17080 37788
rect 13722 37680 13728 37732
rect 13780 37720 13786 37732
rect 17144 37720 17172 37819
rect 17310 37816 17316 37828
rect 17368 37816 17374 37868
rect 17773 37859 17831 37865
rect 17773 37825 17785 37859
rect 17819 37825 17831 37859
rect 17880 37856 17908 37896
rect 18230 37884 18236 37936
rect 18288 37924 18294 37936
rect 18601 37927 18659 37933
rect 18601 37924 18613 37927
rect 18288 37896 18613 37924
rect 18288 37884 18294 37896
rect 18601 37893 18613 37896
rect 18647 37893 18659 37927
rect 21726 37924 21732 37936
rect 18601 37887 18659 37893
rect 18708 37896 21732 37924
rect 18708 37856 18736 37896
rect 21726 37884 21732 37896
rect 21784 37884 21790 37936
rect 24578 37884 24584 37936
rect 24636 37924 24642 37936
rect 24673 37927 24731 37933
rect 24673 37924 24685 37927
rect 24636 37896 24685 37924
rect 24636 37884 24642 37896
rect 24673 37893 24685 37896
rect 24719 37924 24731 37927
rect 24780 37924 24808 37964
rect 25222 37952 25228 37964
rect 25280 37952 25286 38004
rect 26050 37992 26056 38004
rect 26011 37964 26056 37992
rect 26050 37952 26056 37964
rect 26108 37952 26114 38004
rect 27246 37992 27252 38004
rect 27207 37964 27252 37992
rect 27246 37952 27252 37964
rect 27304 37952 27310 38004
rect 27614 37952 27620 38004
rect 27672 37952 27678 38004
rect 28810 37952 28816 38004
rect 28868 37952 28874 38004
rect 29822 37952 29828 38004
rect 29880 37992 29886 38004
rect 29917 37995 29975 38001
rect 29917 37992 29929 37995
rect 29880 37964 29929 37992
rect 29880 37952 29886 37964
rect 29917 37961 29929 37964
rect 29963 37961 29975 37995
rect 29917 37955 29975 37961
rect 24719 37896 24808 37924
rect 24719 37893 24731 37896
rect 24673 37887 24731 37893
rect 24872 37884 24878 37936
rect 24930 37924 24936 37936
rect 25866 37924 25872 37936
rect 24930 37896 24975 37924
rect 25827 37896 25872 37924
rect 24930 37884 24936 37896
rect 25866 37884 25872 37896
rect 25924 37884 25930 37936
rect 26602 37884 26608 37936
rect 26660 37924 26666 37936
rect 27632 37924 27660 37952
rect 28166 37924 28172 37936
rect 26660 37896 27660 37924
rect 27724 37896 28172 37924
rect 26660 37884 26666 37896
rect 17880 37828 18736 37856
rect 17773 37819 17831 37825
rect 17218 37748 17224 37800
rect 17276 37788 17282 37800
rect 17788 37788 17816 37819
rect 19610 37816 19616 37868
rect 19668 37856 19674 37868
rect 19981 37859 20039 37865
rect 19981 37856 19993 37859
rect 19668 37828 19993 37856
rect 19668 37816 19674 37828
rect 19981 37825 19993 37828
rect 20027 37825 20039 37859
rect 23658 37856 23664 37868
rect 23619 37828 23664 37856
rect 19981 37819 20039 37825
rect 23658 37816 23664 37828
rect 23716 37856 23722 37868
rect 24118 37856 24124 37868
rect 23716 37828 24124 37856
rect 23716 37816 23722 37828
rect 24118 37816 24124 37828
rect 24176 37816 24182 37868
rect 24785 37859 24843 37865
rect 24785 37856 24797 37859
rect 24780 37825 24797 37856
rect 24831 37825 24843 37859
rect 25038 37856 25044 37868
rect 24999 37828 25044 37856
rect 24780 37819 24843 37825
rect 17276 37760 17816 37788
rect 17276 37748 17282 37760
rect 24486 37720 24492 37732
rect 13780 37692 17172 37720
rect 24447 37692 24492 37720
rect 13780 37680 13786 37692
rect 24486 37680 24492 37692
rect 24544 37680 24550 37732
rect 24780 37664 24808 37819
rect 25038 37816 25044 37828
rect 25096 37816 25102 37868
rect 26970 37816 26976 37868
rect 27028 37856 27034 37868
rect 27724 37865 27752 37896
rect 28166 37884 28172 37896
rect 28224 37924 28230 37936
rect 28828 37924 28856 37952
rect 28224 37896 28856 37924
rect 28224 37884 28230 37896
rect 27433 37859 27491 37865
rect 27433 37856 27445 37859
rect 27028 37828 27445 37856
rect 27028 37816 27034 37828
rect 27433 37825 27445 37828
rect 27479 37825 27491 37859
rect 27433 37819 27491 37825
rect 27617 37859 27675 37865
rect 27617 37825 27629 37859
rect 27663 37825 27675 37859
rect 27617 37819 27675 37825
rect 27709 37859 27767 37865
rect 27709 37825 27721 37859
rect 27755 37825 27767 37859
rect 28258 37856 28264 37868
rect 28219 37828 28264 37856
rect 27709 37819 27767 37825
rect 25222 37748 25228 37800
rect 25280 37788 25286 37800
rect 26145 37791 26203 37797
rect 26145 37788 26157 37791
rect 25280 37760 26157 37788
rect 25280 37748 25286 37760
rect 26145 37757 26157 37760
rect 26191 37757 26203 37791
rect 26145 37751 26203 37757
rect 26234 37748 26240 37800
rect 26292 37788 26298 37800
rect 27632 37788 27660 37819
rect 28258 37816 28264 37828
rect 28316 37816 28322 37868
rect 29454 37816 29460 37868
rect 29512 37856 29518 37868
rect 29733 37859 29791 37865
rect 29733 37856 29745 37859
rect 29512 37828 29745 37856
rect 29512 37816 29518 37828
rect 29733 37825 29745 37828
rect 29779 37825 29791 37859
rect 29733 37819 29791 37825
rect 29822 37816 29828 37868
rect 29880 37856 29886 37868
rect 30009 37859 30067 37865
rect 30009 37856 30021 37859
rect 29880 37828 30021 37856
rect 29880 37816 29886 37828
rect 30009 37825 30021 37828
rect 30055 37825 30067 37859
rect 30009 37819 30067 37825
rect 26292 37760 27660 37788
rect 28537 37791 28595 37797
rect 26292 37748 26298 37760
rect 28537 37757 28549 37791
rect 28583 37788 28595 37791
rect 29840 37788 29868 37816
rect 28583 37760 29868 37788
rect 28583 37757 28595 37760
rect 28537 37751 28595 37757
rect 1397 37655 1455 37661
rect 1397 37621 1409 37655
rect 1443 37652 1455 37655
rect 9122 37652 9128 37664
rect 1443 37624 9128 37652
rect 1443 37621 1455 37624
rect 1397 37615 1455 37621
rect 9122 37612 9128 37624
rect 9180 37612 9186 37664
rect 10045 37655 10103 37661
rect 10045 37621 10057 37655
rect 10091 37652 10103 37655
rect 12250 37652 12256 37664
rect 10091 37624 12256 37652
rect 10091 37621 10103 37624
rect 10045 37615 10103 37621
rect 12250 37612 12256 37624
rect 12308 37612 12314 37664
rect 15654 37612 15660 37664
rect 15712 37652 15718 37664
rect 16206 37652 16212 37664
rect 15712 37624 16212 37652
rect 15712 37612 15718 37624
rect 16206 37612 16212 37624
rect 16264 37612 16270 37664
rect 17957 37655 18015 37661
rect 17957 37621 17969 37655
rect 18003 37652 18015 37655
rect 18322 37652 18328 37664
rect 18003 37624 18328 37652
rect 18003 37621 18015 37624
rect 17957 37615 18015 37621
rect 18322 37612 18328 37624
rect 18380 37612 18386 37664
rect 20162 37652 20168 37664
rect 20123 37624 20168 37652
rect 20162 37612 20168 37624
rect 20220 37612 20226 37664
rect 24762 37612 24768 37664
rect 24820 37612 24826 37664
rect 25038 37612 25044 37664
rect 25096 37652 25102 37664
rect 25593 37655 25651 37661
rect 25593 37652 25605 37655
rect 25096 37624 25605 37652
rect 25096 37612 25102 37624
rect 25593 37621 25605 37624
rect 25639 37621 25651 37655
rect 25593 37615 25651 37621
rect 28350 37612 28356 37664
rect 28408 37652 28414 37664
rect 28718 37652 28724 37664
rect 28408 37624 28724 37652
rect 28408 37612 28414 37624
rect 28718 37612 28724 37624
rect 28776 37612 28782 37664
rect 28994 37612 29000 37664
rect 29052 37652 29058 37664
rect 29549 37655 29607 37661
rect 29549 37652 29561 37655
rect 29052 37624 29561 37652
rect 29052 37612 29058 37624
rect 29549 37621 29561 37624
rect 29595 37621 29607 37655
rect 29549 37615 29607 37621
rect 1104 37562 30820 37584
rect 1104 37510 5915 37562
rect 5967 37510 5979 37562
rect 6031 37510 6043 37562
rect 6095 37510 6107 37562
rect 6159 37510 6171 37562
rect 6223 37510 15846 37562
rect 15898 37510 15910 37562
rect 15962 37510 15974 37562
rect 16026 37510 16038 37562
rect 16090 37510 16102 37562
rect 16154 37510 25776 37562
rect 25828 37510 25840 37562
rect 25892 37510 25904 37562
rect 25956 37510 25968 37562
rect 26020 37510 26032 37562
rect 26084 37510 30820 37562
rect 1104 37488 30820 37510
rect 2498 37408 2504 37460
rect 2556 37448 2562 37460
rect 4341 37451 4399 37457
rect 4341 37448 4353 37451
rect 2556 37420 4353 37448
rect 2556 37408 2562 37420
rect 4341 37417 4353 37420
rect 4387 37417 4399 37451
rect 9582 37448 9588 37460
rect 9543 37420 9588 37448
rect 4341 37411 4399 37417
rect 9582 37408 9588 37420
rect 9640 37408 9646 37460
rect 12158 37448 12164 37460
rect 11716 37420 12164 37448
rect 8202 37204 8208 37256
rect 8260 37244 8266 37256
rect 11716 37253 11744 37420
rect 12158 37408 12164 37420
rect 12216 37408 12222 37460
rect 12434 37408 12440 37460
rect 12492 37448 12498 37460
rect 12492 37420 12537 37448
rect 12492 37408 12498 37420
rect 13538 37408 13544 37460
rect 13596 37448 13602 37460
rect 17218 37448 17224 37460
rect 13596 37420 17080 37448
rect 17179 37420 17224 37448
rect 13596 37408 13602 37420
rect 11790 37340 11796 37392
rect 11848 37380 11854 37392
rect 11848 37352 12020 37380
rect 11848 37340 11854 37352
rect 11992 37253 12020 37352
rect 12176 37312 12204 37408
rect 12526 37340 12532 37392
rect 12584 37380 12590 37392
rect 17052 37380 17080 37420
rect 17218 37408 17224 37420
rect 17276 37408 17282 37460
rect 21269 37451 21327 37457
rect 21269 37448 21281 37451
rect 17420 37420 21281 37448
rect 17420 37380 17448 37420
rect 21269 37417 21281 37420
rect 21315 37417 21327 37451
rect 21269 37411 21327 37417
rect 26513 37451 26571 37457
rect 26513 37417 26525 37451
rect 26559 37448 26571 37451
rect 27154 37448 27160 37460
rect 26559 37420 27160 37448
rect 26559 37417 26571 37420
rect 26513 37411 26571 37417
rect 27154 37408 27160 37420
rect 27212 37408 27218 37460
rect 27246 37408 27252 37460
rect 27304 37448 27310 37460
rect 27522 37448 27528 37460
rect 27304 37420 27528 37448
rect 27304 37408 27310 37420
rect 27522 37408 27528 37420
rect 27580 37408 27586 37460
rect 28353 37451 28411 37457
rect 28353 37417 28365 37451
rect 28399 37448 28411 37451
rect 29178 37448 29184 37460
rect 28399 37420 29184 37448
rect 28399 37417 28411 37420
rect 28353 37411 28411 37417
rect 29178 37408 29184 37420
rect 29236 37408 29242 37460
rect 29546 37408 29552 37460
rect 29604 37448 29610 37460
rect 29604 37420 30236 37448
rect 29604 37408 29610 37420
rect 12584 37352 12940 37380
rect 17052 37352 17448 37380
rect 12584 37340 12590 37352
rect 12912 37312 12940 37352
rect 17678 37340 17684 37392
rect 17736 37380 17742 37392
rect 17736 37352 18736 37380
rect 17736 37340 17742 37352
rect 13722 37312 13728 37324
rect 12176 37284 12848 37312
rect 8941 37247 8999 37253
rect 8941 37244 8953 37247
rect 8260 37216 8953 37244
rect 8260 37204 8266 37216
rect 8941 37213 8953 37216
rect 8987 37213 8999 37247
rect 8941 37207 8999 37213
rect 11609 37247 11667 37253
rect 11609 37213 11621 37247
rect 11655 37213 11667 37247
rect 11609 37207 11667 37213
rect 11701 37247 11759 37253
rect 11701 37213 11713 37247
rect 11747 37213 11759 37247
rect 11701 37207 11759 37213
rect 11793 37247 11851 37253
rect 11793 37213 11805 37247
rect 11839 37238 11851 37247
rect 11977 37247 12035 37253
rect 11839 37213 11928 37238
rect 11793 37210 11928 37213
rect 11793 37207 11851 37210
rect 4249 37179 4307 37185
rect 4249 37145 4261 37179
rect 4295 37176 4307 37179
rect 8294 37176 8300 37188
rect 4295 37148 8300 37176
rect 4295 37145 4307 37148
rect 4249 37139 4307 37145
rect 8294 37136 8300 37148
rect 8352 37136 8358 37188
rect 11624 37176 11652 37207
rect 11900 37176 11928 37210
rect 11977 37213 11989 37247
rect 12023 37213 12035 37247
rect 12526 37244 12532 37256
rect 11977 37207 12035 37213
rect 12084 37216 12532 37244
rect 12084 37176 12112 37216
rect 12526 37204 12532 37216
rect 12584 37204 12590 37256
rect 12710 37244 12716 37256
rect 12671 37216 12716 37244
rect 12710 37204 12716 37216
rect 12768 37204 12774 37256
rect 12820 37253 12848 37284
rect 12912 37284 13728 37312
rect 12912 37253 12940 37284
rect 13722 37272 13728 37284
rect 13780 37272 13786 37324
rect 18230 37312 18236 37324
rect 18191 37284 18236 37312
rect 18230 37272 18236 37284
rect 18288 37272 18294 37324
rect 18708 37321 18736 37352
rect 21910 37340 21916 37392
rect 21968 37380 21974 37392
rect 24762 37380 24768 37392
rect 21968 37352 22508 37380
rect 21968 37340 21974 37352
rect 18693 37315 18751 37321
rect 18693 37281 18705 37315
rect 18739 37281 18751 37315
rect 18693 37275 18751 37281
rect 18966 37272 18972 37324
rect 19024 37312 19030 37324
rect 21928 37312 21956 37340
rect 19024 37284 19380 37312
rect 19024 37272 19030 37284
rect 12805 37247 12863 37253
rect 12805 37213 12817 37247
rect 12851 37213 12863 37247
rect 12805 37207 12863 37213
rect 12897 37247 12955 37253
rect 12897 37213 12909 37247
rect 12943 37213 12955 37247
rect 12897 37207 12955 37213
rect 13081 37247 13139 37253
rect 13081 37213 13093 37247
rect 13127 37213 13139 37247
rect 13081 37207 13139 37213
rect 15105 37247 15163 37253
rect 15105 37213 15117 37247
rect 15151 37244 15163 37247
rect 15194 37244 15200 37256
rect 15151 37216 15200 37244
rect 15151 37213 15163 37216
rect 15105 37207 15163 37213
rect 11624 37148 11836 37176
rect 11900 37148 12112 37176
rect 11333 37111 11391 37117
rect 11333 37077 11345 37111
rect 11379 37108 11391 37111
rect 11698 37108 11704 37120
rect 11379 37080 11704 37108
rect 11379 37077 11391 37080
rect 11333 37071 11391 37077
rect 11698 37068 11704 37080
rect 11756 37068 11762 37120
rect 11808 37108 11836 37148
rect 12250 37136 12256 37188
rect 12308 37176 12314 37188
rect 13096 37176 13124 37207
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 16666 37244 16672 37256
rect 15488 37216 16672 37244
rect 12308 37148 13124 37176
rect 12308 37136 12314 37148
rect 15010 37136 15016 37188
rect 15068 37176 15074 37188
rect 15350 37179 15408 37185
rect 15350 37176 15362 37179
rect 15068 37148 15362 37176
rect 15068 37136 15074 37148
rect 15350 37145 15362 37148
rect 15396 37145 15408 37179
rect 15350 37139 15408 37145
rect 12802 37108 12808 37120
rect 11808 37080 12808 37108
rect 12802 37068 12808 37080
rect 12860 37068 12866 37120
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 15488 37108 15516 37216
rect 16666 37204 16672 37216
rect 16724 37244 16730 37256
rect 17129 37247 17187 37253
rect 17129 37244 17141 37247
rect 16724 37216 17141 37244
rect 16724 37204 16730 37216
rect 17129 37213 17141 37216
rect 17175 37213 17187 37247
rect 18414 37244 18420 37256
rect 18375 37216 18420 37244
rect 17129 37207 17187 37213
rect 18414 37204 18420 37216
rect 18472 37204 18478 37256
rect 18601 37247 18659 37253
rect 18601 37213 18613 37247
rect 18647 37241 18659 37247
rect 19242 37244 19248 37256
rect 18647 37213 18736 37241
rect 19203 37216 19248 37244
rect 18601 37207 18659 37213
rect 15562 37136 15568 37188
rect 15620 37176 15626 37188
rect 18708 37176 18736 37213
rect 19242 37204 19248 37216
rect 19300 37204 19306 37256
rect 19352 37244 19380 37284
rect 20456 37284 21956 37312
rect 19501 37247 19559 37253
rect 19501 37244 19513 37247
rect 19352 37216 19513 37244
rect 19501 37213 19513 37216
rect 19547 37213 19559 37247
rect 19501 37207 19559 37213
rect 19886 37176 19892 37188
rect 15620 37148 16620 37176
rect 18708 37148 19892 37176
rect 15620 37136 15626 37148
rect 16482 37108 16488 37120
rect 13596 37080 15516 37108
rect 16443 37080 16488 37108
rect 13596 37068 13602 37080
rect 16482 37068 16488 37080
rect 16540 37068 16546 37120
rect 16592 37108 16620 37148
rect 19886 37136 19892 37148
rect 19944 37136 19950 37188
rect 20456 37108 20484 37284
rect 21266 37244 21272 37256
rect 21227 37216 21272 37244
rect 21266 37204 21272 37216
rect 21324 37204 21330 37256
rect 21910 37244 21916 37256
rect 21871 37216 21916 37244
rect 21910 37204 21916 37216
rect 21968 37204 21974 37256
rect 22278 37204 22284 37256
rect 22336 37244 22342 37256
rect 22373 37247 22431 37253
rect 22373 37244 22385 37247
rect 22336 37216 22385 37244
rect 22336 37204 22342 37216
rect 22373 37213 22385 37216
rect 22419 37213 22431 37247
rect 22480 37244 22508 37352
rect 24688 37352 24768 37380
rect 24578 37312 24584 37324
rect 24539 37284 24584 37312
rect 24578 37272 24584 37284
rect 24636 37272 24642 37324
rect 24688 37321 24716 37352
rect 24762 37340 24768 37352
rect 24820 37340 24826 37392
rect 26970 37380 26976 37392
rect 26712 37352 26976 37380
rect 24673 37315 24731 37321
rect 24673 37281 24685 37315
rect 24719 37281 24731 37315
rect 24673 37275 24731 37281
rect 24857 37315 24915 37321
rect 24857 37281 24869 37315
rect 24903 37312 24915 37315
rect 25498 37312 25504 37324
rect 24903 37284 25504 37312
rect 24903 37281 24915 37284
rect 24857 37275 24915 37281
rect 25498 37272 25504 37284
rect 25556 37272 25562 37324
rect 26712 37253 26740 37352
rect 26970 37340 26976 37352
rect 27028 37340 27034 37392
rect 28626 37380 28632 37392
rect 27816 37352 28632 37380
rect 27816 37312 27844 37352
rect 28626 37340 28632 37352
rect 28684 37340 28690 37392
rect 29546 37312 29552 37324
rect 26804 37284 27844 37312
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 22480 37216 24777 37244
rect 22373 37207 22431 37213
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 26697 37247 26755 37253
rect 26697 37213 26709 37247
rect 26743 37213 26755 37247
rect 26697 37207 26755 37213
rect 21726 37136 21732 37188
rect 21784 37176 21790 37188
rect 26804 37176 26832 37284
rect 26973 37247 27031 37253
rect 26973 37213 26985 37247
rect 27019 37213 27031 37247
rect 27614 37244 27620 37256
rect 27575 37216 27620 37244
rect 26973 37207 27031 37213
rect 21784 37148 26832 37176
rect 26988 37176 27016 37207
rect 27614 37204 27620 37216
rect 27672 37204 27678 37256
rect 27816 37253 27844 37284
rect 27908 37284 29552 37312
rect 27908 37253 27936 37284
rect 29546 37272 29552 37284
rect 29604 37312 29610 37324
rect 29822 37312 29828 37324
rect 29604 37284 29828 37312
rect 29604 37272 29610 37284
rect 29822 37272 29828 37284
rect 29880 37312 29886 37324
rect 29880 37284 30052 37312
rect 29880 37272 29886 37284
rect 27801 37247 27859 37253
rect 27801 37213 27813 37247
rect 27847 37213 27859 37247
rect 27801 37207 27859 37213
rect 27893 37247 27951 37253
rect 27893 37213 27905 37247
rect 27939 37244 27951 37247
rect 27982 37244 27988 37256
rect 27939 37216 27988 37244
rect 27939 37213 27951 37216
rect 27893 37207 27951 37213
rect 27982 37204 27988 37216
rect 28040 37204 28046 37256
rect 28626 37244 28632 37256
rect 28587 37216 28632 37244
rect 28626 37204 28632 37216
rect 28684 37204 28690 37256
rect 28721 37247 28779 37253
rect 28721 37213 28733 37247
rect 28767 37213 28779 37247
rect 28721 37207 28779 37213
rect 28813 37247 28871 37253
rect 28813 37213 28825 37247
rect 28859 37213 28871 37247
rect 28813 37207 28871 37213
rect 28997 37247 29055 37253
rect 28997 37213 29009 37247
rect 29043 37244 29055 37247
rect 29086 37244 29092 37256
rect 29043 37216 29092 37244
rect 29043 37213 29055 37216
rect 28997 37207 29055 37213
rect 28166 37176 28172 37188
rect 26988 37148 28172 37176
rect 21784 37136 21790 37148
rect 28166 37136 28172 37148
rect 28224 37136 28230 37188
rect 16592 37080 20484 37108
rect 20625 37111 20683 37117
rect 20625 37077 20637 37111
rect 20671 37108 20683 37111
rect 21818 37108 21824 37120
rect 20671 37080 21824 37108
rect 20671 37077 20683 37080
rect 20625 37071 20683 37077
rect 21818 37068 21824 37080
rect 21876 37068 21882 37120
rect 22002 37068 22008 37120
rect 22060 37108 22066 37120
rect 22557 37111 22615 37117
rect 22557 37108 22569 37111
rect 22060 37080 22569 37108
rect 22060 37068 22066 37080
rect 22557 37077 22569 37080
rect 22603 37077 22615 37111
rect 22557 37071 22615 37077
rect 24397 37111 24455 37117
rect 24397 37077 24409 37111
rect 24443 37108 24455 37111
rect 24578 37108 24584 37120
rect 24443 37080 24584 37108
rect 24443 37077 24455 37080
rect 24397 37071 24455 37077
rect 24578 37068 24584 37080
rect 24636 37068 24642 37120
rect 26050 37068 26056 37120
rect 26108 37108 26114 37120
rect 26881 37111 26939 37117
rect 26881 37108 26893 37111
rect 26108 37080 26893 37108
rect 26108 37068 26114 37080
rect 26881 37077 26893 37080
rect 26927 37077 26939 37111
rect 26881 37071 26939 37077
rect 27433 37111 27491 37117
rect 27433 37077 27445 37111
rect 27479 37108 27491 37111
rect 27522 37108 27528 37120
rect 27479 37080 27528 37108
rect 27479 37077 27491 37080
rect 27433 37071 27491 37077
rect 27522 37068 27528 37080
rect 27580 37068 27586 37120
rect 28258 37068 28264 37120
rect 28316 37108 28322 37120
rect 28736 37108 28764 37207
rect 28316 37080 28764 37108
rect 28828 37108 28856 37207
rect 29086 37204 29092 37216
rect 29144 37204 29150 37256
rect 29454 37204 29460 37256
rect 29512 37244 29518 37256
rect 30024 37253 30052 37284
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 29512 37216 29745 37244
rect 29512 37204 29518 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 30009 37247 30067 37253
rect 30009 37213 30021 37247
rect 30055 37213 30067 37247
rect 30009 37207 30067 37213
rect 29549 37179 29607 37185
rect 29549 37145 29561 37179
rect 29595 37176 29607 37179
rect 30098 37176 30104 37188
rect 29595 37148 30104 37176
rect 29595 37145 29607 37148
rect 29549 37139 29607 37145
rect 30098 37136 30104 37148
rect 30156 37136 30162 37188
rect 29454 37108 29460 37120
rect 28828 37080 29460 37108
rect 28316 37068 28322 37080
rect 29454 37068 29460 37080
rect 29512 37068 29518 37120
rect 29917 37111 29975 37117
rect 29917 37077 29929 37111
rect 29963 37108 29975 37111
rect 30208 37108 30236 37420
rect 29963 37080 30236 37108
rect 29963 37077 29975 37080
rect 29917 37071 29975 37077
rect 1104 37018 30820 37040
rect 1104 36966 10880 37018
rect 10932 36966 10944 37018
rect 10996 36966 11008 37018
rect 11060 36966 11072 37018
rect 11124 36966 11136 37018
rect 11188 36966 20811 37018
rect 20863 36966 20875 37018
rect 20927 36966 20939 37018
rect 20991 36966 21003 37018
rect 21055 36966 21067 37018
rect 21119 36966 30820 37018
rect 1104 36944 30820 36966
rect 1397 36907 1455 36913
rect 1397 36873 1409 36907
rect 1443 36904 1455 36907
rect 9309 36907 9367 36913
rect 1443 36876 2774 36904
rect 1443 36873 1455 36876
rect 1397 36867 1455 36873
rect 2746 36836 2774 36876
rect 9309 36873 9321 36907
rect 9355 36904 9367 36907
rect 13446 36904 13452 36916
rect 9355 36876 13452 36904
rect 9355 36873 9367 36876
rect 9309 36867 9367 36873
rect 13446 36864 13452 36876
rect 13504 36864 13510 36916
rect 15010 36904 15016 36916
rect 14971 36876 15016 36904
rect 15010 36864 15016 36876
rect 15068 36864 15074 36916
rect 16482 36904 16488 36916
rect 15304 36876 16488 36904
rect 8297 36839 8355 36845
rect 8297 36836 8309 36839
rect 2746 36808 8309 36836
rect 8297 36805 8309 36808
rect 8343 36805 8355 36839
rect 9122 36836 9128 36848
rect 9083 36808 9128 36836
rect 8297 36799 8355 36805
rect 9122 36796 9128 36808
rect 9180 36796 9186 36848
rect 1578 36768 1584 36780
rect 1539 36740 1584 36768
rect 1578 36728 1584 36740
rect 1636 36728 1642 36780
rect 8113 36771 8171 36777
rect 8113 36737 8125 36771
rect 8159 36768 8171 36771
rect 8846 36768 8852 36780
rect 8159 36740 8852 36768
rect 8159 36737 8171 36740
rect 8113 36731 8171 36737
rect 8846 36728 8852 36740
rect 8904 36768 8910 36780
rect 8941 36771 8999 36777
rect 8941 36768 8953 36771
rect 8904 36740 8953 36768
rect 8904 36728 8910 36740
rect 8941 36737 8953 36740
rect 8987 36768 8999 36771
rect 9582 36768 9588 36780
rect 8987 36740 9588 36768
rect 8987 36737 8999 36740
rect 8941 36731 8999 36737
rect 9582 36728 9588 36740
rect 9640 36728 9646 36780
rect 13449 36771 13507 36777
rect 13449 36737 13461 36771
rect 13495 36768 13507 36771
rect 13538 36768 13544 36780
rect 13495 36740 13544 36768
rect 13495 36737 13507 36740
rect 13449 36731 13507 36737
rect 13538 36728 13544 36740
rect 13596 36728 13602 36780
rect 13722 36768 13728 36780
rect 13683 36740 13728 36768
rect 13722 36728 13728 36740
rect 13780 36728 13786 36780
rect 15304 36777 15332 36876
rect 16482 36864 16488 36876
rect 16540 36904 16546 36916
rect 23014 36904 23020 36916
rect 16540 36876 23020 36904
rect 16540 36864 16546 36876
rect 23014 36864 23020 36876
rect 23072 36864 23078 36916
rect 26329 36907 26387 36913
rect 26329 36873 26341 36907
rect 26375 36904 26387 36907
rect 26418 36904 26424 36916
rect 26375 36876 26424 36904
rect 26375 36873 26387 36876
rect 26329 36867 26387 36873
rect 26418 36864 26424 36876
rect 26476 36864 26482 36916
rect 28258 36864 28264 36916
rect 28316 36904 28322 36916
rect 28316 36876 28764 36904
rect 28316 36864 28322 36876
rect 15930 36836 15936 36848
rect 15396 36808 15936 36836
rect 15396 36777 15424 36808
rect 15930 36796 15936 36808
rect 15988 36796 15994 36848
rect 16574 36796 16580 36848
rect 16632 36836 16638 36848
rect 22922 36836 22928 36848
rect 16632 36808 22928 36836
rect 16632 36796 16638 36808
rect 22922 36796 22928 36808
rect 22980 36796 22986 36848
rect 27801 36839 27859 36845
rect 27801 36836 27813 36839
rect 24596 36808 27813 36836
rect 15289 36771 15347 36777
rect 15289 36737 15301 36771
rect 15335 36737 15347 36771
rect 15289 36731 15347 36737
rect 15381 36771 15439 36777
rect 15381 36737 15393 36771
rect 15427 36737 15439 36771
rect 15381 36731 15439 36737
rect 15470 36728 15476 36780
rect 15528 36768 15534 36780
rect 15657 36771 15715 36777
rect 15528 36740 15570 36768
rect 15528 36728 15534 36740
rect 15657 36737 15669 36771
rect 15703 36768 15715 36771
rect 15838 36768 15844 36780
rect 15703 36740 15844 36768
rect 15703 36737 15715 36740
rect 15657 36731 15715 36737
rect 15838 36728 15844 36740
rect 15896 36728 15902 36780
rect 17218 36728 17224 36780
rect 17276 36768 17282 36780
rect 17865 36771 17923 36777
rect 17865 36768 17877 36771
rect 17276 36740 17877 36768
rect 17276 36728 17282 36740
rect 17865 36737 17877 36740
rect 17911 36737 17923 36771
rect 18966 36768 18972 36780
rect 18927 36740 18972 36768
rect 17865 36731 17923 36737
rect 18966 36728 18972 36740
rect 19024 36728 19030 36780
rect 21174 36728 21180 36780
rect 21232 36768 21238 36780
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21232 36740 21833 36768
rect 21232 36728 21238 36740
rect 21821 36737 21833 36740
rect 21867 36768 21879 36771
rect 22002 36768 22008 36780
rect 21867 36740 22008 36768
rect 21867 36737 21879 36740
rect 21821 36731 21879 36737
rect 22002 36728 22008 36740
rect 22060 36728 22066 36780
rect 22094 36728 22100 36780
rect 22152 36768 22158 36780
rect 22152 36740 22197 36768
rect 22152 36728 22158 36740
rect 16298 36660 16304 36712
rect 16356 36700 16362 36712
rect 21726 36700 21732 36712
rect 16356 36672 21732 36700
rect 16356 36660 16362 36672
rect 21726 36660 21732 36672
rect 21784 36660 21790 36712
rect 21910 36660 21916 36712
rect 21968 36700 21974 36712
rect 22281 36703 22339 36709
rect 22281 36700 22293 36703
rect 21968 36672 22293 36700
rect 21968 36660 21974 36672
rect 22281 36669 22293 36672
rect 22327 36669 22339 36703
rect 22281 36663 22339 36669
rect 22465 36703 22523 36709
rect 22465 36669 22477 36703
rect 22511 36700 22523 36703
rect 22646 36700 22652 36712
rect 22511 36672 22652 36700
rect 22511 36669 22523 36672
rect 22465 36663 22523 36669
rect 22646 36660 22652 36672
rect 22704 36660 22710 36712
rect 8481 36635 8539 36641
rect 8481 36601 8493 36635
rect 8527 36632 8539 36635
rect 17310 36632 17316 36644
rect 8527 36604 17316 36632
rect 8527 36601 8539 36604
rect 8481 36595 8539 36601
rect 17310 36592 17316 36604
rect 17368 36592 17374 36644
rect 18049 36635 18107 36641
rect 18049 36601 18061 36635
rect 18095 36632 18107 36635
rect 18414 36632 18420 36644
rect 18095 36604 18420 36632
rect 18095 36601 18107 36604
rect 18049 36595 18107 36601
rect 18414 36592 18420 36604
rect 18472 36632 18478 36644
rect 19886 36632 19892 36644
rect 18472 36604 19892 36632
rect 18472 36592 18478 36604
rect 19886 36592 19892 36604
rect 19944 36592 19950 36644
rect 24596 36632 24624 36808
rect 26436 36780 26464 36808
rect 27801 36805 27813 36808
rect 27847 36805 27859 36839
rect 27801 36799 27859 36805
rect 25130 36728 25136 36780
rect 25188 36768 25194 36780
rect 26053 36771 26111 36777
rect 26053 36768 26065 36771
rect 25188 36740 26065 36768
rect 25188 36728 25194 36740
rect 26053 36737 26065 36740
rect 26099 36737 26111 36771
rect 26053 36731 26111 36737
rect 26418 36728 26424 36780
rect 26476 36728 26482 36780
rect 27614 36768 27620 36780
rect 27527 36740 27620 36768
rect 27614 36728 27620 36740
rect 27672 36728 27678 36780
rect 27893 36771 27951 36777
rect 27893 36737 27905 36771
rect 27939 36768 27951 36771
rect 27982 36768 27988 36780
rect 27939 36740 27988 36768
rect 27939 36737 27951 36740
rect 27893 36731 27951 36737
rect 27982 36728 27988 36740
rect 28040 36728 28046 36780
rect 28626 36768 28632 36780
rect 28539 36740 28632 36768
rect 28626 36728 28632 36740
rect 28684 36728 28690 36780
rect 28736 36777 28764 36876
rect 29178 36836 29184 36848
rect 28828 36808 29184 36836
rect 28828 36777 28856 36808
rect 29178 36796 29184 36808
rect 29236 36796 29242 36848
rect 28721 36771 28779 36777
rect 28721 36737 28733 36771
rect 28767 36737 28779 36771
rect 28721 36731 28779 36737
rect 28813 36771 28871 36777
rect 28813 36737 28825 36771
rect 28859 36737 28871 36771
rect 28994 36768 29000 36780
rect 28955 36740 29000 36768
rect 28813 36731 28871 36737
rect 28994 36728 29000 36740
rect 29052 36728 29058 36780
rect 29086 36728 29092 36780
rect 29144 36768 29150 36780
rect 29687 36771 29745 36777
rect 29687 36768 29699 36771
rect 29144 36740 29699 36768
rect 29144 36728 29150 36740
rect 29687 36737 29699 36740
rect 29733 36737 29745 36771
rect 29822 36768 29828 36780
rect 29783 36740 29828 36768
rect 29687 36731 29745 36737
rect 29822 36728 29828 36740
rect 29880 36728 29886 36780
rect 29917 36771 29975 36777
rect 29917 36737 29929 36771
rect 29963 36737 29975 36771
rect 30098 36768 30104 36780
rect 30059 36740 30104 36768
rect 29917 36731 29975 36737
rect 24762 36660 24768 36712
rect 24820 36700 24826 36712
rect 25685 36703 25743 36709
rect 25685 36700 25697 36703
rect 24820 36672 25697 36700
rect 24820 36660 24826 36672
rect 25685 36669 25697 36672
rect 25731 36669 25743 36703
rect 25685 36663 25743 36669
rect 25774 36660 25780 36712
rect 25832 36700 25838 36712
rect 25961 36703 26019 36709
rect 25961 36700 25973 36703
rect 25832 36672 25973 36700
rect 25832 36660 25838 36672
rect 25961 36669 25973 36672
rect 26007 36669 26019 36703
rect 26142 36700 26148 36712
rect 26103 36672 26148 36700
rect 25961 36663 26019 36669
rect 26142 36660 26148 36672
rect 26200 36660 26206 36712
rect 27632 36700 27660 36728
rect 28350 36700 28356 36712
rect 27632 36672 28356 36700
rect 28350 36660 28356 36672
rect 28408 36660 28414 36712
rect 28644 36700 28672 36728
rect 29104 36700 29132 36728
rect 28644 36672 29132 36700
rect 22487 36604 24624 36632
rect 14918 36524 14924 36576
rect 14976 36564 14982 36576
rect 16574 36564 16580 36576
rect 14976 36536 16580 36564
rect 14976 36524 14982 36536
rect 16574 36524 16580 36536
rect 16632 36524 16638 36576
rect 19334 36524 19340 36576
rect 19392 36564 19398 36576
rect 19794 36564 19800 36576
rect 19392 36536 19800 36564
rect 19392 36524 19398 36536
rect 19794 36524 19800 36536
rect 19852 36524 19858 36576
rect 20070 36524 20076 36576
rect 20128 36564 20134 36576
rect 20257 36567 20315 36573
rect 20257 36564 20269 36567
rect 20128 36536 20269 36564
rect 20128 36524 20134 36536
rect 20257 36533 20269 36536
rect 20303 36533 20315 36567
rect 20257 36527 20315 36533
rect 21818 36524 21824 36576
rect 21876 36564 21882 36576
rect 22487 36564 22515 36604
rect 26050 36592 26056 36644
rect 26108 36632 26114 36644
rect 26878 36632 26884 36644
rect 26108 36604 26884 36632
rect 26108 36592 26114 36604
rect 26878 36592 26884 36604
rect 26936 36592 26942 36644
rect 27433 36635 27491 36641
rect 27433 36601 27445 36635
rect 27479 36632 27491 36635
rect 28994 36632 29000 36644
rect 27479 36604 29000 36632
rect 27479 36601 27491 36604
rect 27433 36595 27491 36601
rect 28994 36592 29000 36604
rect 29052 36592 29058 36644
rect 29932 36632 29960 36731
rect 30098 36728 30104 36740
rect 30156 36728 30162 36780
rect 30098 36632 30104 36644
rect 29932 36604 30104 36632
rect 30098 36592 30104 36604
rect 30156 36592 30162 36644
rect 31294 36592 31300 36644
rect 31352 36632 31358 36644
rect 31352 36604 31524 36632
rect 31352 36592 31358 36604
rect 21876 36536 22515 36564
rect 21876 36524 21882 36536
rect 22554 36524 22560 36576
rect 22612 36564 22618 36576
rect 23382 36564 23388 36576
rect 22612 36536 23388 36564
rect 22612 36524 22618 36536
rect 23382 36524 23388 36536
rect 23440 36524 23446 36576
rect 25222 36524 25228 36576
rect 25280 36564 25286 36576
rect 25590 36564 25596 36576
rect 25280 36536 25596 36564
rect 25280 36524 25286 36536
rect 25590 36524 25596 36536
rect 25648 36524 25654 36576
rect 27614 36524 27620 36576
rect 27672 36564 27678 36576
rect 28353 36567 28411 36573
rect 28353 36564 28365 36567
rect 27672 36536 28365 36564
rect 27672 36524 27678 36536
rect 28353 36533 28365 36536
rect 28399 36533 28411 36567
rect 28353 36527 28411 36533
rect 28718 36524 28724 36576
rect 28776 36564 28782 36576
rect 29457 36567 29515 36573
rect 29457 36564 29469 36567
rect 28776 36536 29469 36564
rect 28776 36524 28782 36536
rect 29457 36533 29469 36536
rect 29503 36533 29515 36567
rect 29457 36527 29515 36533
rect 1104 36474 30820 36496
rect 1104 36422 5915 36474
rect 5967 36422 5979 36474
rect 6031 36422 6043 36474
rect 6095 36422 6107 36474
rect 6159 36422 6171 36474
rect 6223 36422 15846 36474
rect 15898 36422 15910 36474
rect 15962 36422 15974 36474
rect 16026 36422 16038 36474
rect 16090 36422 16102 36474
rect 16154 36422 25776 36474
rect 25828 36422 25840 36474
rect 25892 36422 25904 36474
rect 25956 36422 25968 36474
rect 26020 36422 26032 36474
rect 26084 36422 30820 36474
rect 1104 36400 30820 36422
rect 8202 36360 8208 36372
rect 8163 36332 8208 36360
rect 8202 36320 8208 36332
rect 8260 36320 8266 36372
rect 11057 36363 11115 36369
rect 11057 36329 11069 36363
rect 11103 36360 11115 36363
rect 11330 36360 11336 36372
rect 11103 36332 11336 36360
rect 11103 36329 11115 36332
rect 11057 36323 11115 36329
rect 11330 36320 11336 36332
rect 11388 36360 11394 36372
rect 15194 36360 15200 36372
rect 11388 36332 12434 36360
rect 15155 36332 15200 36360
rect 11388 36320 11394 36332
rect 1397 36295 1455 36301
rect 1397 36261 1409 36295
rect 1443 36292 1455 36295
rect 9030 36292 9036 36304
rect 1443 36264 9036 36292
rect 1443 36261 1455 36264
rect 1397 36255 1455 36261
rect 9030 36252 9036 36264
rect 9088 36252 9094 36304
rect 9674 36252 9680 36304
rect 9732 36252 9738 36304
rect 9692 36224 9720 36252
rect 12406 36224 12434 36332
rect 15194 36320 15200 36332
rect 15252 36320 15258 36372
rect 15746 36320 15752 36372
rect 15804 36360 15810 36372
rect 18233 36363 18291 36369
rect 18233 36360 18245 36363
rect 15804 36332 18245 36360
rect 15804 36320 15810 36332
rect 18233 36329 18245 36332
rect 18279 36329 18291 36363
rect 18233 36323 18291 36329
rect 19242 36320 19248 36372
rect 19300 36360 19306 36372
rect 19429 36363 19487 36369
rect 19429 36360 19441 36363
rect 19300 36332 19441 36360
rect 19300 36320 19306 36332
rect 19429 36329 19441 36332
rect 19475 36329 19487 36363
rect 25133 36363 25191 36369
rect 19429 36323 19487 36329
rect 19536 36332 20944 36360
rect 19536 36224 19564 36332
rect 20809 36295 20867 36301
rect 20809 36261 20821 36295
rect 20855 36261 20867 36295
rect 20916 36292 20944 36332
rect 25133 36329 25145 36363
rect 25179 36360 25191 36363
rect 26878 36360 26884 36372
rect 25179 36332 26884 36360
rect 25179 36329 25191 36332
rect 25133 36323 25191 36329
rect 25976 36304 26004 36332
rect 26878 36320 26884 36332
rect 26936 36320 26942 36372
rect 20916 36264 23612 36292
rect 20809 36255 20867 36261
rect 9692 36196 9812 36224
rect 12406 36196 19564 36224
rect 19981 36227 20039 36233
rect 1578 36156 1584 36168
rect 1539 36128 1584 36156
rect 1578 36116 1584 36128
rect 1636 36116 1642 36168
rect 8294 36116 8300 36168
rect 8352 36156 8358 36168
rect 8389 36159 8447 36165
rect 8389 36156 8401 36159
rect 8352 36128 8401 36156
rect 8352 36116 8358 36128
rect 8389 36125 8401 36128
rect 8435 36125 8447 36159
rect 9674 36156 9680 36168
rect 9635 36128 9680 36156
rect 8389 36119 8447 36125
rect 8404 36088 8432 36119
rect 9674 36116 9680 36128
rect 9732 36116 9738 36168
rect 9784 36156 9812 36196
rect 19981 36193 19993 36227
rect 20027 36224 20039 36227
rect 20346 36224 20352 36236
rect 20027 36196 20352 36224
rect 20027 36193 20039 36196
rect 19981 36187 20039 36193
rect 20346 36184 20352 36196
rect 20404 36224 20410 36236
rect 20622 36224 20628 36236
rect 20404 36196 20628 36224
rect 20404 36184 20410 36196
rect 20622 36184 20628 36196
rect 20680 36184 20686 36236
rect 9933 36159 9991 36165
rect 9933 36156 9945 36159
rect 9784 36128 9945 36156
rect 9933 36125 9945 36128
rect 9979 36125 9991 36159
rect 15010 36156 15016 36168
rect 14971 36128 15016 36156
rect 9933 36119 9991 36125
rect 15010 36116 15016 36128
rect 15068 36116 15074 36168
rect 16850 36116 16856 36168
rect 16908 36156 16914 36168
rect 16945 36159 17003 36165
rect 16945 36156 16957 36159
rect 16908 36128 16957 36156
rect 16908 36116 16914 36128
rect 16945 36125 16957 36128
rect 16991 36125 17003 36159
rect 19242 36156 19248 36168
rect 19203 36128 19248 36156
rect 16945 36119 17003 36125
rect 19242 36116 19248 36128
rect 19300 36116 19306 36168
rect 20165 36159 20223 36165
rect 20165 36125 20177 36159
rect 20211 36156 20223 36159
rect 20824 36156 20852 36255
rect 21450 36224 21456 36236
rect 21411 36196 21456 36224
rect 21450 36184 21456 36196
rect 21508 36184 21514 36236
rect 21174 36156 21180 36168
rect 20211 36128 20852 36156
rect 21135 36128 21180 36156
rect 20211 36125 20223 36128
rect 20165 36119 20223 36125
rect 21174 36116 21180 36128
rect 21232 36116 21238 36168
rect 22005 36159 22063 36165
rect 22005 36125 22017 36159
rect 22051 36156 22063 36159
rect 22094 36156 22100 36168
rect 22051 36128 22100 36156
rect 22051 36125 22063 36128
rect 22005 36119 22063 36125
rect 22094 36116 22100 36128
rect 22152 36156 22158 36168
rect 22833 36159 22891 36165
rect 22833 36156 22845 36159
rect 22152 36128 22845 36156
rect 22152 36116 22158 36128
rect 22833 36125 22845 36128
rect 22879 36125 22891 36159
rect 23584 36156 23612 36264
rect 23658 36252 23664 36304
rect 23716 36292 23722 36304
rect 24762 36292 24768 36304
rect 23716 36264 24768 36292
rect 23716 36252 23722 36264
rect 24762 36252 24768 36264
rect 24820 36292 24826 36304
rect 25685 36295 25743 36301
rect 25685 36292 25697 36295
rect 24820 36264 25697 36292
rect 24820 36252 24826 36264
rect 25685 36261 25697 36264
rect 25731 36261 25743 36295
rect 25685 36255 25743 36261
rect 25958 36252 25964 36304
rect 26016 36252 26022 36304
rect 26510 36252 26516 36304
rect 26568 36292 26574 36304
rect 29914 36292 29920 36304
rect 26568 36264 29920 36292
rect 26568 36252 26574 36264
rect 29914 36252 29920 36264
rect 29972 36252 29978 36304
rect 30558 36252 30564 36304
rect 30616 36292 30622 36304
rect 31386 36292 31392 36304
rect 30616 36264 31392 36292
rect 30616 36252 30622 36264
rect 31386 36252 31392 36264
rect 31444 36252 31450 36304
rect 24026 36184 24032 36236
rect 24084 36224 24090 36236
rect 26237 36227 26295 36233
rect 26237 36224 26249 36227
rect 24084 36196 26249 36224
rect 24084 36184 24090 36196
rect 26237 36193 26249 36196
rect 26283 36193 26295 36227
rect 28077 36227 28135 36233
rect 28077 36224 28089 36227
rect 26237 36187 26295 36193
rect 27448 36196 28089 36224
rect 27448 36168 27476 36196
rect 28077 36193 28089 36196
rect 28123 36224 28135 36227
rect 28166 36224 28172 36236
rect 28123 36196 28172 36224
rect 28123 36193 28135 36196
rect 28077 36187 28135 36193
rect 28166 36184 28172 36196
rect 28224 36184 28230 36236
rect 29362 36184 29368 36236
rect 29420 36184 29426 36236
rect 29546 36184 29552 36236
rect 29604 36224 29610 36236
rect 29604 36196 30052 36224
rect 29604 36184 29610 36196
rect 24762 36156 24768 36168
rect 23584 36128 24768 36156
rect 22833 36119 22891 36125
rect 24762 36116 24768 36128
rect 24820 36116 24826 36168
rect 24946 36156 24952 36168
rect 24907 36128 24952 36156
rect 24946 36116 24952 36128
rect 25004 36116 25010 36168
rect 25130 36116 25136 36168
rect 25188 36156 25194 36168
rect 25774 36156 25780 36168
rect 25188 36128 25780 36156
rect 25188 36116 25194 36128
rect 25774 36116 25780 36128
rect 25832 36156 25838 36168
rect 25961 36159 26019 36165
rect 25961 36156 25973 36159
rect 25832 36128 25973 36156
rect 25832 36116 25838 36128
rect 25961 36125 25973 36128
rect 26007 36125 26019 36159
rect 25961 36119 26019 36125
rect 26878 36116 26884 36168
rect 26936 36156 26942 36168
rect 27341 36159 27399 36165
rect 27341 36156 27353 36159
rect 26936 36128 27353 36156
rect 26936 36116 26942 36128
rect 27341 36125 27353 36128
rect 27387 36156 27399 36159
rect 27430 36156 27436 36168
rect 27387 36128 27436 36156
rect 27387 36125 27399 36128
rect 27341 36119 27399 36125
rect 27430 36116 27436 36128
rect 27488 36116 27494 36168
rect 27617 36159 27675 36165
rect 27617 36125 27629 36159
rect 27663 36125 27675 36159
rect 28350 36156 28356 36168
rect 28263 36128 28356 36156
rect 27617 36119 27675 36125
rect 10042 36088 10048 36100
rect 8404 36060 10048 36088
rect 10042 36048 10048 36060
rect 10100 36048 10106 36100
rect 11974 36048 11980 36100
rect 12032 36088 12038 36100
rect 21818 36088 21824 36100
rect 12032 36060 21824 36088
rect 12032 36048 12038 36060
rect 21818 36048 21824 36060
rect 21876 36048 21882 36100
rect 22189 36091 22247 36097
rect 22189 36057 22201 36091
rect 22235 36088 22247 36091
rect 22278 36088 22284 36100
rect 22235 36060 22284 36088
rect 22235 36057 22247 36060
rect 22189 36051 22247 36057
rect 22278 36048 22284 36060
rect 22336 36048 22342 36100
rect 22373 36091 22431 36097
rect 22373 36057 22385 36091
rect 22419 36088 22431 36091
rect 22554 36088 22560 36100
rect 22419 36060 22560 36088
rect 22419 36057 22431 36060
rect 22373 36051 22431 36057
rect 22554 36048 22560 36060
rect 22612 36048 22618 36100
rect 22922 36048 22928 36100
rect 22980 36088 22986 36100
rect 25866 36088 25872 36100
rect 22980 36060 24900 36088
rect 25827 36060 25872 36088
rect 22980 36048 22986 36060
rect 20346 36020 20352 36032
rect 20307 35992 20352 36020
rect 20346 35980 20352 35992
rect 20404 35980 20410 36032
rect 21269 36023 21327 36029
rect 21269 35989 21281 36023
rect 21315 36020 21327 36023
rect 21910 36020 21916 36032
rect 21315 35992 21916 36020
rect 21315 35989 21327 35992
rect 21269 35983 21327 35989
rect 21910 35980 21916 35992
rect 21968 36020 21974 36032
rect 23017 36023 23075 36029
rect 23017 36020 23029 36023
rect 21968 35992 23029 36020
rect 21968 35980 21974 35992
rect 23017 35989 23029 35992
rect 23063 35989 23075 36023
rect 24872 36020 24900 36060
rect 25866 36048 25872 36060
rect 25924 36048 25930 36100
rect 26234 36088 26240 36100
rect 25976 36060 26240 36088
rect 25976 36020 26004 36060
rect 26234 36048 26240 36060
rect 26292 36088 26298 36100
rect 27525 36091 27583 36097
rect 27525 36088 27537 36091
rect 26292 36060 27537 36088
rect 26292 36048 26298 36060
rect 27525 36057 27537 36060
rect 27571 36057 27583 36091
rect 27632 36088 27660 36119
rect 28350 36116 28356 36128
rect 28408 36156 28414 36168
rect 29380 36156 29408 36184
rect 29733 36159 29791 36165
rect 29733 36156 29745 36159
rect 28408 36128 29745 36156
rect 28408 36116 28414 36128
rect 29733 36125 29745 36128
rect 29779 36125 29791 36159
rect 29914 36156 29920 36168
rect 29875 36128 29920 36156
rect 29733 36119 29791 36125
rect 29914 36116 29920 36128
rect 29972 36116 29978 36168
rect 30024 36165 30052 36196
rect 30009 36159 30067 36165
rect 30009 36125 30021 36159
rect 30055 36125 30067 36159
rect 30009 36119 30067 36125
rect 28258 36088 28264 36100
rect 27632 36060 28264 36088
rect 27525 36051 27583 36057
rect 28258 36048 28264 36060
rect 28316 36048 28322 36100
rect 24872 35992 26004 36020
rect 23017 35983 23075 35989
rect 26050 35980 26056 36032
rect 26108 36020 26114 36032
rect 27157 36023 27215 36029
rect 26108 35992 26153 36020
rect 26108 35980 26114 35992
rect 27157 35989 27169 36023
rect 27203 36020 27215 36023
rect 27430 36020 27436 36032
rect 27203 35992 27436 36020
rect 27203 35989 27215 35992
rect 27157 35983 27215 35989
rect 27430 35980 27436 35992
rect 27488 35980 27494 36032
rect 28350 35980 28356 36032
rect 28408 36020 28414 36032
rect 28626 36020 28632 36032
rect 28408 35992 28632 36020
rect 28408 35980 28414 35992
rect 28626 35980 28632 35992
rect 28684 35980 28690 36032
rect 29178 35980 29184 36032
rect 29236 36020 29242 36032
rect 29362 36020 29368 36032
rect 29236 35992 29368 36020
rect 29236 35980 29242 35992
rect 29362 35980 29368 35992
rect 29420 35980 29426 36032
rect 29546 36020 29552 36032
rect 29507 35992 29552 36020
rect 29546 35980 29552 35992
rect 29604 35980 29610 36032
rect 1104 35930 30820 35952
rect 1104 35878 10880 35930
rect 10932 35878 10944 35930
rect 10996 35878 11008 35930
rect 11060 35878 11072 35930
rect 11124 35878 11136 35930
rect 11188 35878 20811 35930
rect 20863 35878 20875 35930
rect 20927 35878 20939 35930
rect 20991 35878 21003 35930
rect 21055 35878 21067 35930
rect 21119 35878 30820 35930
rect 31496 35884 31524 36604
rect 1104 35856 30820 35878
rect 30852 35856 31524 35884
rect 30852 35828 30880 35856
rect 20530 35776 20536 35828
rect 20588 35816 20594 35828
rect 21177 35819 21235 35825
rect 21177 35816 21189 35819
rect 20588 35788 21189 35816
rect 20588 35776 20594 35788
rect 21177 35785 21189 35788
rect 21223 35785 21235 35819
rect 21177 35779 21235 35785
rect 23658 35776 23664 35828
rect 23716 35816 23722 35828
rect 23753 35819 23811 35825
rect 23753 35816 23765 35819
rect 23716 35788 23765 35816
rect 23716 35776 23722 35788
rect 23753 35785 23765 35788
rect 23799 35785 23811 35819
rect 23753 35779 23811 35785
rect 24026 35776 24032 35828
rect 24084 35816 24090 35828
rect 24762 35816 24768 35828
rect 24084 35788 24768 35816
rect 24084 35776 24090 35788
rect 24762 35776 24768 35788
rect 24820 35816 24826 35828
rect 25958 35816 25964 35828
rect 24820 35788 25964 35816
rect 24820 35776 24826 35788
rect 25958 35776 25964 35788
rect 26016 35776 26022 35828
rect 27709 35819 27767 35825
rect 27709 35785 27721 35819
rect 27755 35816 27767 35819
rect 27982 35816 27988 35828
rect 27755 35788 27988 35816
rect 27755 35785 27767 35788
rect 27709 35779 27767 35785
rect 27982 35776 27988 35788
rect 28040 35776 28046 35828
rect 30282 35776 30288 35828
rect 30340 35776 30346 35828
rect 30834 35776 30840 35828
rect 30892 35776 30898 35828
rect 8846 35748 8852 35760
rect 8807 35720 8852 35748
rect 8846 35708 8852 35720
rect 8904 35708 8910 35760
rect 9030 35748 9036 35760
rect 8991 35720 9036 35748
rect 9030 35708 9036 35720
rect 9088 35708 9094 35760
rect 16666 35708 16672 35760
rect 16724 35748 16730 35760
rect 25317 35751 25375 35757
rect 25317 35748 25329 35751
rect 16724 35720 25329 35748
rect 16724 35708 16730 35720
rect 25317 35717 25329 35720
rect 25363 35717 25375 35751
rect 28810 35748 28816 35760
rect 25317 35711 25375 35717
rect 28092 35720 28816 35748
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 19245 35683 19303 35689
rect 19245 35649 19257 35683
rect 19291 35680 19303 35683
rect 19518 35680 19524 35692
rect 19291 35652 19524 35680
rect 19291 35649 19303 35652
rect 19245 35643 19303 35649
rect 19518 35640 19524 35652
rect 19576 35640 19582 35692
rect 20165 35683 20223 35689
rect 20165 35649 20177 35683
rect 20211 35680 20223 35683
rect 20346 35680 20352 35692
rect 20211 35652 20352 35680
rect 20211 35649 20223 35652
rect 20165 35643 20223 35649
rect 20346 35640 20352 35652
rect 20404 35640 20410 35692
rect 20993 35683 21051 35689
rect 20993 35649 21005 35683
rect 21039 35680 21051 35683
rect 21266 35680 21272 35692
rect 21039 35652 21272 35680
rect 21039 35649 21051 35652
rect 20993 35643 21051 35649
rect 21266 35640 21272 35652
rect 21324 35640 21330 35692
rect 22370 35680 22376 35692
rect 22331 35652 22376 35680
rect 22370 35640 22376 35652
rect 22428 35640 22434 35692
rect 22629 35683 22687 35689
rect 22629 35680 22641 35683
rect 22480 35652 22641 35680
rect 15470 35572 15476 35624
rect 15528 35612 15534 35624
rect 20806 35612 20812 35624
rect 15528 35584 19840 35612
rect 20719 35584 20812 35612
rect 15528 35572 15534 35584
rect 19429 35547 19487 35553
rect 19429 35513 19441 35547
rect 19475 35544 19487 35547
rect 19702 35544 19708 35556
rect 19475 35516 19708 35544
rect 19475 35513 19487 35516
rect 19429 35507 19487 35513
rect 19702 35504 19708 35516
rect 19760 35504 19766 35556
rect 19812 35544 19840 35584
rect 20806 35572 20812 35584
rect 20864 35612 20870 35624
rect 22094 35612 22100 35624
rect 20864 35584 22100 35612
rect 20864 35572 20870 35584
rect 22094 35572 22100 35584
rect 22152 35572 22158 35624
rect 22278 35572 22284 35624
rect 22336 35612 22342 35624
rect 22480 35612 22508 35652
rect 22629 35649 22641 35652
rect 22675 35649 22687 35683
rect 22629 35643 22687 35649
rect 23198 35640 23204 35692
rect 23256 35680 23262 35692
rect 24762 35680 24768 35692
rect 23256 35652 23980 35680
rect 24723 35652 24768 35680
rect 23256 35640 23262 35652
rect 22336 35584 22508 35612
rect 22336 35572 22342 35584
rect 21358 35544 21364 35556
rect 19812 35516 21364 35544
rect 21358 35504 21364 35516
rect 21416 35504 21422 35556
rect 23952 35544 23980 35652
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 25041 35683 25099 35689
rect 25041 35649 25053 35683
rect 25087 35649 25099 35683
rect 25041 35643 25099 35649
rect 26973 35683 27031 35689
rect 26973 35649 26985 35683
rect 27019 35680 27031 35683
rect 27614 35680 27620 35692
rect 27019 35652 27620 35680
rect 27019 35649 27031 35652
rect 26973 35643 27031 35649
rect 24302 35612 24308 35624
rect 24263 35584 24308 35612
rect 24302 35572 24308 35584
rect 24360 35572 24366 35624
rect 25056 35544 25084 35643
rect 27614 35640 27620 35652
rect 27672 35640 27678 35692
rect 28092 35689 28120 35720
rect 28810 35708 28816 35720
rect 28868 35708 28874 35760
rect 27985 35683 28043 35689
rect 27985 35649 27997 35683
rect 28031 35649 28043 35683
rect 27985 35643 28043 35649
rect 28077 35683 28135 35689
rect 28077 35649 28089 35683
rect 28123 35649 28135 35683
rect 28077 35643 28135 35649
rect 28169 35683 28227 35689
rect 28169 35649 28181 35683
rect 28215 35649 28227 35683
rect 28169 35643 28227 35649
rect 28000 35612 28028 35643
rect 28184 35612 28212 35643
rect 28258 35640 28264 35692
rect 28316 35680 28322 35692
rect 28353 35683 28411 35689
rect 28353 35680 28365 35683
rect 28316 35652 28365 35680
rect 28316 35640 28322 35652
rect 28353 35649 28365 35652
rect 28399 35649 28411 35683
rect 29914 35680 29920 35692
rect 28353 35643 28411 35649
rect 28552 35652 29920 35680
rect 28552 35612 28580 35652
rect 29914 35640 29920 35652
rect 29972 35640 29978 35692
rect 30300 35624 30328 35776
rect 28810 35612 28816 35624
rect 28000 35584 28120 35612
rect 28184 35584 28580 35612
rect 28771 35584 28816 35612
rect 23952 35516 25084 35544
rect 28092 35544 28120 35584
rect 28810 35572 28816 35584
rect 28868 35572 28874 35624
rect 29086 35612 29092 35624
rect 29047 35584 29092 35612
rect 29086 35572 29092 35584
rect 29144 35572 29150 35624
rect 30282 35572 30288 35624
rect 30340 35572 30346 35624
rect 29104 35544 29132 35572
rect 28092 35516 29132 35544
rect 1397 35479 1455 35485
rect 1397 35445 1409 35479
rect 1443 35476 1455 35479
rect 3970 35476 3976 35488
rect 1443 35448 3976 35476
rect 1443 35445 1455 35448
rect 1397 35439 1455 35445
rect 3970 35436 3976 35448
rect 4028 35436 4034 35488
rect 9217 35479 9275 35485
rect 9217 35445 9229 35479
rect 9263 35476 9275 35479
rect 13354 35476 13360 35488
rect 9263 35448 13360 35476
rect 9263 35445 9275 35448
rect 9217 35439 9275 35445
rect 13354 35436 13360 35448
rect 13412 35436 13418 35488
rect 19794 35436 19800 35488
rect 19852 35476 19858 35488
rect 19981 35479 20039 35485
rect 19981 35476 19993 35479
rect 19852 35448 19993 35476
rect 19852 35436 19858 35448
rect 19981 35445 19993 35448
rect 20027 35445 20039 35479
rect 19981 35439 20039 35445
rect 26326 35436 26332 35488
rect 26384 35476 26390 35488
rect 26510 35476 26516 35488
rect 26384 35448 26516 35476
rect 26384 35436 26390 35448
rect 26510 35436 26516 35448
rect 26568 35436 26574 35488
rect 27157 35479 27215 35485
rect 27157 35445 27169 35479
rect 27203 35476 27215 35479
rect 27614 35476 27620 35488
rect 27203 35448 27620 35476
rect 27203 35445 27215 35448
rect 27157 35439 27215 35445
rect 27614 35436 27620 35448
rect 27672 35436 27678 35488
rect 1104 35386 30820 35408
rect 1104 35334 5915 35386
rect 5967 35334 5979 35386
rect 6031 35334 6043 35386
rect 6095 35334 6107 35386
rect 6159 35334 6171 35386
rect 6223 35334 15846 35386
rect 15898 35334 15910 35386
rect 15962 35334 15974 35386
rect 16026 35334 16038 35386
rect 16090 35334 16102 35386
rect 16154 35334 25776 35386
rect 25828 35334 25840 35386
rect 25892 35334 25904 35386
rect 25956 35334 25968 35386
rect 26020 35334 26032 35386
rect 26084 35334 30820 35386
rect 1104 35312 30820 35334
rect 9674 35232 9680 35284
rect 9732 35272 9738 35284
rect 10873 35275 10931 35281
rect 10873 35272 10885 35275
rect 9732 35244 10885 35272
rect 9732 35232 9738 35244
rect 10873 35241 10885 35244
rect 10919 35241 10931 35275
rect 10873 35235 10931 35241
rect 11606 35232 11612 35284
rect 11664 35272 11670 35284
rect 11701 35275 11759 35281
rect 11701 35272 11713 35275
rect 11664 35244 11713 35272
rect 11664 35232 11670 35244
rect 11701 35241 11713 35244
rect 11747 35241 11759 35275
rect 12342 35272 12348 35284
rect 12303 35244 12348 35272
rect 11701 35235 11759 35241
rect 12342 35232 12348 35244
rect 12400 35232 12406 35284
rect 13449 35275 13507 35281
rect 13449 35241 13461 35275
rect 13495 35272 13507 35275
rect 14090 35272 14096 35284
rect 13495 35244 14096 35272
rect 13495 35241 13507 35244
rect 13449 35235 13507 35241
rect 14090 35232 14096 35244
rect 14148 35232 14154 35284
rect 18049 35275 18107 35281
rect 18049 35241 18061 35275
rect 18095 35272 18107 35275
rect 19242 35272 19248 35284
rect 18095 35244 19248 35272
rect 18095 35241 18107 35244
rect 18049 35235 18107 35241
rect 19242 35232 19248 35244
rect 19300 35232 19306 35284
rect 19702 35272 19708 35284
rect 19352 35244 19708 35272
rect 16390 35164 16396 35216
rect 16448 35204 16454 35216
rect 16577 35207 16635 35213
rect 16577 35204 16589 35207
rect 16448 35176 16589 35204
rect 16448 35164 16454 35176
rect 16577 35173 16589 35176
rect 16623 35173 16635 35207
rect 16577 35167 16635 35173
rect 17037 35139 17095 35145
rect 17037 35105 17049 35139
rect 17083 35136 17095 35139
rect 17310 35136 17316 35148
rect 17083 35108 17316 35136
rect 17083 35105 17095 35108
rect 17037 35099 17095 35105
rect 17310 35096 17316 35108
rect 17368 35096 17374 35148
rect 18509 35139 18567 35145
rect 18509 35105 18521 35139
rect 18555 35136 18567 35139
rect 19352 35136 19380 35244
rect 19702 35232 19708 35244
rect 19760 35232 19766 35284
rect 20806 35272 20812 35284
rect 20767 35244 20812 35272
rect 20806 35232 20812 35244
rect 20864 35232 20870 35284
rect 23106 35232 23112 35284
rect 23164 35272 23170 35284
rect 23753 35275 23811 35281
rect 23753 35272 23765 35275
rect 23164 35244 23765 35272
rect 23164 35232 23170 35244
rect 23753 35241 23765 35244
rect 23799 35241 23811 35275
rect 23753 35235 23811 35241
rect 18555 35108 19380 35136
rect 23768 35136 23796 35235
rect 24118 35232 24124 35284
rect 24176 35272 24182 35284
rect 24581 35275 24639 35281
rect 24581 35272 24593 35275
rect 24176 35244 24593 35272
rect 24176 35232 24182 35244
rect 24581 35241 24593 35244
rect 24627 35272 24639 35275
rect 28810 35272 28816 35284
rect 24627 35244 28816 35272
rect 24627 35241 24639 35244
rect 24581 35235 24639 35241
rect 28810 35232 28816 35244
rect 28868 35232 28874 35284
rect 24762 35164 24768 35216
rect 24820 35204 24826 35216
rect 26973 35207 27031 35213
rect 26973 35204 26985 35207
rect 24820 35176 26985 35204
rect 24820 35164 24826 35176
rect 26973 35173 26985 35176
rect 27019 35173 27031 35207
rect 26973 35167 27031 35173
rect 23768 35108 24440 35136
rect 18555 35105 18567 35108
rect 18509 35099 18567 35105
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35028 1642 35080
rect 10318 35028 10324 35080
rect 10376 35068 10382 35080
rect 10689 35071 10747 35077
rect 10689 35068 10701 35071
rect 10376 35040 10701 35068
rect 10376 35028 10382 35040
rect 10689 35037 10701 35040
rect 10735 35037 10747 35071
rect 10689 35031 10747 35037
rect 11517 35071 11575 35077
rect 11517 35037 11529 35071
rect 11563 35037 11575 35071
rect 11517 35031 11575 35037
rect 12161 35071 12219 35077
rect 12161 35037 12173 35071
rect 12207 35068 12219 35071
rect 12207 35040 12434 35068
rect 12207 35037 12219 35040
rect 12161 35031 12219 35037
rect 10594 34960 10600 35012
rect 10652 35000 10658 35012
rect 11532 35000 11560 35031
rect 10652 34972 11560 35000
rect 12406 35000 12434 35040
rect 12618 35028 12624 35080
rect 12676 35068 12682 35080
rect 13265 35071 13323 35077
rect 13265 35068 13277 35071
rect 12676 35040 13277 35068
rect 12676 35028 12682 35040
rect 13265 35037 13277 35040
rect 13311 35037 13323 35071
rect 14550 35068 14556 35080
rect 14511 35040 14556 35068
rect 13265 35031 13323 35037
rect 14550 35028 14556 35040
rect 14608 35028 14614 35080
rect 14737 35071 14795 35077
rect 14737 35037 14749 35071
rect 14783 35068 14795 35071
rect 15102 35068 15108 35080
rect 14783 35040 15108 35068
rect 14783 35037 14795 35040
rect 14737 35031 14795 35037
rect 15102 35028 15108 35040
rect 15160 35068 15166 35080
rect 15841 35071 15899 35077
rect 15841 35068 15853 35071
rect 15160 35040 15853 35068
rect 15160 35028 15166 35040
rect 15841 35037 15853 35040
rect 15887 35037 15899 35071
rect 18598 35068 18604 35080
rect 18511 35040 18604 35068
rect 15841 35031 15899 35037
rect 18598 35028 18604 35040
rect 18656 35068 18662 35080
rect 18782 35068 18788 35080
rect 18656 35040 18788 35068
rect 18656 35028 18662 35040
rect 18782 35028 18788 35040
rect 18840 35028 18846 35080
rect 19429 35071 19487 35077
rect 19429 35037 19441 35071
rect 19475 35068 19487 35071
rect 20438 35068 20444 35080
rect 19475 35040 20444 35068
rect 19475 35037 19487 35040
rect 19429 35031 19487 35037
rect 20438 35028 20444 35040
rect 20496 35028 20502 35080
rect 21174 35028 21180 35080
rect 21232 35068 21238 35080
rect 21821 35071 21879 35077
rect 21821 35068 21833 35071
rect 21232 35040 21833 35068
rect 21232 35028 21238 35040
rect 21821 35037 21833 35040
rect 21867 35037 21879 35071
rect 22094 35068 22100 35080
rect 22055 35040 22100 35068
rect 21821 35031 21879 35037
rect 22094 35028 22100 35040
rect 22152 35028 22158 35080
rect 23661 35071 23719 35077
rect 23661 35037 23673 35071
rect 23707 35068 23719 35071
rect 23845 35071 23903 35077
rect 23707 35040 23796 35068
rect 23707 35037 23719 35040
rect 23661 35031 23719 35037
rect 14090 35000 14096 35012
rect 12406 34972 14096 35000
rect 10652 34960 10658 34972
rect 14090 34960 14096 34972
rect 14148 34960 14154 35012
rect 17129 35003 17187 35009
rect 17129 34969 17141 35003
rect 17175 35000 17187 35003
rect 17402 35000 17408 35012
rect 17175 34972 17408 35000
rect 17175 34969 17187 34972
rect 17129 34963 17187 34969
rect 17402 34960 17408 34972
rect 17460 34960 17466 35012
rect 19696 35003 19754 35009
rect 19696 34969 19708 35003
rect 19742 35000 19754 35003
rect 19794 35000 19800 35012
rect 19742 34972 19800 35000
rect 19742 34969 19754 34972
rect 19696 34963 19754 34969
rect 19794 34960 19800 34972
rect 19852 34960 19858 35012
rect 1397 34935 1455 34941
rect 1397 34901 1409 34935
rect 1443 34932 1455 34935
rect 4062 34932 4068 34944
rect 1443 34904 4068 34932
rect 1443 34901 1455 34904
rect 1397 34895 1455 34901
rect 4062 34892 4068 34904
rect 4120 34892 4126 34944
rect 16025 34935 16083 34941
rect 16025 34901 16037 34935
rect 16071 34932 16083 34935
rect 16942 34932 16948 34944
rect 16071 34904 16948 34932
rect 16071 34901 16083 34904
rect 16025 34895 16083 34901
rect 16942 34892 16948 34904
rect 17000 34892 17006 34944
rect 17037 34935 17095 34941
rect 17037 34901 17049 34935
rect 17083 34932 17095 34935
rect 17954 34932 17960 34944
rect 17083 34904 17960 34932
rect 17083 34901 17095 34904
rect 17037 34895 17095 34901
rect 17954 34892 17960 34904
rect 18012 34932 18018 34944
rect 18414 34932 18420 34944
rect 18012 34904 18420 34932
rect 18012 34892 18018 34904
rect 18414 34892 18420 34904
rect 18472 34892 18478 34944
rect 18509 34935 18567 34941
rect 18509 34901 18521 34935
rect 18555 34932 18567 34935
rect 19058 34932 19064 34944
rect 18555 34904 19064 34932
rect 18555 34901 18567 34904
rect 18509 34895 18567 34901
rect 19058 34892 19064 34904
rect 19116 34892 19122 34944
rect 21818 34892 21824 34944
rect 21876 34932 21882 34944
rect 21913 34935 21971 34941
rect 21913 34932 21925 34935
rect 21876 34904 21925 34932
rect 21876 34892 21882 34904
rect 21913 34901 21925 34904
rect 21959 34901 21971 34935
rect 23768 34932 23796 35040
rect 23845 35037 23857 35071
rect 23891 35068 23903 35071
rect 24026 35068 24032 35080
rect 23891 35040 24032 35068
rect 23891 35037 23903 35040
rect 23845 35031 23903 35037
rect 24026 35028 24032 35040
rect 24084 35028 24090 35080
rect 24412 35077 24440 35108
rect 26326 35096 26332 35148
rect 26384 35136 26390 35148
rect 26384 35108 29868 35136
rect 26384 35096 26390 35108
rect 24397 35071 24455 35077
rect 24397 35037 24409 35071
rect 24443 35037 24455 35071
rect 27062 35068 27068 35080
rect 27023 35040 27068 35068
rect 24397 35031 24455 35037
rect 27062 35028 27068 35040
rect 27120 35028 27126 35080
rect 27617 35071 27675 35077
rect 27617 35037 27629 35071
rect 27663 35037 27675 35071
rect 28166 35068 28172 35080
rect 28127 35040 28172 35068
rect 27617 35031 27675 35037
rect 27632 35000 27660 35031
rect 28166 35028 28172 35040
rect 28224 35028 28230 35080
rect 29840 35077 29868 35108
rect 29825 35071 29883 35077
rect 29825 35037 29837 35071
rect 29871 35037 29883 35071
rect 29825 35031 29883 35037
rect 30006 35028 30012 35080
rect 30064 35068 30070 35080
rect 30374 35068 30380 35080
rect 30064 35040 30380 35068
rect 30064 35028 30070 35040
rect 30374 35028 30380 35040
rect 30432 35028 30438 35080
rect 28258 35000 28264 35012
rect 27632 34972 28264 35000
rect 28258 34960 28264 34972
rect 28316 35000 28322 35012
rect 28353 35003 28411 35009
rect 28353 35000 28365 35003
rect 28316 34972 28365 35000
rect 28316 34960 28322 34972
rect 28353 34969 28365 34972
rect 28399 34969 28411 35003
rect 28353 34963 28411 34969
rect 27614 34932 27620 34944
rect 23768 34904 27620 34932
rect 21913 34895 21971 34901
rect 27614 34892 27620 34904
rect 27672 34892 27678 34944
rect 30006 34932 30012 34944
rect 29967 34904 30012 34932
rect 30006 34892 30012 34904
rect 30064 34892 30070 34944
rect 1104 34842 30820 34864
rect 1104 34790 10880 34842
rect 10932 34790 10944 34842
rect 10996 34790 11008 34842
rect 11060 34790 11072 34842
rect 11124 34790 11136 34842
rect 11188 34790 20811 34842
rect 20863 34790 20875 34842
rect 20927 34790 20939 34842
rect 20991 34790 21003 34842
rect 21055 34790 21067 34842
rect 21119 34790 30820 34842
rect 1104 34768 30820 34790
rect 1397 34731 1455 34737
rect 1397 34697 1409 34731
rect 1443 34728 1455 34731
rect 1443 34700 2774 34728
rect 1443 34697 1455 34700
rect 1397 34691 1455 34697
rect 2746 34660 2774 34700
rect 9766 34688 9772 34740
rect 9824 34728 9830 34740
rect 9861 34731 9919 34737
rect 9861 34728 9873 34731
rect 9824 34700 9873 34728
rect 9824 34688 9830 34700
rect 9861 34697 9873 34700
rect 9907 34697 9919 34731
rect 9861 34691 9919 34697
rect 13906 34688 13912 34740
rect 13964 34728 13970 34740
rect 14277 34731 14335 34737
rect 14277 34728 14289 34731
rect 13964 34700 14289 34728
rect 13964 34688 13970 34700
rect 14277 34697 14289 34700
rect 14323 34697 14335 34731
rect 14277 34691 14335 34697
rect 17313 34731 17371 34737
rect 17313 34697 17325 34731
rect 17359 34728 17371 34731
rect 17954 34728 17960 34740
rect 17359 34700 17960 34728
rect 17359 34697 17371 34700
rect 17313 34691 17371 34697
rect 17954 34688 17960 34700
rect 18012 34688 18018 34740
rect 19058 34728 19064 34740
rect 19019 34700 19064 34728
rect 19058 34688 19064 34700
rect 19116 34688 19122 34740
rect 20438 34728 20444 34740
rect 20399 34700 20444 34728
rect 20438 34688 20444 34700
rect 20496 34688 20502 34740
rect 27614 34688 27620 34740
rect 27672 34728 27678 34740
rect 28169 34731 28227 34737
rect 28169 34728 28181 34731
rect 27672 34700 28181 34728
rect 27672 34688 27678 34700
rect 28169 34697 28181 34700
rect 28215 34697 28227 34731
rect 28902 34728 28908 34740
rect 28863 34700 28908 34728
rect 28169 34691 28227 34697
rect 28902 34688 28908 34700
rect 28960 34688 28966 34740
rect 29178 34688 29184 34740
rect 29236 34728 29242 34740
rect 29546 34728 29552 34740
rect 29236 34700 29552 34728
rect 29236 34688 29242 34700
rect 29546 34688 29552 34700
rect 29604 34688 29610 34740
rect 30834 34728 30840 34740
rect 29840 34700 30840 34728
rect 10413 34663 10471 34669
rect 2746 34632 9904 34660
rect 9876 34604 9904 34632
rect 10413 34629 10425 34663
rect 10459 34660 10471 34663
rect 13170 34660 13176 34672
rect 10459 34632 13176 34660
rect 10459 34629 10471 34632
rect 10413 34623 10471 34629
rect 13170 34620 13176 34632
rect 13228 34620 13234 34672
rect 15746 34620 15752 34672
rect 15804 34660 15810 34672
rect 15933 34663 15991 34669
rect 15933 34660 15945 34663
rect 15804 34632 15945 34660
rect 15804 34620 15810 34632
rect 15933 34629 15945 34632
rect 15979 34629 15991 34663
rect 15933 34623 15991 34629
rect 18141 34663 18199 34669
rect 18141 34629 18153 34663
rect 18187 34660 18199 34663
rect 18690 34660 18696 34672
rect 18187 34632 18696 34660
rect 18187 34629 18199 34632
rect 18141 34623 18199 34629
rect 18690 34620 18696 34632
rect 18748 34620 18754 34672
rect 18969 34663 19027 34669
rect 18969 34629 18981 34663
rect 19015 34660 19027 34663
rect 20070 34660 20076 34672
rect 19015 34632 20076 34660
rect 19015 34629 19027 34632
rect 18969 34623 19027 34629
rect 20070 34620 20076 34632
rect 20128 34620 20134 34672
rect 24946 34620 24952 34672
rect 25004 34660 25010 34672
rect 27341 34663 27399 34669
rect 27341 34660 27353 34663
rect 25004 34632 27353 34660
rect 25004 34620 25010 34632
rect 27341 34629 27353 34632
rect 27387 34629 27399 34663
rect 27341 34623 27399 34629
rect 27448 34632 28028 34660
rect 1394 34552 1400 34604
rect 1452 34592 1458 34604
rect 1581 34595 1639 34601
rect 1581 34592 1593 34595
rect 1452 34564 1593 34592
rect 1452 34552 1458 34564
rect 1581 34561 1593 34564
rect 1627 34561 1639 34595
rect 9674 34592 9680 34604
rect 9635 34564 9680 34592
rect 1581 34555 1639 34561
rect 9674 34552 9680 34564
rect 9732 34552 9738 34604
rect 9858 34552 9864 34604
rect 9916 34552 9922 34604
rect 11609 34595 11667 34601
rect 11609 34561 11621 34595
rect 11655 34561 11667 34595
rect 11609 34555 11667 34561
rect 12345 34595 12403 34601
rect 12345 34561 12357 34595
rect 12391 34592 12403 34595
rect 12986 34592 12992 34604
rect 12391 34564 12992 34592
rect 12391 34561 12403 34564
rect 12345 34555 12403 34561
rect 11624 34524 11652 34555
rect 12986 34552 12992 34564
rect 13044 34552 13050 34604
rect 13081 34595 13139 34601
rect 13081 34561 13093 34595
rect 13127 34592 13139 34595
rect 13998 34592 14004 34604
rect 13127 34564 14004 34592
rect 13127 34561 13139 34564
rect 13081 34555 13139 34561
rect 13998 34552 14004 34564
rect 14056 34552 14062 34604
rect 14090 34552 14096 34604
rect 14148 34592 14154 34604
rect 14734 34592 14740 34604
rect 14148 34564 14193 34592
rect 14695 34564 14740 34592
rect 14148 34552 14154 34564
rect 14734 34552 14740 34564
rect 14792 34552 14798 34604
rect 19610 34592 19616 34604
rect 19571 34564 19616 34592
rect 19610 34552 19616 34564
rect 19668 34552 19674 34604
rect 20254 34592 20260 34604
rect 20215 34564 20260 34592
rect 20254 34552 20260 34564
rect 20312 34552 20318 34604
rect 27062 34552 27068 34604
rect 27120 34592 27126 34604
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 27120 34564 27169 34592
rect 27120 34552 27126 34564
rect 27157 34561 27169 34564
rect 27203 34592 27215 34595
rect 27448 34592 27476 34632
rect 28000 34601 28028 34632
rect 27203 34564 27476 34592
rect 27985 34595 28043 34601
rect 27203 34561 27215 34564
rect 27157 34555 27215 34561
rect 27985 34561 27997 34595
rect 28031 34561 28043 34595
rect 27985 34555 28043 34561
rect 28721 34595 28779 34601
rect 28721 34561 28733 34595
rect 28767 34561 28779 34595
rect 28721 34555 28779 34561
rect 13265 34527 13323 34533
rect 11624 34496 12434 34524
rect 10597 34459 10655 34465
rect 10597 34425 10609 34459
rect 10643 34456 10655 34459
rect 10778 34456 10784 34468
rect 10643 34428 10784 34456
rect 10643 34425 10655 34428
rect 10597 34419 10655 34425
rect 10778 34416 10784 34428
rect 10836 34416 10842 34468
rect 12406 34456 12434 34496
rect 13265 34493 13277 34527
rect 13311 34524 13323 34527
rect 14108 34524 14136 34552
rect 13311 34496 14136 34524
rect 16117 34527 16175 34533
rect 13311 34493 13323 34496
rect 13265 34487 13323 34493
rect 16117 34493 16129 34527
rect 16163 34524 16175 34527
rect 17310 34524 17316 34536
rect 16163 34496 17316 34524
rect 16163 34493 16175 34496
rect 16117 34487 16175 34493
rect 17310 34484 17316 34496
rect 17368 34484 17374 34536
rect 17402 34484 17408 34536
rect 17460 34524 17466 34536
rect 18322 34524 18328 34536
rect 17460 34496 17505 34524
rect 18283 34496 18328 34524
rect 17460 34484 17466 34496
rect 18322 34484 18328 34496
rect 18380 34484 18386 34536
rect 19886 34484 19892 34536
rect 19944 34524 19950 34536
rect 20438 34524 20444 34536
rect 19944 34496 20444 34524
rect 19944 34484 19950 34496
rect 20438 34484 20444 34496
rect 20496 34484 20502 34536
rect 26234 34484 26240 34536
rect 26292 34524 26298 34536
rect 28736 34524 28764 34555
rect 29086 34552 29092 34604
rect 29144 34592 29150 34604
rect 29840 34601 29868 34700
rect 30834 34688 30840 34700
rect 30892 34688 30898 34740
rect 29733 34595 29791 34601
rect 29733 34592 29745 34595
rect 29144 34564 29745 34592
rect 29144 34552 29150 34564
rect 29733 34561 29745 34564
rect 29779 34561 29791 34595
rect 29733 34555 29791 34561
rect 29825 34595 29883 34601
rect 29825 34561 29837 34595
rect 29871 34561 29883 34595
rect 29825 34555 29883 34561
rect 29917 34595 29975 34601
rect 29917 34561 29929 34595
rect 29963 34561 29975 34595
rect 30101 34595 30159 34601
rect 30101 34592 30113 34595
rect 29917 34555 29975 34561
rect 30024 34564 30113 34592
rect 26292 34496 28764 34524
rect 26292 34484 26298 34496
rect 28994 34484 29000 34536
rect 29052 34524 29058 34536
rect 29052 34496 29500 34524
rect 29052 34484 29058 34496
rect 13814 34456 13820 34468
rect 12406 34428 13820 34456
rect 13814 34416 13820 34428
rect 13872 34416 13878 34468
rect 27154 34416 27160 34468
rect 27212 34456 27218 34468
rect 27522 34456 27528 34468
rect 27212 34428 27528 34456
rect 27212 34416 27218 34428
rect 27522 34416 27528 34428
rect 27580 34416 27586 34468
rect 29472 34456 29500 34496
rect 29546 34484 29552 34536
rect 29604 34524 29610 34536
rect 29932 34524 29960 34555
rect 29604 34496 29960 34524
rect 29604 34484 29610 34496
rect 30024 34456 30052 34564
rect 30101 34561 30113 34564
rect 30147 34561 30159 34595
rect 30101 34555 30159 34561
rect 29472 34428 30052 34456
rect 11790 34388 11796 34400
rect 11751 34360 11796 34388
rect 11790 34348 11796 34360
rect 11848 34348 11854 34400
rect 11882 34348 11888 34400
rect 11940 34388 11946 34400
rect 12437 34391 12495 34397
rect 12437 34388 12449 34391
rect 11940 34360 12449 34388
rect 11940 34348 11946 34360
rect 12437 34357 12449 34360
rect 12483 34357 12495 34391
rect 14918 34388 14924 34400
rect 14879 34360 14924 34388
rect 12437 34351 12495 34357
rect 14918 34348 14924 34360
rect 14976 34348 14982 34400
rect 16853 34391 16911 34397
rect 16853 34357 16865 34391
rect 16899 34388 16911 34391
rect 17218 34388 17224 34400
rect 16899 34360 17224 34388
rect 16899 34357 16911 34360
rect 16853 34351 16911 34357
rect 17218 34348 17224 34360
rect 17276 34348 17282 34400
rect 17494 34348 17500 34400
rect 17552 34388 17558 34400
rect 19797 34391 19855 34397
rect 19797 34388 19809 34391
rect 17552 34360 19809 34388
rect 17552 34348 17558 34360
rect 19797 34357 19809 34360
rect 19843 34357 19855 34391
rect 19797 34351 19855 34357
rect 21726 34348 21732 34400
rect 21784 34388 21790 34400
rect 24762 34388 24768 34400
rect 21784 34360 24768 34388
rect 21784 34348 21790 34360
rect 24762 34348 24768 34360
rect 24820 34348 24826 34400
rect 26878 34348 26884 34400
rect 26936 34388 26942 34400
rect 27433 34391 27491 34397
rect 27433 34388 27445 34391
rect 26936 34360 27445 34388
rect 26936 34348 26942 34360
rect 27433 34357 27445 34360
rect 27479 34357 27491 34391
rect 27433 34351 27491 34357
rect 29457 34391 29515 34397
rect 29457 34357 29469 34391
rect 29503 34388 29515 34391
rect 29822 34388 29828 34400
rect 29503 34360 29828 34388
rect 29503 34357 29515 34360
rect 29457 34351 29515 34357
rect 29822 34348 29828 34360
rect 29880 34348 29886 34400
rect 1104 34298 30820 34320
rect 1104 34246 5915 34298
rect 5967 34246 5979 34298
rect 6031 34246 6043 34298
rect 6095 34246 6107 34298
rect 6159 34246 6171 34298
rect 6223 34246 15846 34298
rect 15898 34246 15910 34298
rect 15962 34246 15974 34298
rect 16026 34246 16038 34298
rect 16090 34246 16102 34298
rect 16154 34246 25776 34298
rect 25828 34246 25840 34298
rect 25892 34246 25904 34298
rect 25956 34246 25968 34298
rect 26020 34246 26032 34298
rect 26084 34246 30820 34298
rect 1104 34224 30820 34246
rect 9674 34144 9680 34196
rect 9732 34184 9738 34196
rect 10505 34187 10563 34193
rect 10505 34184 10517 34187
rect 9732 34156 10517 34184
rect 9732 34144 9738 34156
rect 10505 34153 10517 34156
rect 10551 34153 10563 34187
rect 10505 34147 10563 34153
rect 13998 34144 14004 34196
rect 14056 34184 14062 34196
rect 16577 34187 16635 34193
rect 16577 34184 16589 34187
rect 14056 34156 16589 34184
rect 14056 34144 14062 34156
rect 16577 34153 16589 34156
rect 16623 34184 16635 34187
rect 16623 34156 19380 34184
rect 16623 34153 16635 34156
rect 16577 34147 16635 34153
rect 12986 34076 12992 34128
rect 13044 34116 13050 34128
rect 13722 34116 13728 34128
rect 13044 34088 13728 34116
rect 13044 34076 13050 34088
rect 13722 34076 13728 34088
rect 13780 34076 13786 34128
rect 17589 34119 17647 34125
rect 17589 34085 17601 34119
rect 17635 34116 17647 34119
rect 17862 34116 17868 34128
rect 17635 34088 17868 34116
rect 17635 34085 17647 34088
rect 17589 34079 17647 34085
rect 17862 34076 17868 34088
rect 17920 34076 17926 34128
rect 11057 34051 11115 34057
rect 11057 34017 11069 34051
rect 11103 34048 11115 34051
rect 11238 34048 11244 34060
rect 11103 34020 11244 34048
rect 11103 34017 11115 34020
rect 11057 34011 11115 34017
rect 11238 34008 11244 34020
rect 11296 34048 11302 34060
rect 11882 34048 11888 34060
rect 11296 34020 11888 34048
rect 11296 34008 11302 34020
rect 11882 34008 11888 34020
rect 11940 34008 11946 34060
rect 12713 34051 12771 34057
rect 12713 34017 12725 34051
rect 12759 34048 12771 34051
rect 13078 34048 13084 34060
rect 12759 34020 13084 34048
rect 12759 34017 12771 34020
rect 12713 34011 12771 34017
rect 13078 34008 13084 34020
rect 13136 34008 13142 34060
rect 17310 34008 17316 34060
rect 17368 34048 17374 34060
rect 17957 34051 18015 34057
rect 17957 34048 17969 34051
rect 17368 34020 17969 34048
rect 17368 34008 17374 34020
rect 17957 34017 17969 34020
rect 18003 34017 18015 34051
rect 17957 34011 18015 34017
rect 1578 33980 1584 33992
rect 1539 33952 1584 33980
rect 1578 33940 1584 33952
rect 1636 33940 1642 33992
rect 10778 33980 10784 33992
rect 10739 33952 10784 33980
rect 10778 33940 10784 33952
rect 10836 33940 10842 33992
rect 13357 33983 13415 33989
rect 13357 33949 13369 33983
rect 13403 33980 13415 33983
rect 13814 33980 13820 33992
rect 13403 33952 13820 33980
rect 13403 33949 13415 33952
rect 13357 33943 13415 33949
rect 13814 33940 13820 33952
rect 13872 33980 13878 33992
rect 15102 33980 15108 33992
rect 13872 33952 15108 33980
rect 13872 33940 13878 33952
rect 15102 33940 15108 33952
rect 15160 33940 15166 33992
rect 15289 33983 15347 33989
rect 15289 33949 15301 33983
rect 15335 33980 15347 33983
rect 17494 33980 17500 33992
rect 15335 33952 17500 33980
rect 15335 33949 15347 33952
rect 15289 33943 15347 33949
rect 17494 33940 17500 33952
rect 17552 33940 17558 33992
rect 12805 33915 12863 33921
rect 12805 33881 12817 33915
rect 12851 33912 12863 33915
rect 12986 33912 12992 33924
rect 12851 33884 12992 33912
rect 12851 33881 12863 33884
rect 12805 33875 12863 33881
rect 12986 33872 12992 33884
rect 13044 33912 13050 33924
rect 13044 33884 13676 33912
rect 13044 33872 13050 33884
rect 1397 33847 1455 33853
rect 1397 33813 1409 33847
rect 1443 33844 1455 33847
rect 9950 33844 9956 33856
rect 1443 33816 9956 33844
rect 1443 33813 1455 33816
rect 1397 33807 1455 33813
rect 9950 33804 9956 33816
rect 10008 33804 10014 33856
rect 10965 33847 11023 33853
rect 10965 33813 10977 33847
rect 11011 33844 11023 33847
rect 11514 33844 11520 33856
rect 11011 33816 11520 33844
rect 11011 33813 11023 33816
rect 10965 33807 11023 33813
rect 11514 33804 11520 33816
rect 11572 33804 11578 33856
rect 11606 33804 11612 33856
rect 11664 33844 11670 33856
rect 12235 33847 12293 33853
rect 12235 33844 12247 33847
rect 11664 33816 12247 33844
rect 11664 33804 11670 33816
rect 12235 33813 12247 33816
rect 12281 33813 12293 33847
rect 12235 33807 12293 33813
rect 12342 33804 12348 33856
rect 12400 33844 12406 33856
rect 12713 33847 12771 33853
rect 12713 33844 12725 33847
rect 12400 33816 12725 33844
rect 12400 33804 12406 33816
rect 12713 33813 12725 33816
rect 12759 33813 12771 33847
rect 13538 33844 13544 33856
rect 13499 33816 13544 33844
rect 12713 33807 12771 33813
rect 13538 33804 13544 33816
rect 13596 33804 13602 33856
rect 13648 33844 13676 33884
rect 13722 33872 13728 33924
rect 13780 33912 13786 33924
rect 14185 33915 14243 33921
rect 14185 33912 14197 33915
rect 13780 33884 14197 33912
rect 13780 33872 13786 33884
rect 14185 33881 14197 33884
rect 14231 33881 14243 33915
rect 18046 33912 18052 33924
rect 18007 33884 18052 33912
rect 14185 33875 14243 33881
rect 18046 33872 18052 33884
rect 18104 33872 18110 33924
rect 19352 33921 19380 34156
rect 19610 34144 19616 34196
rect 19668 34184 19674 34196
rect 20073 34187 20131 34193
rect 20073 34184 20085 34187
rect 19668 34156 20085 34184
rect 19668 34144 19674 34156
rect 20073 34153 20085 34156
rect 20119 34153 20131 34187
rect 20073 34147 20131 34153
rect 25038 34144 25044 34196
rect 25096 34184 25102 34196
rect 26694 34184 26700 34196
rect 25096 34156 26004 34184
rect 25096 34144 25102 34156
rect 25976 34128 26004 34156
rect 26344 34156 26700 34184
rect 19518 34076 19524 34128
rect 19576 34116 19582 34128
rect 19886 34116 19892 34128
rect 19576 34088 19892 34116
rect 19576 34076 19582 34088
rect 19886 34076 19892 34088
rect 19944 34076 19950 34128
rect 25133 34119 25191 34125
rect 25133 34085 25145 34119
rect 25179 34116 25191 34119
rect 25590 34116 25596 34128
rect 25179 34088 25596 34116
rect 25179 34085 25191 34088
rect 25133 34079 25191 34085
rect 25590 34076 25596 34088
rect 25648 34076 25654 34128
rect 25958 34076 25964 34128
rect 26016 34076 26022 34128
rect 26344 34125 26372 34156
rect 26694 34144 26700 34156
rect 26752 34144 26758 34196
rect 28166 34184 28172 34196
rect 28127 34156 28172 34184
rect 28166 34144 28172 34156
rect 28224 34144 28230 34196
rect 26329 34119 26387 34125
rect 26329 34085 26341 34119
rect 26375 34085 26387 34119
rect 26329 34079 26387 34085
rect 24854 34008 24860 34060
rect 24912 34008 24918 34060
rect 26694 34048 26700 34060
rect 25608 34020 26700 34048
rect 19978 33980 19984 33992
rect 19939 33952 19984 33980
rect 19978 33940 19984 33952
rect 20036 33940 20042 33992
rect 23290 33940 23296 33992
rect 23348 33980 23354 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 23348 33952 24593 33980
rect 23348 33940 23354 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33980 24823 33983
rect 24872 33980 24900 34008
rect 24811 33952 24900 33980
rect 24949 33983 25007 33989
rect 24811 33949 24823 33952
rect 24765 33943 24823 33949
rect 24949 33949 24961 33983
rect 24995 33980 25007 33983
rect 25038 33980 25044 33992
rect 24995 33952 25044 33980
rect 24995 33949 25007 33952
rect 24949 33943 25007 33949
rect 25038 33940 25044 33952
rect 25096 33940 25102 33992
rect 18141 33915 18199 33921
rect 18141 33881 18153 33915
rect 18187 33881 18199 33915
rect 18141 33875 18199 33881
rect 19337 33915 19395 33921
rect 19337 33881 19349 33915
rect 19383 33881 19395 33915
rect 19337 33875 19395 33881
rect 24857 33915 24915 33921
rect 24857 33881 24869 33915
rect 24903 33912 24915 33915
rect 25608 33912 25636 34020
rect 26694 34008 26700 34020
rect 26752 34008 26758 34060
rect 25774 33980 25780 33992
rect 25735 33952 25780 33980
rect 25774 33940 25780 33952
rect 25832 33940 25838 33992
rect 26145 33983 26203 33989
rect 26145 33949 26157 33983
rect 26191 33980 26203 33983
rect 26878 33980 26884 33992
rect 26191 33952 26884 33980
rect 26191 33949 26203 33952
rect 26145 33943 26203 33949
rect 26878 33940 26884 33952
rect 26936 33940 26942 33992
rect 27982 33980 27988 33992
rect 27943 33952 27988 33980
rect 27982 33940 27988 33952
rect 28040 33940 28046 33992
rect 28721 33983 28779 33989
rect 28721 33949 28733 33983
rect 28767 33980 28779 33983
rect 28810 33980 28816 33992
rect 28767 33952 28816 33980
rect 28767 33949 28779 33952
rect 28721 33943 28779 33949
rect 28810 33940 28816 33952
rect 28868 33940 28874 33992
rect 29822 33980 29828 33992
rect 29783 33952 29828 33980
rect 29822 33940 29828 33952
rect 29880 33940 29886 33992
rect 24903 33884 25636 33912
rect 24903 33881 24915 33884
rect 24857 33875 24915 33881
rect 14277 33847 14335 33853
rect 14277 33844 14289 33847
rect 13648 33816 14289 33844
rect 14277 33813 14289 33816
rect 14323 33813 14335 33847
rect 14277 33807 14335 33813
rect 17402 33804 17408 33856
rect 17460 33844 17466 33856
rect 18156 33844 18184 33875
rect 25682 33872 25688 33924
rect 25740 33912 25746 33924
rect 25961 33915 26019 33921
rect 25961 33912 25973 33915
rect 25740 33884 25973 33912
rect 25740 33872 25746 33884
rect 25961 33881 25973 33884
rect 26007 33881 26019 33915
rect 25961 33875 26019 33881
rect 26053 33915 26111 33921
rect 26053 33881 26065 33915
rect 26099 33912 26111 33915
rect 27246 33912 27252 33924
rect 26099 33884 27252 33912
rect 26099 33881 26111 33884
rect 26053 33875 26111 33881
rect 27246 33872 27252 33884
rect 27304 33872 27310 33924
rect 19426 33844 19432 33856
rect 17460 33816 18184 33844
rect 19387 33816 19432 33844
rect 17460 33804 17466 33816
rect 19426 33804 19432 33816
rect 19484 33804 19490 33856
rect 28902 33844 28908 33856
rect 28863 33816 28908 33844
rect 28902 33804 28908 33816
rect 28960 33804 28966 33856
rect 29362 33804 29368 33856
rect 29420 33844 29426 33856
rect 29822 33844 29828 33856
rect 29420 33816 29828 33844
rect 29420 33804 29426 33816
rect 29822 33804 29828 33816
rect 29880 33804 29886 33856
rect 30006 33844 30012 33856
rect 29967 33816 30012 33844
rect 30006 33804 30012 33816
rect 30064 33804 30070 33856
rect 1104 33754 30820 33776
rect 1104 33702 10880 33754
rect 10932 33702 10944 33754
rect 10996 33702 11008 33754
rect 11060 33702 11072 33754
rect 11124 33702 11136 33754
rect 11188 33702 20811 33754
rect 20863 33702 20875 33754
rect 20927 33702 20939 33754
rect 20991 33702 21003 33754
rect 21055 33702 21067 33754
rect 21119 33702 30820 33754
rect 1104 33680 30820 33702
rect 11793 33643 11851 33649
rect 11793 33609 11805 33643
rect 11839 33640 11851 33643
rect 12066 33640 12072 33652
rect 11839 33612 12072 33640
rect 11839 33609 11851 33612
rect 11793 33603 11851 33609
rect 12066 33600 12072 33612
rect 12124 33600 12130 33652
rect 13722 33600 13728 33652
rect 13780 33640 13786 33652
rect 15473 33643 15531 33649
rect 13780 33612 15424 33640
rect 13780 33600 13786 33612
rect 9769 33575 9827 33581
rect 9769 33541 9781 33575
rect 9815 33572 9827 33575
rect 10781 33575 10839 33581
rect 10781 33572 10793 33575
rect 9815 33544 10793 33572
rect 9815 33541 9827 33544
rect 9769 33535 9827 33541
rect 10781 33541 10793 33544
rect 10827 33572 10839 33575
rect 11514 33572 11520 33584
rect 10827 33544 11520 33572
rect 10827 33541 10839 33544
rect 10781 33535 10839 33541
rect 11514 33532 11520 33544
rect 11572 33532 11578 33584
rect 13081 33575 13139 33581
rect 13081 33541 13093 33575
rect 13127 33572 13139 33575
rect 13262 33572 13268 33584
rect 13127 33544 13268 33572
rect 13127 33541 13139 33544
rect 13081 33535 13139 33541
rect 13262 33532 13268 33544
rect 13320 33572 13326 33584
rect 14277 33575 14335 33581
rect 14277 33572 14289 33575
rect 13320 33544 14289 33572
rect 13320 33532 13326 33544
rect 14277 33541 14289 33544
rect 14323 33541 14335 33575
rect 15396 33572 15424 33612
rect 15473 33609 15485 33643
rect 15519 33640 15531 33643
rect 17310 33640 17316 33652
rect 15519 33612 17316 33640
rect 15519 33609 15531 33612
rect 15473 33603 15531 33609
rect 17310 33600 17316 33612
rect 17368 33640 17374 33652
rect 17589 33643 17647 33649
rect 17589 33640 17601 33643
rect 17368 33612 17601 33640
rect 17368 33600 17374 33612
rect 17589 33609 17601 33612
rect 17635 33609 17647 33643
rect 17589 33603 17647 33609
rect 24762 33600 24768 33652
rect 24820 33640 24826 33652
rect 26234 33640 26240 33652
rect 24820 33612 25728 33640
rect 26195 33612 26240 33640
rect 24820 33600 24826 33612
rect 16761 33575 16819 33581
rect 16761 33572 16773 33575
rect 15396 33544 16773 33572
rect 14277 33535 14335 33541
rect 16761 33541 16773 33544
rect 16807 33541 16819 33575
rect 16761 33535 16819 33541
rect 1394 33464 1400 33516
rect 1452 33504 1458 33516
rect 1581 33507 1639 33513
rect 1581 33504 1593 33507
rect 1452 33476 1593 33504
rect 1452 33464 1458 33476
rect 1581 33473 1593 33476
rect 1627 33473 1639 33507
rect 1581 33467 1639 33473
rect 9585 33507 9643 33513
rect 9585 33473 9597 33507
rect 9631 33473 9643 33507
rect 9585 33467 9643 33473
rect 10873 33507 10931 33513
rect 10873 33473 10885 33507
rect 10919 33504 10931 33507
rect 11238 33504 11244 33516
rect 10919 33476 11244 33504
rect 10919 33473 10931 33476
rect 10873 33467 10931 33473
rect 9600 33436 9628 33467
rect 11238 33464 11244 33476
rect 11296 33464 11302 33516
rect 11606 33504 11612 33516
rect 11567 33476 11612 33504
rect 11606 33464 11612 33476
rect 11664 33464 11670 33516
rect 12986 33464 12992 33516
rect 13044 33504 13050 33516
rect 13173 33507 13231 33513
rect 13173 33504 13185 33507
rect 13044 33476 13185 33504
rect 13044 33464 13050 33476
rect 13173 33473 13185 33476
rect 13219 33473 13231 33507
rect 13173 33467 13231 33473
rect 14093 33507 14151 33513
rect 14093 33473 14105 33507
rect 14139 33504 14151 33507
rect 15289 33507 15347 33513
rect 15289 33504 15301 33507
rect 14139 33476 15301 33504
rect 14139 33473 14151 33476
rect 14093 33467 14151 33473
rect 15289 33473 15301 33476
rect 15335 33504 15347 33507
rect 16206 33504 16212 33516
rect 15335 33476 16212 33504
rect 15335 33473 15347 33476
rect 15289 33467 15347 33473
rect 16206 33464 16212 33476
rect 16264 33464 16270 33516
rect 16776 33504 16804 33535
rect 16942 33532 16948 33584
rect 17000 33572 17006 33584
rect 18233 33575 18291 33581
rect 18233 33572 18245 33575
rect 17000 33544 18245 33572
rect 17000 33532 17006 33544
rect 18233 33541 18245 33544
rect 18279 33541 18291 33575
rect 18233 33535 18291 33541
rect 19518 33532 19524 33584
rect 19576 33572 19582 33584
rect 19886 33572 19892 33584
rect 19576 33544 19892 33572
rect 19576 33532 19582 33544
rect 19886 33532 19892 33544
rect 19944 33532 19950 33584
rect 24949 33575 25007 33581
rect 24949 33541 24961 33575
rect 24995 33572 25007 33575
rect 25130 33572 25136 33584
rect 24995 33544 25136 33572
rect 24995 33541 25007 33544
rect 24949 33535 25007 33541
rect 25130 33532 25136 33544
rect 25188 33532 25194 33584
rect 17494 33504 17500 33516
rect 16776 33476 17356 33504
rect 17455 33476 17500 33504
rect 10778 33436 10784 33448
rect 9600 33408 10640 33436
rect 10739 33408 10784 33436
rect 10318 33368 10324 33380
rect 10279 33340 10324 33368
rect 10318 33328 10324 33340
rect 10376 33328 10382 33380
rect 10612 33368 10640 33408
rect 10778 33396 10784 33408
rect 10836 33396 10842 33448
rect 13078 33436 13084 33448
rect 13039 33408 13084 33436
rect 13078 33396 13084 33408
rect 13136 33396 13142 33448
rect 14369 33439 14427 33445
rect 14369 33405 14381 33439
rect 14415 33436 14427 33439
rect 15194 33436 15200 33448
rect 14415 33408 15200 33436
rect 14415 33405 14427 33408
rect 14369 33399 14427 33405
rect 15194 33396 15200 33408
rect 15252 33436 15258 33448
rect 15565 33439 15623 33445
rect 15565 33436 15577 33439
rect 15252 33408 15577 33436
rect 15252 33396 15258 33408
rect 15565 33405 15577 33408
rect 15611 33436 15623 33439
rect 16945 33439 17003 33445
rect 16945 33436 16957 33439
rect 15611 33408 16957 33436
rect 15611 33405 15623 33408
rect 15565 33399 15623 33405
rect 16945 33405 16957 33408
rect 16991 33405 17003 33439
rect 17328 33436 17356 33476
rect 17494 33464 17500 33476
rect 17552 33464 17558 33516
rect 19426 33464 19432 33516
rect 19484 33504 19490 33516
rect 20441 33507 20499 33513
rect 20441 33504 20453 33507
rect 19484 33476 20453 33504
rect 19484 33464 19490 33476
rect 20441 33473 20453 33476
rect 20487 33473 20499 33507
rect 24670 33504 24676 33516
rect 24631 33476 24676 33504
rect 20441 33467 20499 33473
rect 24670 33464 24676 33476
rect 24728 33464 24734 33516
rect 24762 33464 24768 33516
rect 24820 33504 24826 33516
rect 24857 33507 24915 33513
rect 24857 33504 24869 33507
rect 24820 33476 24869 33504
rect 24820 33464 24826 33476
rect 24857 33473 24869 33476
rect 24903 33473 24915 33507
rect 24857 33467 24915 33473
rect 25038 33464 25044 33516
rect 25096 33504 25102 33516
rect 25700 33513 25728 33612
rect 26234 33600 26240 33612
rect 26292 33600 26298 33652
rect 25866 33572 25872 33584
rect 25827 33544 25872 33572
rect 25866 33532 25872 33544
rect 25924 33532 25930 33584
rect 25961 33575 26019 33581
rect 25961 33541 25973 33575
rect 26007 33572 26019 33575
rect 26142 33572 26148 33584
rect 26007 33544 26148 33572
rect 26007 33541 26019 33544
rect 25961 33535 26019 33541
rect 26142 33532 26148 33544
rect 26200 33532 26206 33584
rect 26878 33572 26884 33584
rect 26252 33544 26884 33572
rect 25685 33507 25743 33513
rect 25096 33476 25189 33504
rect 25096 33464 25102 33476
rect 25685 33473 25697 33507
rect 25731 33473 25743 33507
rect 26053 33507 26111 33513
rect 26053 33504 26065 33507
rect 25685 33467 25743 33473
rect 25792 33476 26065 33504
rect 17402 33436 17408 33448
rect 17328 33408 17408 33436
rect 16945 33399 17003 33405
rect 17402 33396 17408 33408
rect 17460 33436 17466 33448
rect 18322 33436 18328 33448
rect 17460 33408 18328 33436
rect 17460 33396 17466 33408
rect 18322 33396 18328 33408
rect 18380 33396 18386 33448
rect 25056 33436 25084 33464
rect 25792 33436 25820 33476
rect 26053 33473 26065 33476
rect 26099 33504 26111 33507
rect 26252 33504 26280 33544
rect 26878 33532 26884 33544
rect 26936 33532 26942 33584
rect 26099 33476 26280 33504
rect 26099 33473 26111 33476
rect 26053 33467 26111 33473
rect 27982 33464 27988 33516
rect 28040 33504 28046 33516
rect 29089 33507 29147 33513
rect 29089 33504 29101 33507
rect 28040 33476 29101 33504
rect 28040 33464 28046 33476
rect 29089 33473 29101 33476
rect 29135 33473 29147 33507
rect 29089 33467 29147 33473
rect 29825 33507 29883 33513
rect 29825 33473 29837 33507
rect 29871 33473 29883 33507
rect 29825 33467 29883 33473
rect 25056 33408 25820 33436
rect 25958 33396 25964 33448
rect 26016 33436 26022 33448
rect 27154 33436 27160 33448
rect 26016 33408 27160 33436
rect 26016 33396 26022 33408
rect 27154 33396 27160 33408
rect 27212 33396 27218 33448
rect 28258 33396 28264 33448
rect 28316 33436 28322 33448
rect 29840 33436 29868 33467
rect 28316 33408 29868 33436
rect 28316 33396 28322 33408
rect 11606 33368 11612 33380
rect 10612 33340 11612 33368
rect 11606 33328 11612 33340
rect 11664 33328 11670 33380
rect 12618 33368 12624 33380
rect 12579 33340 12624 33368
rect 12618 33328 12624 33340
rect 12676 33328 12682 33380
rect 13817 33371 13875 33377
rect 13817 33337 13829 33371
rect 13863 33368 13875 33371
rect 14734 33368 14740 33380
rect 13863 33340 14740 33368
rect 13863 33337 13875 33340
rect 13817 33331 13875 33337
rect 14734 33328 14740 33340
rect 14792 33328 14798 33380
rect 15010 33368 15016 33380
rect 14971 33340 15016 33368
rect 15010 33328 15016 33340
rect 15068 33328 15074 33380
rect 24670 33328 24676 33380
rect 24728 33368 24734 33380
rect 25866 33368 25872 33380
rect 24728 33340 25872 33368
rect 24728 33328 24734 33340
rect 25866 33328 25872 33340
rect 25924 33328 25930 33380
rect 1397 33303 1455 33309
rect 1397 33269 1409 33303
rect 1443 33300 1455 33303
rect 9766 33300 9772 33312
rect 1443 33272 9772 33300
rect 1443 33269 1455 33272
rect 1397 33263 1455 33269
rect 9766 33260 9772 33272
rect 9824 33260 9830 33312
rect 20622 33300 20628 33312
rect 20583 33272 20628 33300
rect 20622 33260 20628 33272
rect 20680 33260 20686 33312
rect 25225 33303 25283 33309
rect 25225 33269 25237 33303
rect 25271 33300 25283 33303
rect 26326 33300 26332 33312
rect 25271 33272 26332 33300
rect 25271 33269 25283 33272
rect 25225 33263 25283 33269
rect 26326 33260 26332 33272
rect 26384 33260 26390 33312
rect 29270 33300 29276 33312
rect 29231 33272 29276 33300
rect 29270 33260 29276 33272
rect 29328 33260 29334 33312
rect 30009 33303 30067 33309
rect 30009 33269 30021 33303
rect 30055 33300 30067 33303
rect 30834 33300 30840 33312
rect 30055 33272 30840 33300
rect 30055 33269 30067 33272
rect 30009 33263 30067 33269
rect 30834 33260 30840 33272
rect 30892 33260 30898 33312
rect 1104 33210 30820 33232
rect 1104 33158 5915 33210
rect 5967 33158 5979 33210
rect 6031 33158 6043 33210
rect 6095 33158 6107 33210
rect 6159 33158 6171 33210
rect 6223 33158 15846 33210
rect 15898 33158 15910 33210
rect 15962 33158 15974 33210
rect 16026 33158 16038 33210
rect 16090 33158 16102 33210
rect 16154 33158 25776 33210
rect 25828 33158 25840 33210
rect 25892 33158 25904 33210
rect 25956 33158 25968 33210
rect 26020 33158 26032 33210
rect 26084 33158 30820 33210
rect 1104 33136 30820 33158
rect 10594 33056 10600 33108
rect 10652 33096 10658 33108
rect 10689 33099 10747 33105
rect 10689 33096 10701 33099
rect 10652 33068 10701 33096
rect 10652 33056 10658 33068
rect 10689 33065 10701 33068
rect 10735 33065 10747 33099
rect 11330 33096 11336 33108
rect 10689 33059 10747 33065
rect 11164 33068 11336 33096
rect 11164 32969 11192 33068
rect 11330 33056 11336 33068
rect 11388 33056 11394 33108
rect 14366 33056 14372 33108
rect 14424 33096 14430 33108
rect 16206 33096 16212 33108
rect 14424 33068 15608 33096
rect 16167 33068 16212 33096
rect 14424 33056 14430 33068
rect 11238 32988 11244 33040
rect 11296 32988 11302 33040
rect 15580 33037 15608 33068
rect 16206 33056 16212 33068
rect 16264 33056 16270 33108
rect 18325 33099 18383 33105
rect 18325 33065 18337 33099
rect 18371 33096 18383 33099
rect 18966 33096 18972 33108
rect 18371 33068 18972 33096
rect 18371 33065 18383 33068
rect 18325 33059 18383 33065
rect 18966 33056 18972 33068
rect 19024 33056 19030 33108
rect 19337 33099 19395 33105
rect 19337 33065 19349 33099
rect 19383 33096 19395 33099
rect 20254 33096 20260 33108
rect 19383 33068 20260 33096
rect 19383 33065 19395 33068
rect 19337 33059 19395 33065
rect 20254 33056 20260 33068
rect 20312 33056 20318 33108
rect 22922 33096 22928 33108
rect 20456 33068 22928 33096
rect 15565 33031 15623 33037
rect 15565 32997 15577 33031
rect 15611 32997 15623 33031
rect 15565 32991 15623 32997
rect 11149 32963 11207 32969
rect 11149 32929 11161 32963
rect 11195 32929 11207 32963
rect 11149 32923 11207 32929
rect 1486 32852 1492 32904
rect 1544 32892 1550 32904
rect 1581 32895 1639 32901
rect 1581 32892 1593 32895
rect 1544 32864 1593 32892
rect 1544 32852 1550 32864
rect 1581 32861 1593 32864
rect 1627 32861 1639 32895
rect 1581 32855 1639 32861
rect 9769 32895 9827 32901
rect 9769 32861 9781 32895
rect 9815 32892 9827 32895
rect 9858 32892 9864 32904
rect 9815 32864 9864 32892
rect 9815 32861 9827 32864
rect 9769 32855 9827 32861
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 11256 32901 11284 32988
rect 15580 32960 15608 32991
rect 16574 32988 16580 33040
rect 16632 33028 16638 33040
rect 16853 33031 16911 33037
rect 16853 33028 16865 33031
rect 16632 33000 16865 33028
rect 16632 32988 16638 33000
rect 16853 32997 16865 33000
rect 16899 32997 16911 33031
rect 20456 33028 20484 33068
rect 22922 33056 22928 33068
rect 22980 33056 22986 33108
rect 16853 32991 16911 32997
rect 17328 33000 20484 33028
rect 17328 32960 17356 33000
rect 20530 32988 20536 33040
rect 20588 32988 20594 33040
rect 25685 33031 25743 33037
rect 25685 32997 25697 33031
rect 25731 33028 25743 33031
rect 25774 33028 25780 33040
rect 25731 33000 25780 33028
rect 25731 32997 25743 33000
rect 25685 32991 25743 32997
rect 25774 32988 25780 33000
rect 25832 32988 25838 33040
rect 15580 32932 17356 32960
rect 17402 32920 17408 32972
rect 17460 32960 17466 32972
rect 19702 32960 19708 32972
rect 17460 32932 17505 32960
rect 19663 32932 19708 32960
rect 17460 32920 17466 32932
rect 19702 32920 19708 32932
rect 19760 32920 19766 32972
rect 20548 32960 20576 32988
rect 21910 32960 21916 32972
rect 20548 32932 20668 32960
rect 11241 32895 11299 32901
rect 11241 32861 11253 32895
rect 11287 32861 11299 32895
rect 11241 32855 11299 32861
rect 11606 32852 11612 32904
rect 11664 32892 11670 32904
rect 13541 32895 13599 32901
rect 13541 32892 13553 32895
rect 11664 32864 13553 32892
rect 11664 32852 11670 32864
rect 13541 32861 13553 32864
rect 13587 32892 13599 32895
rect 13630 32892 13636 32904
rect 13587 32864 13636 32892
rect 13587 32861 13599 32864
rect 13541 32855 13599 32861
rect 13630 32852 13636 32864
rect 13688 32852 13694 32904
rect 14185 32895 14243 32901
rect 14185 32861 14197 32895
rect 14231 32892 14243 32895
rect 14918 32892 14924 32904
rect 14231 32864 14924 32892
rect 14231 32861 14243 32864
rect 14185 32855 14243 32861
rect 14918 32852 14924 32864
rect 14976 32852 14982 32904
rect 17126 32892 17132 32904
rect 17087 32864 17132 32892
rect 17126 32852 17132 32864
rect 17184 32852 17190 32904
rect 18141 32895 18199 32901
rect 18141 32861 18153 32895
rect 18187 32892 18199 32895
rect 19426 32892 19432 32904
rect 18187 32864 19432 32892
rect 18187 32861 18199 32864
rect 18141 32855 18199 32861
rect 19426 32852 19432 32864
rect 19484 32852 19490 32904
rect 20530 32892 20536 32904
rect 20491 32864 20536 32892
rect 20530 32852 20536 32864
rect 20588 32852 20594 32904
rect 20640 32901 20668 32932
rect 21468 32932 21916 32960
rect 20625 32895 20683 32901
rect 20625 32861 20637 32895
rect 20671 32861 20683 32895
rect 21266 32892 21272 32904
rect 21227 32864 21272 32892
rect 20625 32855 20683 32861
rect 21266 32852 21272 32864
rect 21324 32852 21330 32904
rect 21468 32901 21496 32932
rect 21910 32920 21916 32932
rect 21968 32960 21974 32972
rect 21968 32932 22692 32960
rect 21968 32920 21974 32932
rect 21453 32895 21511 32901
rect 21453 32861 21465 32895
rect 21499 32861 21511 32895
rect 21453 32855 21511 32861
rect 21821 32895 21879 32901
rect 21821 32861 21833 32895
rect 21867 32892 21879 32895
rect 22462 32892 22468 32904
rect 21867 32864 22468 32892
rect 21867 32861 21879 32864
rect 21821 32855 21879 32861
rect 22462 32852 22468 32864
rect 22520 32852 22526 32904
rect 22664 32901 22692 32932
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 29788 32932 30972 32960
rect 29788 32920 29794 32932
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32861 22707 32895
rect 22649 32855 22707 32861
rect 22741 32895 22799 32901
rect 22741 32861 22753 32895
rect 22787 32892 22799 32895
rect 22922 32892 22928 32904
rect 22787 32864 22928 32892
rect 22787 32861 22799 32864
rect 22741 32855 22799 32861
rect 22922 32852 22928 32864
rect 22980 32852 22986 32904
rect 23934 32852 23940 32904
rect 23992 32892 23998 32904
rect 25133 32895 25191 32901
rect 25133 32892 25145 32895
rect 23992 32864 25145 32892
rect 23992 32852 23998 32864
rect 25133 32861 25145 32864
rect 25179 32861 25191 32895
rect 25133 32855 25191 32861
rect 25501 32895 25559 32901
rect 25501 32861 25513 32895
rect 25547 32892 25559 32895
rect 25866 32892 25872 32904
rect 25547 32864 25872 32892
rect 25547 32861 25559 32864
rect 25501 32855 25559 32861
rect 25866 32852 25872 32864
rect 25924 32892 25930 32904
rect 26878 32892 26884 32904
rect 25924 32864 26884 32892
rect 25924 32852 25930 32864
rect 26878 32852 26884 32864
rect 26936 32852 26942 32904
rect 28718 32892 28724 32904
rect 28679 32864 28724 32892
rect 28718 32852 28724 32864
rect 28776 32852 28782 32904
rect 29825 32895 29883 32901
rect 29825 32861 29837 32895
rect 29871 32892 29883 32895
rect 29871 32864 30880 32892
rect 29871 32861 29883 32864
rect 29825 32855 29883 32861
rect 9585 32827 9643 32833
rect 9585 32793 9597 32827
rect 9631 32824 9643 32827
rect 9674 32824 9680 32836
rect 9631 32796 9680 32824
rect 9631 32793 9643 32796
rect 9585 32787 9643 32793
rect 9674 32784 9680 32796
rect 9732 32784 9738 32836
rect 9953 32827 10011 32833
rect 9953 32793 9965 32827
rect 9999 32824 10011 32827
rect 11793 32827 11851 32833
rect 9999 32796 11652 32824
rect 9999 32793 10011 32796
rect 9953 32787 10011 32793
rect 1397 32759 1455 32765
rect 1397 32725 1409 32759
rect 1443 32756 1455 32759
rect 2590 32756 2596 32768
rect 1443 32728 2596 32756
rect 1443 32725 1455 32728
rect 1397 32719 1455 32725
rect 2590 32716 2596 32728
rect 2648 32716 2654 32768
rect 11149 32759 11207 32765
rect 11149 32725 11161 32759
rect 11195 32756 11207 32759
rect 11514 32756 11520 32768
rect 11195 32728 11520 32756
rect 11195 32725 11207 32728
rect 11149 32719 11207 32725
rect 11514 32716 11520 32728
rect 11572 32716 11578 32768
rect 11624 32756 11652 32796
rect 11793 32793 11805 32827
rect 11839 32824 11851 32827
rect 14274 32824 14280 32836
rect 11839 32796 14280 32824
rect 11839 32793 11851 32796
rect 11793 32787 11851 32793
rect 14274 32784 14280 32796
rect 14332 32784 14338 32836
rect 14458 32833 14464 32836
rect 14452 32787 14464 32833
rect 14516 32824 14522 32836
rect 16117 32827 16175 32833
rect 14516 32796 14552 32824
rect 14458 32784 14464 32787
rect 14516 32784 14522 32796
rect 16117 32793 16129 32827
rect 16163 32824 16175 32827
rect 17034 32824 17040 32836
rect 16163 32796 17040 32824
rect 16163 32793 16175 32796
rect 16117 32787 16175 32793
rect 17034 32784 17040 32796
rect 17092 32784 17098 32836
rect 19058 32784 19064 32836
rect 19116 32824 19122 32836
rect 19797 32827 19855 32833
rect 19797 32824 19809 32827
rect 19116 32796 19809 32824
rect 19116 32784 19122 32796
rect 19797 32793 19809 32796
rect 19843 32793 19855 32827
rect 19797 32787 19855 32793
rect 19889 32827 19947 32833
rect 19889 32793 19901 32827
rect 19935 32824 19947 32827
rect 24026 32824 24032 32836
rect 19935 32796 24032 32824
rect 19935 32793 19947 32796
rect 19889 32787 19947 32793
rect 24026 32784 24032 32796
rect 24084 32784 24090 32836
rect 24946 32784 24952 32836
rect 25004 32824 25010 32836
rect 25317 32827 25375 32833
rect 25317 32824 25329 32827
rect 25004 32796 25329 32824
rect 25004 32784 25010 32796
rect 25317 32793 25329 32796
rect 25363 32793 25375 32827
rect 25317 32787 25375 32793
rect 25409 32827 25467 32833
rect 25409 32793 25421 32827
rect 25455 32793 25467 32827
rect 25409 32787 25467 32793
rect 14734 32756 14740 32768
rect 11624 32728 14740 32756
rect 14734 32716 14740 32728
rect 14792 32716 14798 32768
rect 17313 32759 17371 32765
rect 17313 32725 17325 32759
rect 17359 32756 17371 32759
rect 18046 32756 18052 32768
rect 17359 32728 18052 32756
rect 17359 32725 17371 32728
rect 17313 32719 17371 32725
rect 18046 32716 18052 32728
rect 18104 32716 18110 32768
rect 20714 32716 20720 32768
rect 20772 32756 20778 32768
rect 20809 32759 20867 32765
rect 20809 32756 20821 32759
rect 20772 32728 20821 32756
rect 20772 32716 20778 32728
rect 20809 32725 20821 32728
rect 20855 32725 20867 32759
rect 20809 32719 20867 32725
rect 21729 32759 21787 32765
rect 21729 32725 21741 32759
rect 21775 32756 21787 32759
rect 22002 32756 22008 32768
rect 21775 32728 22008 32756
rect 21775 32725 21787 32728
rect 21729 32719 21787 32725
rect 22002 32716 22008 32728
rect 22060 32716 22066 32768
rect 22281 32759 22339 32765
rect 22281 32725 22293 32759
rect 22327 32756 22339 32759
rect 23290 32756 23296 32768
rect 22327 32728 23296 32756
rect 22327 32725 22339 32728
rect 22281 32719 22339 32725
rect 23290 32716 23296 32728
rect 23348 32716 23354 32768
rect 25038 32716 25044 32768
rect 25096 32756 25102 32768
rect 25424 32756 25452 32787
rect 29730 32784 29736 32836
rect 29788 32824 29794 32836
rect 30558 32824 30564 32836
rect 29788 32796 30564 32824
rect 29788 32784 29794 32796
rect 30558 32784 30564 32796
rect 30616 32784 30622 32836
rect 25096 32728 25452 32756
rect 25096 32716 25102 32728
rect 25590 32716 25596 32768
rect 25648 32756 25654 32768
rect 27982 32756 27988 32768
rect 25648 32728 27988 32756
rect 25648 32716 25654 32728
rect 27982 32716 27988 32728
rect 28040 32716 28046 32768
rect 28442 32716 28448 32768
rect 28500 32756 28506 32768
rect 28626 32756 28632 32768
rect 28500 32728 28632 32756
rect 28500 32716 28506 32728
rect 28626 32716 28632 32728
rect 28684 32716 28690 32768
rect 28902 32756 28908 32768
rect 28863 32728 28908 32756
rect 28902 32716 28908 32728
rect 28960 32716 28966 32768
rect 30009 32759 30067 32765
rect 30009 32725 30021 32759
rect 30055 32756 30067 32759
rect 30190 32756 30196 32768
rect 30055 32728 30196 32756
rect 30055 32725 30067 32728
rect 30009 32719 30067 32725
rect 30190 32716 30196 32728
rect 30248 32716 30254 32768
rect 1104 32666 30820 32688
rect 1104 32614 10880 32666
rect 10932 32614 10944 32666
rect 10996 32614 11008 32666
rect 11060 32614 11072 32666
rect 11124 32614 11136 32666
rect 11188 32614 20811 32666
rect 20863 32614 20875 32666
rect 20927 32614 20939 32666
rect 20991 32614 21003 32666
rect 21055 32614 21067 32666
rect 21119 32614 30820 32666
rect 1104 32592 30820 32614
rect 9953 32555 10011 32561
rect 9953 32521 9965 32555
rect 9999 32552 10011 32555
rect 10410 32552 10416 32564
rect 9999 32524 10416 32552
rect 9999 32521 10011 32524
rect 9953 32515 10011 32521
rect 10410 32512 10416 32524
rect 10468 32512 10474 32564
rect 13170 32552 13176 32564
rect 13131 32524 13176 32552
rect 13170 32512 13176 32524
rect 13228 32512 13234 32564
rect 14093 32555 14151 32561
rect 14093 32521 14105 32555
rect 14139 32552 14151 32555
rect 14458 32552 14464 32564
rect 14139 32524 14464 32552
rect 14139 32521 14151 32524
rect 14093 32515 14151 32521
rect 14458 32512 14464 32524
rect 14516 32512 14522 32564
rect 17221 32555 17279 32561
rect 17221 32521 17233 32555
rect 17267 32552 17279 32555
rect 18046 32552 18052 32564
rect 17267 32524 18052 32552
rect 17267 32521 17279 32524
rect 17221 32515 17279 32521
rect 18046 32512 18052 32524
rect 18104 32512 18110 32564
rect 18690 32512 18696 32564
rect 18748 32552 18754 32564
rect 18969 32555 19027 32561
rect 18969 32552 18981 32555
rect 18748 32524 18981 32552
rect 18748 32512 18754 32524
rect 18969 32521 18981 32524
rect 19015 32552 19027 32555
rect 19058 32552 19064 32564
rect 19015 32524 19064 32552
rect 19015 32521 19027 32524
rect 18969 32515 19027 32521
rect 19058 32512 19064 32524
rect 19116 32512 19122 32564
rect 20530 32512 20536 32564
rect 20588 32552 20594 32564
rect 21821 32555 21879 32561
rect 21821 32552 21833 32555
rect 20588 32524 21833 32552
rect 20588 32512 20594 32524
rect 21821 32521 21833 32524
rect 21867 32521 21879 32555
rect 21821 32515 21879 32521
rect 23658 32512 23664 32564
rect 23716 32552 23722 32564
rect 30852 32552 30880 32864
rect 23716 32524 28212 32552
rect 23716 32512 23722 32524
rect 9766 32484 9772 32496
rect 9727 32456 9772 32484
rect 9766 32444 9772 32456
rect 9824 32444 9830 32496
rect 11146 32444 11152 32496
rect 11204 32484 11210 32496
rect 11514 32484 11520 32496
rect 11204 32456 11520 32484
rect 11204 32444 11210 32456
rect 11514 32444 11520 32456
rect 11572 32444 11578 32496
rect 11790 32444 11796 32496
rect 11848 32484 11854 32496
rect 11885 32487 11943 32493
rect 11885 32484 11897 32487
rect 11848 32456 11897 32484
rect 11848 32444 11854 32456
rect 11885 32453 11897 32456
rect 11931 32453 11943 32487
rect 11885 32447 11943 32453
rect 13630 32444 13636 32496
rect 13688 32484 13694 32496
rect 15289 32487 15347 32493
rect 15289 32484 15301 32487
rect 13688 32456 15301 32484
rect 13688 32444 13694 32456
rect 15289 32453 15301 32456
rect 15335 32453 15347 32487
rect 15289 32447 15347 32453
rect 17037 32487 17095 32493
rect 17037 32453 17049 32487
rect 17083 32484 17095 32487
rect 17126 32484 17132 32496
rect 17083 32456 17132 32484
rect 17083 32453 17095 32456
rect 17037 32447 17095 32453
rect 17126 32444 17132 32456
rect 17184 32444 17190 32496
rect 17313 32487 17371 32493
rect 17313 32453 17325 32487
rect 17359 32484 17371 32487
rect 17402 32484 17408 32496
rect 17359 32456 17408 32484
rect 17359 32453 17371 32456
rect 17313 32447 17371 32453
rect 17402 32444 17408 32456
rect 17460 32444 17466 32496
rect 20162 32484 20168 32496
rect 19628 32456 20168 32484
rect 1578 32416 1584 32428
rect 1539 32388 1584 32416
rect 1578 32376 1584 32388
rect 1636 32376 1642 32428
rect 9585 32419 9643 32425
rect 9585 32385 9597 32419
rect 9631 32416 9643 32419
rect 9674 32416 9680 32428
rect 9631 32388 9680 32416
rect 9631 32385 9643 32388
rect 9585 32379 9643 32385
rect 9674 32376 9680 32388
rect 9732 32376 9738 32428
rect 14366 32416 14372 32428
rect 14327 32388 14372 32416
rect 14366 32376 14372 32388
rect 14424 32376 14430 32428
rect 14458 32419 14516 32425
rect 14458 32412 14470 32419
rect 14504 32412 14516 32419
rect 14458 32360 14464 32412
rect 14516 32360 14522 32412
rect 14550 32376 14556 32428
rect 14608 32425 14614 32428
rect 14608 32416 14616 32425
rect 14608 32388 14653 32416
rect 14608 32379 14616 32388
rect 14608 32376 14614 32379
rect 14734 32376 14740 32428
rect 14792 32416 14798 32428
rect 14792 32388 14837 32416
rect 14792 32376 14798 32388
rect 15102 32376 15108 32428
rect 15160 32416 15166 32428
rect 15933 32419 15991 32425
rect 15933 32416 15945 32419
rect 15160 32388 15945 32416
rect 15160 32376 15166 32388
rect 15933 32385 15945 32388
rect 15979 32385 15991 32419
rect 18782 32416 18788 32428
rect 18743 32388 18788 32416
rect 15933 32379 15991 32385
rect 18782 32376 18788 32388
rect 18840 32376 18846 32428
rect 19628 32425 19656 32456
rect 20162 32444 20168 32456
rect 20220 32444 20226 32496
rect 22186 32484 22192 32496
rect 22147 32456 22192 32484
rect 22186 32444 22192 32456
rect 22244 32444 22250 32496
rect 22327 32487 22385 32493
rect 22327 32453 22339 32487
rect 22373 32484 22385 32487
rect 22462 32484 22468 32496
rect 22373 32456 22468 32484
rect 22373 32453 22385 32456
rect 22327 32447 22385 32453
rect 22462 32444 22468 32456
rect 22520 32444 22526 32496
rect 28184 32493 28212 32524
rect 29472 32524 30880 32552
rect 28169 32487 28227 32493
rect 28169 32453 28181 32487
rect 28215 32484 28227 32487
rect 29089 32487 29147 32493
rect 28215 32456 28580 32484
rect 28215 32453 28227 32456
rect 28169 32447 28227 32453
rect 19886 32425 19892 32428
rect 19613 32419 19671 32425
rect 19613 32385 19625 32419
rect 19659 32385 19671 32419
rect 19613 32379 19671 32385
rect 19880 32379 19892 32425
rect 19944 32416 19950 32428
rect 19944 32388 19980 32416
rect 19886 32376 19892 32379
rect 19944 32376 19950 32388
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 21876 32388 22017 32416
rect 21876 32376 21882 32388
rect 22005 32385 22017 32388
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 22094 32376 22100 32428
rect 22152 32416 22158 32428
rect 22152 32388 22197 32416
rect 22152 32376 22158 32388
rect 22738 32376 22744 32428
rect 22796 32416 22802 32428
rect 23385 32419 23443 32425
rect 23385 32416 23397 32419
rect 22796 32388 23397 32416
rect 22796 32376 22802 32388
rect 23385 32385 23397 32388
rect 23431 32416 23443 32419
rect 23753 32419 23811 32425
rect 23431 32388 23704 32416
rect 23431 32385 23443 32388
rect 23385 32379 23443 32385
rect 18322 32308 18328 32360
rect 18380 32348 18386 32360
rect 18598 32348 18604 32360
rect 18380 32320 18604 32348
rect 18380 32308 18386 32320
rect 18598 32308 18604 32320
rect 18656 32348 18662 32360
rect 19061 32351 19119 32357
rect 19061 32348 19073 32351
rect 18656 32320 19073 32348
rect 18656 32308 18662 32320
rect 19061 32317 19073 32320
rect 19107 32317 19119 32351
rect 22370 32348 22376 32360
rect 19061 32311 19119 32317
rect 21008 32320 22376 32348
rect 11054 32240 11060 32292
rect 11112 32280 11118 32292
rect 11238 32280 11244 32292
rect 11112 32252 11244 32280
rect 11112 32240 11118 32252
rect 11238 32240 11244 32252
rect 11296 32240 11302 32292
rect 21008 32289 21036 32320
rect 22370 32308 22376 32320
rect 22428 32348 22434 32360
rect 22465 32351 22523 32357
rect 22465 32348 22477 32351
rect 22428 32320 22477 32348
rect 22428 32308 22434 32320
rect 22465 32317 22477 32320
rect 22511 32317 22523 32351
rect 22465 32311 22523 32317
rect 20993 32283 21051 32289
rect 20993 32249 21005 32283
rect 21039 32249 21051 32283
rect 20993 32243 21051 32249
rect 22738 32240 22744 32292
rect 22796 32280 22802 32292
rect 23014 32280 23020 32292
rect 22796 32252 23020 32280
rect 22796 32240 22802 32252
rect 23014 32240 23020 32252
rect 23072 32240 23078 32292
rect 1397 32215 1455 32221
rect 1397 32181 1409 32215
rect 1443 32212 1455 32215
rect 2314 32212 2320 32224
rect 1443 32184 2320 32212
rect 1443 32181 1455 32184
rect 1397 32175 1455 32181
rect 2314 32172 2320 32184
rect 2372 32172 2378 32224
rect 12342 32172 12348 32224
rect 12400 32212 12406 32224
rect 15381 32215 15439 32221
rect 15381 32212 15393 32215
rect 12400 32184 15393 32212
rect 12400 32172 12406 32184
rect 15381 32181 15393 32184
rect 15427 32181 15439 32215
rect 15381 32175 15439 32181
rect 15746 32172 15752 32224
rect 15804 32212 15810 32224
rect 16117 32215 16175 32221
rect 16117 32212 16129 32215
rect 15804 32184 16129 32212
rect 15804 32172 15810 32184
rect 16117 32181 16129 32184
rect 16163 32181 16175 32215
rect 16117 32175 16175 32181
rect 16298 32172 16304 32224
rect 16356 32212 16362 32224
rect 16761 32215 16819 32221
rect 16761 32212 16773 32215
rect 16356 32184 16773 32212
rect 16356 32172 16362 32184
rect 16761 32181 16773 32184
rect 16807 32181 16819 32215
rect 16761 32175 16819 32181
rect 18414 32172 18420 32224
rect 18472 32212 18478 32224
rect 18509 32215 18567 32221
rect 18509 32212 18521 32215
rect 18472 32184 18521 32212
rect 18472 32172 18478 32184
rect 18509 32181 18521 32184
rect 18555 32181 18567 32215
rect 23676 32212 23704 32388
rect 23753 32385 23765 32419
rect 23799 32416 23811 32419
rect 24026 32416 24032 32428
rect 23799 32388 24032 32416
rect 23799 32385 23811 32388
rect 23753 32379 23811 32385
rect 24026 32376 24032 32388
rect 24084 32416 24090 32428
rect 25593 32419 25651 32425
rect 24084 32388 24532 32416
rect 24084 32376 24090 32388
rect 24504 32280 24532 32388
rect 25593 32385 25605 32419
rect 25639 32416 25651 32419
rect 26326 32416 26332 32428
rect 25639 32388 26332 32416
rect 25639 32385 25651 32388
rect 25593 32379 25651 32385
rect 26326 32376 26332 32388
rect 26384 32376 26390 32428
rect 27985 32419 28043 32425
rect 27985 32385 27997 32419
rect 28031 32385 28043 32419
rect 27985 32379 28043 32385
rect 25866 32348 25872 32360
rect 25827 32320 25872 32348
rect 25866 32308 25872 32320
rect 25924 32308 25930 32360
rect 28000 32348 28028 32379
rect 28074 32376 28080 32428
rect 28132 32416 28138 32428
rect 28245 32419 28303 32425
rect 28245 32416 28257 32419
rect 28132 32388 28257 32416
rect 28132 32376 28138 32388
rect 28245 32385 28257 32388
rect 28291 32385 28303 32419
rect 28245 32379 28303 32385
rect 28000 32320 28212 32348
rect 28184 32292 28212 32320
rect 24504 32252 27752 32280
rect 27724 32224 27752 32252
rect 28166 32240 28172 32292
rect 28224 32240 28230 32292
rect 28552 32280 28580 32456
rect 29089 32453 29101 32487
rect 29135 32484 29147 32487
rect 29472 32484 29500 32524
rect 30944 32484 30972 32932
rect 29135 32456 29500 32484
rect 30852 32456 30972 32484
rect 29135 32453 29147 32456
rect 29089 32447 29147 32453
rect 28718 32416 28724 32428
rect 28679 32388 28724 32416
rect 28718 32376 28724 32388
rect 28776 32376 28782 32428
rect 28994 32376 29000 32428
rect 29052 32416 29058 32428
rect 29365 32419 29423 32425
rect 29365 32416 29377 32419
rect 29052 32388 29377 32416
rect 29052 32376 29058 32388
rect 29365 32385 29377 32388
rect 29411 32385 29423 32419
rect 29365 32379 29423 32385
rect 29457 32419 29515 32425
rect 29457 32385 29469 32419
rect 29503 32385 29515 32419
rect 29457 32379 29515 32385
rect 29549 32419 29607 32425
rect 29549 32385 29561 32419
rect 29595 32385 29607 32419
rect 29549 32379 29607 32385
rect 29733 32419 29791 32425
rect 29733 32385 29745 32419
rect 29779 32416 29868 32419
rect 29779 32391 30052 32416
rect 29779 32385 29791 32391
rect 29840 32388 30052 32391
rect 29733 32379 29791 32385
rect 28736 32348 28764 32376
rect 29472 32348 29500 32379
rect 28736 32320 29500 32348
rect 29564 32348 29592 32379
rect 29822 32348 29828 32360
rect 29564 32320 29828 32348
rect 29822 32308 29828 32320
rect 29880 32308 29886 32360
rect 29362 32280 29368 32292
rect 28552 32252 29368 32280
rect 29362 32240 29368 32252
rect 29420 32240 29426 32292
rect 26234 32212 26240 32224
rect 23676 32184 26240 32212
rect 18509 32175 18567 32181
rect 26234 32172 26240 32184
rect 26292 32172 26298 32224
rect 27706 32172 27712 32224
rect 27764 32172 27770 32224
rect 27801 32215 27859 32221
rect 27801 32181 27813 32215
rect 27847 32212 27859 32215
rect 30024 32212 30052 32388
rect 27847 32184 30052 32212
rect 27847 32181 27859 32184
rect 27801 32175 27859 32181
rect 1104 32122 30820 32144
rect 1104 32070 5915 32122
rect 5967 32070 5979 32122
rect 6031 32070 6043 32122
rect 6095 32070 6107 32122
rect 6159 32070 6171 32122
rect 6223 32070 15846 32122
rect 15898 32070 15910 32122
rect 15962 32070 15974 32122
rect 16026 32070 16038 32122
rect 16090 32070 16102 32122
rect 16154 32070 25776 32122
rect 25828 32070 25840 32122
rect 25892 32070 25904 32122
rect 25956 32070 25968 32122
rect 26020 32070 26032 32122
rect 26084 32070 30820 32122
rect 1104 32048 30820 32070
rect 2777 32011 2835 32017
rect 2777 31977 2789 32011
rect 2823 32008 2835 32011
rect 2823 31980 11376 32008
rect 2823 31977 2835 31980
rect 2777 31971 2835 31977
rect 9493 31943 9551 31949
rect 9493 31909 9505 31943
rect 9539 31940 9551 31943
rect 9674 31940 9680 31952
rect 9539 31912 9680 31940
rect 9539 31909 9551 31912
rect 9493 31903 9551 31909
rect 9674 31900 9680 31912
rect 9732 31900 9738 31952
rect 10413 31943 10471 31949
rect 10413 31909 10425 31943
rect 10459 31940 10471 31943
rect 11238 31940 11244 31952
rect 10459 31912 11244 31940
rect 10459 31909 10471 31912
rect 10413 31903 10471 31909
rect 11238 31900 11244 31912
rect 11296 31900 11302 31952
rect 11348 31940 11376 31980
rect 11422 31968 11428 32020
rect 11480 32008 11486 32020
rect 11609 32011 11667 32017
rect 11609 32008 11621 32011
rect 11480 31980 11621 32008
rect 11480 31968 11486 31980
rect 11609 31977 11621 31980
rect 11655 31977 11667 32011
rect 11609 31971 11667 31977
rect 13078 31968 13084 32020
rect 13136 32008 13142 32020
rect 13357 32011 13415 32017
rect 13357 32008 13369 32011
rect 13136 31980 13369 32008
rect 13136 31968 13142 31980
rect 13357 31977 13369 31980
rect 13403 31977 13415 32011
rect 14274 32008 14280 32020
rect 14235 31980 14280 32008
rect 13357 31971 13415 31977
rect 14274 31968 14280 31980
rect 14332 31968 14338 32020
rect 15562 31968 15568 32020
rect 15620 32008 15626 32020
rect 16301 32011 16359 32017
rect 16301 32008 16313 32011
rect 15620 31980 16313 32008
rect 15620 31968 15626 31980
rect 15948 31952 15976 31980
rect 16301 31977 16313 31980
rect 16347 31977 16359 32011
rect 16301 31971 16359 31977
rect 19886 31968 19892 32020
rect 19944 32008 19950 32020
rect 20073 32011 20131 32017
rect 20073 32008 20085 32011
rect 19944 31980 20085 32008
rect 19944 31968 19950 31980
rect 20073 31977 20085 31980
rect 20119 31977 20131 32011
rect 20073 31971 20131 31977
rect 21453 32011 21511 32017
rect 21453 31977 21465 32011
rect 21499 32008 21511 32011
rect 22186 32008 22192 32020
rect 21499 31980 22192 32008
rect 21499 31977 21511 31980
rect 21453 31971 21511 31977
rect 22186 31968 22192 31980
rect 22244 31968 22250 32020
rect 22646 32008 22652 32020
rect 22388 31980 22652 32008
rect 11348 31912 13952 31940
rect 10873 31875 10931 31881
rect 10873 31841 10885 31875
rect 10919 31872 10931 31875
rect 11330 31872 11336 31884
rect 10919 31844 11336 31872
rect 10919 31841 10931 31844
rect 10873 31835 10931 31841
rect 11330 31832 11336 31844
rect 11388 31872 11394 31884
rect 11977 31875 12035 31881
rect 11977 31872 11989 31875
rect 11388 31844 11989 31872
rect 11388 31832 11394 31844
rect 11977 31841 11989 31844
rect 12023 31872 12035 31875
rect 12066 31872 12072 31884
rect 12023 31844 12072 31872
rect 12023 31841 12035 31844
rect 11977 31835 12035 31841
rect 12066 31832 12072 31844
rect 12124 31832 12130 31884
rect 13814 31872 13820 31884
rect 13280 31844 13820 31872
rect 1854 31804 1860 31816
rect 1815 31776 1860 31804
rect 1854 31764 1860 31776
rect 1912 31764 1918 31816
rect 2409 31807 2467 31813
rect 2409 31773 2421 31807
rect 2455 31804 2467 31807
rect 2498 31804 2504 31816
rect 2455 31776 2504 31804
rect 2455 31773 2467 31776
rect 2409 31767 2467 31773
rect 2498 31764 2504 31776
rect 2556 31764 2562 31816
rect 2590 31764 2596 31816
rect 2648 31804 2654 31816
rect 9677 31807 9735 31813
rect 2648 31776 2693 31804
rect 2648 31764 2654 31776
rect 9677 31773 9689 31807
rect 9723 31804 9735 31807
rect 9766 31804 9772 31816
rect 9723 31776 9772 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 9766 31764 9772 31776
rect 9824 31804 9830 31816
rect 10042 31804 10048 31816
rect 9824 31776 10048 31804
rect 9824 31764 9830 31776
rect 10042 31764 10048 31776
rect 10100 31764 10106 31816
rect 10965 31807 11023 31813
rect 10965 31773 10977 31807
rect 11011 31804 11023 31807
rect 11054 31804 11060 31816
rect 11011 31776 11060 31804
rect 11011 31773 11023 31776
rect 10965 31767 11023 31773
rect 11054 31764 11060 31776
rect 11112 31804 11118 31816
rect 13280 31813 13308 31844
rect 13814 31832 13820 31844
rect 13872 31832 13878 31884
rect 12161 31807 12219 31813
rect 12161 31804 12173 31807
rect 11112 31776 12173 31804
rect 11112 31764 11118 31776
rect 12161 31773 12173 31776
rect 12207 31773 12219 31807
rect 12161 31767 12219 31773
rect 13265 31807 13323 31813
rect 13265 31773 13277 31807
rect 13311 31773 13323 31807
rect 13265 31767 13323 31773
rect 11146 31696 11152 31748
rect 11204 31696 11210 31748
rect 13924 31736 13952 31912
rect 15930 31900 15936 31952
rect 15988 31900 15994 31952
rect 17865 31943 17923 31949
rect 17865 31909 17877 31943
rect 17911 31940 17923 31943
rect 18966 31940 18972 31952
rect 17911 31912 18972 31940
rect 17911 31909 17923 31912
rect 17865 31903 17923 31909
rect 18966 31900 18972 31912
rect 19024 31900 19030 31952
rect 21910 31900 21916 31952
rect 21968 31940 21974 31952
rect 22094 31940 22100 31952
rect 21968 31912 22100 31940
rect 21968 31900 21974 31912
rect 22094 31900 22100 31912
rect 22152 31940 22158 31952
rect 22388 31940 22416 31980
rect 22646 31968 22652 31980
rect 22704 31968 22710 32020
rect 23198 31968 23204 32020
rect 23256 32008 23262 32020
rect 23256 31980 23428 32008
rect 23256 31968 23262 31980
rect 22152 31912 22416 31940
rect 23400 31940 23428 31980
rect 23566 31968 23572 32020
rect 23624 32008 23630 32020
rect 24026 32008 24032 32020
rect 23624 31980 24032 32008
rect 23624 31968 23630 31980
rect 24026 31968 24032 31980
rect 24084 31968 24090 32020
rect 24397 32011 24455 32017
rect 24397 31977 24409 32011
rect 24443 32008 24455 32011
rect 24670 32008 24676 32020
rect 24443 31980 24676 32008
rect 24443 31977 24455 31980
rect 24397 31971 24455 31977
rect 24670 31968 24676 31980
rect 24728 31968 24734 32020
rect 26881 32011 26939 32017
rect 26881 32008 26893 32011
rect 24780 31980 26893 32008
rect 24780 31940 24808 31980
rect 26881 31977 26893 31980
rect 26927 31977 26939 32011
rect 28077 32011 28135 32017
rect 28077 32008 28089 32011
rect 26881 31971 26939 31977
rect 26988 31980 28089 32008
rect 23400 31912 24808 31940
rect 22152 31900 22158 31912
rect 26050 31900 26056 31952
rect 26108 31940 26114 31952
rect 26988 31940 27016 31980
rect 28077 31977 28089 31980
rect 28123 31977 28135 32011
rect 28077 31971 28135 31977
rect 28442 31968 28448 32020
rect 28500 32008 28506 32020
rect 30101 32011 30159 32017
rect 30101 32008 30113 32011
rect 28500 31980 30113 32008
rect 28500 31968 28506 31980
rect 30101 31977 30113 31980
rect 30147 31977 30159 32011
rect 30101 31971 30159 31977
rect 30374 31968 30380 32020
rect 30432 32008 30438 32020
rect 30432 31980 30512 32008
rect 30432 31968 30438 31980
rect 26108 31912 27016 31940
rect 26108 31900 26114 31912
rect 28258 31900 28264 31952
rect 28316 31940 28322 31952
rect 29730 31940 29736 31952
rect 28316 31912 29736 31940
rect 28316 31900 28322 31912
rect 29730 31900 29736 31912
rect 29788 31900 29794 31952
rect 18138 31832 18144 31884
rect 18196 31872 18202 31884
rect 18325 31875 18383 31881
rect 18325 31872 18337 31875
rect 18196 31844 18337 31872
rect 18196 31832 18202 31844
rect 18325 31841 18337 31844
rect 18371 31872 18383 31875
rect 18782 31872 18788 31884
rect 18371 31844 18788 31872
rect 18371 31841 18383 31844
rect 18325 31835 18383 31841
rect 18782 31832 18788 31844
rect 18840 31832 18846 31884
rect 19978 31832 19984 31884
rect 20036 31872 20042 31884
rect 22462 31872 22468 31884
rect 20036 31844 22468 31872
rect 20036 31832 20042 31844
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 24118 31832 24124 31884
rect 24176 31872 24182 31884
rect 24176 31844 24624 31872
rect 24176 31832 24182 31844
rect 14090 31804 14096 31816
rect 14051 31776 14096 31804
rect 14090 31764 14096 31776
rect 14148 31764 14154 31816
rect 16209 31807 16267 31813
rect 16209 31773 16221 31807
rect 16255 31804 16267 31807
rect 16666 31804 16672 31816
rect 16255 31776 16672 31804
rect 16255 31773 16267 31776
rect 16209 31767 16267 31773
rect 16666 31764 16672 31776
rect 16724 31804 16730 31816
rect 17678 31804 17684 31816
rect 16724 31776 17684 31804
rect 16724 31764 16730 31776
rect 17678 31764 17684 31776
rect 17736 31764 17742 31816
rect 18230 31764 18236 31816
rect 18288 31804 18294 31816
rect 18417 31807 18475 31813
rect 18417 31804 18429 31807
rect 18288 31776 18429 31804
rect 18288 31764 18294 31776
rect 18417 31773 18429 31776
rect 18463 31773 18475 31807
rect 18417 31767 18475 31773
rect 20257 31807 20315 31813
rect 20257 31773 20269 31807
rect 20303 31804 20315 31807
rect 20714 31804 20720 31816
rect 20303 31776 20720 31804
rect 20303 31773 20315 31776
rect 20257 31767 20315 31773
rect 20714 31764 20720 31776
rect 20772 31764 20778 31816
rect 21266 31764 21272 31816
rect 21324 31804 21330 31816
rect 21637 31807 21695 31813
rect 21637 31804 21649 31807
rect 21324 31776 21649 31804
rect 21324 31764 21330 31776
rect 21637 31773 21649 31776
rect 21683 31773 21695 31807
rect 21637 31767 21695 31773
rect 21729 31807 21787 31813
rect 21729 31773 21741 31807
rect 21775 31773 21787 31807
rect 21910 31804 21916 31816
rect 21871 31776 21916 31804
rect 21729 31767 21787 31773
rect 15010 31736 15016 31748
rect 13924 31708 15016 31736
rect 15010 31696 15016 31708
rect 15068 31696 15074 31748
rect 18325 31739 18383 31745
rect 15120 31708 16896 31736
rect 1670 31668 1676 31680
rect 1631 31640 1676 31668
rect 1670 31628 1676 31640
rect 1728 31628 1734 31680
rect 10873 31671 10931 31677
rect 10873 31637 10885 31671
rect 10919 31668 10931 31671
rect 11164 31668 11192 31696
rect 10919 31640 11192 31668
rect 12069 31671 12127 31677
rect 10919 31637 10931 31640
rect 10873 31631 10931 31637
rect 12069 31637 12081 31671
rect 12115 31668 12127 31671
rect 12158 31668 12164 31680
rect 12115 31640 12164 31668
rect 12115 31637 12127 31640
rect 12069 31631 12127 31637
rect 12158 31628 12164 31640
rect 12216 31628 12222 31680
rect 12802 31628 12808 31680
rect 12860 31668 12866 31680
rect 15120 31668 15148 31708
rect 12860 31640 15148 31668
rect 12860 31628 12866 31640
rect 15286 31628 15292 31680
rect 15344 31668 15350 31680
rect 15562 31668 15568 31680
rect 15344 31640 15568 31668
rect 15344 31628 15350 31640
rect 15562 31628 15568 31640
rect 15620 31628 15626 31680
rect 15654 31628 15660 31680
rect 15712 31668 15718 31680
rect 16758 31668 16764 31680
rect 15712 31640 16764 31668
rect 15712 31628 15718 31640
rect 16758 31628 16764 31640
rect 16816 31628 16822 31680
rect 16868 31668 16896 31708
rect 18325 31705 18337 31739
rect 18371 31736 18383 31739
rect 18690 31736 18696 31748
rect 18371 31708 18696 31736
rect 18371 31705 18383 31708
rect 18325 31699 18383 31705
rect 18690 31696 18696 31708
rect 18748 31696 18754 31748
rect 21744 31736 21772 31767
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 22005 31807 22063 31813
rect 22005 31773 22017 31807
rect 22051 31804 22063 31807
rect 22094 31804 22100 31816
rect 22051 31776 22100 31804
rect 22051 31773 22063 31776
rect 22005 31767 22063 31773
rect 22094 31764 22100 31776
rect 22152 31764 22158 31816
rect 24596 31813 24624 31844
rect 25406 31832 25412 31884
rect 25464 31872 25470 31884
rect 25590 31872 25596 31884
rect 25464 31844 25596 31872
rect 25464 31832 25470 31844
rect 25590 31832 25596 31844
rect 25648 31832 25654 31884
rect 27246 31872 27252 31884
rect 27207 31844 27252 31872
rect 27246 31832 27252 31844
rect 27304 31832 27310 31884
rect 27706 31832 27712 31884
rect 27764 31872 27770 31884
rect 28074 31872 28080 31884
rect 27764 31844 28080 31872
rect 27764 31832 27770 31844
rect 28074 31832 28080 31844
rect 28132 31832 28138 31884
rect 28537 31875 28595 31881
rect 28537 31841 28549 31875
rect 28583 31872 28595 31875
rect 28718 31872 28724 31884
rect 28583 31844 28724 31872
rect 28583 31841 28595 31844
rect 28537 31835 28595 31841
rect 28718 31832 28724 31844
rect 28776 31832 28782 31884
rect 30374 31872 30380 31884
rect 29748 31844 30380 31872
rect 24581 31807 24639 31813
rect 22204 31776 23520 31804
rect 22204 31736 22232 31776
rect 21744 31708 22232 31736
rect 22732 31739 22790 31745
rect 22732 31705 22744 31739
rect 22778 31736 22790 31739
rect 23106 31736 23112 31748
rect 22778 31708 23112 31736
rect 22778 31705 22790 31708
rect 22732 31699 22790 31705
rect 23106 31696 23112 31708
rect 23164 31696 23170 31748
rect 23492 31736 23520 31776
rect 24581 31773 24593 31807
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 24670 31764 24676 31816
rect 24728 31804 24734 31816
rect 24765 31807 24823 31813
rect 24765 31804 24777 31807
rect 24728 31776 24777 31804
rect 24728 31764 24734 31776
rect 24765 31773 24777 31776
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31773 24915 31807
rect 24857 31767 24915 31773
rect 26145 31807 26203 31813
rect 26145 31773 26157 31807
rect 26191 31804 26203 31807
rect 26234 31804 26240 31816
rect 26191 31776 26240 31804
rect 26191 31773 26203 31776
rect 26145 31767 26203 31773
rect 23566 31736 23572 31748
rect 23479 31708 23572 31736
rect 23566 31696 23572 31708
rect 23624 31736 23630 31748
rect 24872 31736 24900 31767
rect 26234 31764 26240 31776
rect 26292 31764 26298 31816
rect 29748 31813 29776 31844
rect 30374 31832 30380 31844
rect 30432 31832 30438 31884
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31804 26387 31807
rect 27433 31807 27491 31813
rect 26375 31776 27016 31804
rect 26375 31773 26387 31776
rect 26329 31767 26387 31773
rect 23624 31708 24900 31736
rect 26988 31736 27016 31776
rect 27433 31773 27445 31807
rect 27479 31804 27491 31807
rect 29733 31807 29791 31813
rect 27479 31776 28488 31804
rect 27479 31773 27491 31776
rect 27433 31767 27491 31773
rect 27062 31736 27068 31748
rect 26988 31708 27068 31736
rect 23624 31696 23630 31708
rect 23658 31668 23664 31680
rect 16868 31640 23664 31668
rect 23658 31628 23664 31640
rect 23716 31628 23722 31680
rect 23860 31677 23888 31708
rect 27062 31696 27068 31708
rect 27120 31696 27126 31748
rect 27338 31736 27344 31748
rect 27299 31708 27344 31736
rect 27338 31696 27344 31708
rect 27396 31696 27402 31748
rect 28460 31736 28488 31776
rect 29733 31773 29745 31807
rect 29779 31773 29791 31807
rect 29733 31767 29791 31773
rect 30098 31764 30104 31816
rect 30156 31804 30162 31816
rect 30484 31804 30512 31980
rect 30852 31952 30880 32456
rect 30834 31900 30840 31952
rect 30892 31900 30898 31952
rect 30156 31776 30512 31804
rect 30156 31764 30162 31776
rect 28629 31739 28687 31745
rect 28629 31736 28641 31739
rect 28460 31708 28641 31736
rect 28629 31705 28641 31708
rect 28675 31705 28687 31739
rect 29362 31736 29368 31748
rect 28629 31699 28687 31705
rect 28966 31708 29368 31736
rect 23845 31671 23903 31677
rect 23845 31637 23857 31671
rect 23891 31637 23903 31671
rect 23845 31631 23903 31637
rect 26786 31628 26792 31680
rect 26844 31668 26850 31680
rect 28537 31671 28595 31677
rect 28537 31668 28549 31671
rect 26844 31640 28549 31668
rect 26844 31628 26850 31640
rect 28537 31637 28549 31640
rect 28583 31637 28595 31671
rect 28644 31668 28672 31699
rect 28966 31668 28994 31708
rect 29362 31696 29368 31708
rect 29420 31696 29426 31748
rect 29917 31739 29975 31745
rect 29917 31705 29929 31739
rect 29963 31705 29975 31739
rect 29917 31699 29975 31705
rect 28644 31640 28994 31668
rect 29932 31668 29960 31699
rect 30006 31668 30012 31680
rect 29932 31640 30012 31668
rect 28537 31631 28595 31637
rect 30006 31628 30012 31640
rect 30064 31628 30070 31680
rect 30190 31628 30196 31680
rect 30248 31668 30254 31680
rect 30558 31668 30564 31680
rect 30248 31640 30564 31668
rect 30248 31628 30254 31640
rect 30558 31628 30564 31640
rect 30616 31628 30622 31680
rect 1104 31578 30820 31600
rect 1104 31526 10880 31578
rect 10932 31526 10944 31578
rect 10996 31526 11008 31578
rect 11060 31526 11072 31578
rect 11124 31526 11136 31578
rect 11188 31526 20811 31578
rect 20863 31526 20875 31578
rect 20927 31526 20939 31578
rect 20991 31526 21003 31578
rect 21055 31526 21067 31578
rect 21119 31526 30820 31578
rect 1104 31504 30820 31526
rect 4062 31424 4068 31476
rect 4120 31464 4126 31476
rect 4120 31436 10732 31464
rect 4120 31424 4126 31436
rect 2409 31399 2467 31405
rect 2409 31365 2421 31399
rect 2455 31396 2467 31399
rect 2498 31396 2504 31408
rect 2455 31368 2504 31396
rect 2455 31365 2467 31368
rect 2409 31359 2467 31365
rect 2498 31356 2504 31368
rect 2556 31356 2562 31408
rect 3970 31356 3976 31408
rect 4028 31396 4034 31408
rect 10704 31405 10732 31436
rect 12066 31424 12072 31476
rect 12124 31464 12130 31476
rect 12437 31467 12495 31473
rect 12437 31464 12449 31467
rect 12124 31436 12449 31464
rect 12124 31424 12130 31436
rect 12437 31433 12449 31436
rect 12483 31433 12495 31467
rect 13262 31464 13268 31476
rect 13223 31436 13268 31464
rect 12437 31427 12495 31433
rect 13262 31424 13268 31436
rect 13320 31424 13326 31476
rect 13998 31464 14004 31476
rect 13957 31436 14004 31464
rect 13998 31424 14004 31436
rect 14056 31473 14062 31476
rect 14056 31467 14105 31473
rect 14056 31433 14059 31467
rect 14093 31464 14105 31467
rect 14550 31464 14556 31476
rect 14093 31436 14556 31464
rect 14093 31433 14105 31436
rect 14056 31427 14105 31433
rect 14056 31424 14062 31427
rect 14550 31424 14556 31436
rect 14608 31424 14614 31476
rect 15010 31424 15016 31476
rect 15068 31464 15074 31476
rect 17221 31467 17279 31473
rect 15068 31436 16160 31464
rect 15068 31424 15074 31436
rect 9861 31399 9919 31405
rect 9861 31396 9873 31399
rect 4028 31368 9873 31396
rect 4028 31356 4034 31368
rect 9861 31365 9873 31368
rect 9907 31365 9919 31399
rect 9861 31359 9919 31365
rect 10689 31399 10747 31405
rect 10689 31365 10701 31399
rect 10735 31365 10747 31399
rect 10689 31359 10747 31365
rect 12345 31399 12403 31405
rect 12345 31365 12357 31399
rect 12391 31396 12403 31399
rect 13078 31396 13084 31408
rect 12391 31368 13084 31396
rect 12391 31365 12403 31368
rect 12345 31359 12403 31365
rect 13078 31356 13084 31368
rect 13136 31356 13142 31408
rect 15378 31356 15384 31408
rect 15436 31396 15442 31408
rect 15562 31396 15568 31408
rect 15436 31368 15568 31396
rect 15436 31356 15442 31368
rect 15562 31356 15568 31368
rect 15620 31396 15626 31408
rect 15620 31368 15884 31396
rect 15620 31356 15626 31368
rect 1854 31328 1860 31340
rect 1815 31300 1860 31328
rect 1854 31288 1860 31300
rect 1912 31288 1918 31340
rect 2314 31288 2320 31340
rect 2372 31328 2378 31340
rect 2593 31331 2651 31337
rect 2593 31328 2605 31331
rect 2372 31300 2605 31328
rect 2372 31288 2378 31300
rect 2593 31297 2605 31300
rect 2639 31297 2651 31331
rect 9674 31328 9680 31340
rect 9635 31300 9680 31328
rect 2593 31291 2651 31297
rect 9674 31288 9680 31300
rect 9732 31328 9738 31340
rect 10505 31331 10563 31337
rect 10505 31328 10517 31331
rect 9732 31300 10517 31328
rect 9732 31288 9738 31300
rect 10505 31297 10517 31300
rect 10551 31297 10563 31331
rect 10505 31291 10563 31297
rect 13173 31331 13231 31337
rect 13173 31297 13185 31331
rect 13219 31328 13231 31331
rect 15102 31328 15108 31340
rect 13219 31300 15108 31328
rect 13219 31297 13231 31300
rect 13173 31291 13231 31297
rect 15102 31288 15108 31300
rect 15160 31288 15166 31340
rect 15654 31288 15660 31340
rect 15712 31328 15718 31340
rect 15856 31337 15884 31368
rect 15749 31331 15807 31337
rect 15749 31328 15761 31331
rect 15712 31300 15761 31328
rect 15712 31288 15718 31300
rect 15749 31297 15761 31300
rect 15795 31297 15807 31331
rect 15749 31291 15807 31297
rect 15841 31331 15899 31337
rect 15841 31297 15853 31331
rect 15887 31297 15899 31331
rect 15841 31291 15899 31297
rect 15930 31288 15936 31340
rect 15988 31328 15994 31340
rect 16132 31337 16160 31436
rect 17221 31433 17233 31467
rect 17267 31464 17279 31467
rect 17310 31464 17316 31476
rect 17267 31436 17316 31464
rect 17267 31433 17279 31436
rect 17221 31427 17279 31433
rect 17310 31424 17316 31436
rect 17368 31424 17374 31476
rect 21818 31424 21824 31476
rect 21876 31464 21882 31476
rect 22649 31467 22707 31473
rect 22649 31464 22661 31467
rect 21876 31436 22661 31464
rect 21876 31424 21882 31436
rect 22649 31433 22661 31436
rect 22695 31433 22707 31467
rect 23106 31464 23112 31476
rect 23067 31436 23112 31464
rect 22649 31427 22707 31433
rect 23106 31424 23112 31436
rect 23164 31424 23170 31476
rect 24029 31467 24087 31473
rect 24029 31433 24041 31467
rect 24075 31464 24087 31467
rect 24762 31464 24768 31476
rect 24075 31436 24768 31464
rect 24075 31433 24087 31436
rect 24029 31427 24087 31433
rect 24762 31424 24768 31436
rect 24820 31424 24826 31476
rect 24854 31424 24860 31476
rect 24912 31464 24918 31476
rect 24949 31467 25007 31473
rect 24949 31464 24961 31467
rect 24912 31436 24961 31464
rect 24912 31424 24918 31436
rect 24949 31433 24961 31436
rect 24995 31433 25007 31467
rect 26421 31467 26479 31473
rect 24949 31427 25007 31433
rect 25332 31436 26096 31464
rect 19337 31399 19395 31405
rect 19337 31365 19349 31399
rect 19383 31396 19395 31399
rect 19518 31396 19524 31408
rect 19383 31368 19524 31396
rect 19383 31365 19395 31368
rect 19337 31359 19395 31365
rect 19518 31356 19524 31368
rect 19576 31356 19582 31408
rect 22554 31396 22560 31408
rect 22296 31368 22560 31396
rect 16117 31331 16175 31337
rect 15988 31300 16033 31328
rect 15988 31288 15994 31300
rect 16117 31297 16129 31331
rect 16163 31297 16175 31331
rect 16117 31291 16175 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31328 17371 31331
rect 18322 31328 18328 31340
rect 17359 31300 18328 31328
rect 17359 31297 17371 31300
rect 17313 31291 17371 31297
rect 18322 31288 18328 31300
rect 18380 31288 18386 31340
rect 22094 31288 22100 31340
rect 22152 31328 22158 31340
rect 22296 31337 22324 31368
rect 22554 31356 22560 31368
rect 22612 31356 22618 31408
rect 25332 31396 25360 31436
rect 22940 31368 25360 31396
rect 26068 31396 26096 31436
rect 26421 31433 26433 31467
rect 26467 31464 26479 31467
rect 26970 31464 26976 31476
rect 26467 31436 26976 31464
rect 26467 31433 26479 31436
rect 26421 31427 26479 31433
rect 26970 31424 26976 31436
rect 27028 31424 27034 31476
rect 27617 31467 27675 31473
rect 27617 31433 27629 31467
rect 27663 31464 27675 31467
rect 27706 31464 27712 31476
rect 27663 31436 27712 31464
rect 27663 31433 27675 31436
rect 27617 31427 27675 31433
rect 27706 31424 27712 31436
rect 27764 31424 27770 31476
rect 26068 31368 27016 31396
rect 22281 31331 22339 31337
rect 22281 31328 22293 31331
rect 22152 31300 22293 31328
rect 22152 31288 22158 31300
rect 22281 31297 22293 31300
rect 22327 31297 22339 31331
rect 22281 31291 22339 31297
rect 22465 31331 22523 31337
rect 22465 31297 22477 31331
rect 22511 31328 22523 31331
rect 22940 31328 22968 31368
rect 26988 31340 27016 31368
rect 27522 31356 27528 31408
rect 27580 31396 27586 31408
rect 28721 31399 28779 31405
rect 28721 31396 28733 31399
rect 27580 31368 28733 31396
rect 27580 31356 27586 31368
rect 28721 31365 28733 31368
rect 28767 31396 28779 31399
rect 29641 31399 29699 31405
rect 29641 31396 29653 31399
rect 28767 31368 29653 31396
rect 28767 31365 28779 31368
rect 28721 31359 28779 31365
rect 29641 31365 29653 31368
rect 29687 31365 29699 31399
rect 29641 31359 29699 31365
rect 30006 31356 30012 31408
rect 30064 31396 30070 31408
rect 30064 31368 30144 31396
rect 30064 31356 30070 31368
rect 22511 31300 22968 31328
rect 22511 31297 22523 31300
rect 22465 31291 22523 31297
rect 23014 31288 23020 31340
rect 23072 31328 23078 31340
rect 23293 31331 23351 31337
rect 23293 31328 23305 31331
rect 23072 31300 23305 31328
rect 23072 31288 23078 31300
rect 23293 31297 23305 31300
rect 23339 31297 23351 31331
rect 23566 31328 23572 31340
rect 23527 31300 23572 31328
rect 23293 31291 23351 31297
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 23934 31288 23940 31340
rect 23992 31328 23998 31340
rect 24118 31328 24124 31340
rect 23992 31300 24124 31328
rect 23992 31288 23998 31300
rect 24118 31288 24124 31300
rect 24176 31328 24182 31340
rect 24213 31331 24271 31337
rect 24213 31328 24225 31331
rect 24176 31300 24225 31328
rect 24176 31288 24182 31300
rect 24213 31297 24225 31300
rect 24259 31328 24271 31331
rect 25133 31331 25191 31337
rect 25133 31328 25145 31331
rect 24259 31300 25145 31328
rect 24259 31297 24271 31300
rect 24213 31291 24271 31297
rect 25133 31297 25145 31300
rect 25179 31297 25191 31331
rect 25133 31291 25191 31297
rect 25498 31288 25504 31340
rect 25556 31328 25562 31340
rect 25869 31331 25927 31337
rect 25869 31328 25881 31331
rect 25556 31300 25881 31328
rect 25556 31288 25562 31300
rect 25869 31297 25881 31300
rect 25915 31297 25927 31331
rect 25869 31291 25927 31297
rect 26053 31331 26111 31337
rect 26053 31297 26065 31331
rect 26099 31297 26111 31331
rect 26053 31291 26111 31297
rect 26145 31331 26203 31337
rect 26145 31297 26157 31331
rect 26191 31297 26203 31331
rect 26145 31291 26203 31297
rect 26237 31331 26295 31337
rect 26237 31297 26249 31331
rect 26283 31328 26295 31331
rect 26326 31328 26332 31340
rect 26283 31300 26332 31328
rect 26283 31297 26295 31300
rect 26237 31291 26295 31297
rect 13817 31263 13875 31269
rect 13817 31229 13829 31263
rect 13863 31229 13875 31263
rect 16666 31260 16672 31272
rect 13817 31223 13875 31229
rect 14200 31232 16672 31260
rect 2777 31195 2835 31201
rect 2777 31161 2789 31195
rect 2823 31192 2835 31195
rect 9950 31192 9956 31204
rect 2823 31164 9956 31192
rect 2823 31161 2835 31164
rect 2777 31155 2835 31161
rect 9950 31152 9956 31164
rect 10008 31152 10014 31204
rect 10045 31195 10103 31201
rect 10045 31161 10057 31195
rect 10091 31192 10103 31195
rect 13832 31192 13860 31223
rect 14200 31192 14228 31232
rect 16666 31220 16672 31232
rect 16724 31220 16730 31272
rect 17221 31263 17279 31269
rect 17221 31229 17233 31263
rect 17267 31229 17279 31263
rect 17221 31223 17279 31229
rect 18233 31263 18291 31269
rect 18233 31229 18245 31263
rect 18279 31260 18291 31263
rect 18506 31260 18512 31272
rect 18279 31232 18512 31260
rect 18279 31229 18291 31232
rect 18233 31223 18291 31229
rect 10091 31164 13768 31192
rect 13832 31164 14228 31192
rect 15473 31195 15531 31201
rect 10091 31161 10103 31164
rect 10045 31155 10103 31161
rect 1394 31084 1400 31136
rect 1452 31124 1458 31136
rect 1673 31127 1731 31133
rect 1673 31124 1685 31127
rect 1452 31096 1685 31124
rect 1452 31084 1458 31096
rect 1673 31093 1685 31096
rect 1719 31093 1731 31127
rect 1673 31087 1731 31093
rect 10873 31127 10931 31133
rect 10873 31093 10885 31127
rect 10919 31124 10931 31127
rect 13446 31124 13452 31136
rect 10919 31096 13452 31124
rect 10919 31093 10931 31096
rect 10873 31087 10931 31093
rect 13446 31084 13452 31096
rect 13504 31084 13510 31136
rect 13740 31124 13768 31164
rect 15473 31161 15485 31195
rect 15519 31192 15531 31195
rect 16942 31192 16948 31204
rect 15519 31164 16948 31192
rect 15519 31161 15531 31164
rect 15473 31155 15531 31161
rect 16942 31152 16948 31164
rect 17000 31152 17006 31204
rect 17236 31192 17264 31223
rect 18506 31220 18512 31232
rect 18564 31220 18570 31272
rect 22186 31220 22192 31272
rect 22244 31260 22250 31272
rect 24489 31263 24547 31269
rect 24489 31260 24501 31263
rect 22244 31232 24501 31260
rect 22244 31220 22250 31232
rect 24489 31229 24501 31232
rect 24535 31229 24547 31263
rect 24489 31223 24547 31229
rect 25409 31263 25467 31269
rect 25409 31229 25421 31263
rect 25455 31229 25467 31263
rect 25409 31223 25467 31229
rect 19521 31195 19579 31201
rect 19521 31192 19533 31195
rect 17236 31164 19533 31192
rect 18156 31136 18184 31164
rect 19521 31161 19533 31164
rect 19567 31161 19579 31195
rect 25424 31192 25452 31223
rect 19521 31155 19579 31161
rect 24136 31164 25452 31192
rect 26068 31192 26096 31291
rect 26160 31260 26188 31291
rect 26326 31288 26332 31300
rect 26384 31328 26390 31340
rect 26694 31328 26700 31340
rect 26384 31300 26700 31328
rect 26384 31288 26390 31300
rect 26694 31288 26700 31300
rect 26752 31288 26758 31340
rect 26970 31288 26976 31340
rect 27028 31288 27034 31340
rect 27062 31288 27068 31340
rect 27120 31328 27126 31340
rect 27246 31328 27252 31340
rect 27120 31300 27252 31328
rect 27120 31288 27126 31300
rect 27246 31288 27252 31300
rect 27304 31328 27310 31340
rect 28261 31331 28319 31337
rect 28261 31328 28273 31331
rect 27304 31300 28273 31328
rect 27304 31288 27310 31300
rect 28261 31297 28273 31300
rect 28307 31297 28319 31331
rect 28261 31291 28319 31297
rect 28445 31331 28503 31337
rect 28445 31297 28457 31331
rect 28491 31328 28503 31331
rect 29362 31328 29368 31340
rect 28491 31300 29368 31328
rect 28491 31297 28503 31300
rect 28445 31291 28503 31297
rect 27522 31260 27528 31272
rect 26160 31232 27528 31260
rect 27522 31220 27528 31232
rect 27580 31220 27586 31272
rect 27709 31263 27767 31269
rect 27709 31229 27721 31263
rect 27755 31260 27767 31263
rect 28460 31260 28488 31291
rect 29362 31288 29368 31300
rect 29420 31328 29426 31340
rect 29420 31300 29776 31328
rect 29420 31288 29426 31300
rect 29546 31260 29552 31272
rect 27755 31232 28488 31260
rect 29507 31232 29552 31260
rect 27755 31229 27767 31232
rect 27709 31223 27767 31229
rect 29546 31220 29552 31232
rect 29604 31220 29610 31272
rect 29748 31269 29776 31300
rect 29733 31263 29791 31269
rect 29733 31229 29745 31263
rect 29779 31260 29791 31263
rect 30006 31260 30012 31272
rect 29779 31232 30012 31260
rect 29779 31229 29791 31232
rect 29733 31223 29791 31229
rect 30006 31220 30012 31232
rect 30064 31220 30070 31272
rect 26142 31192 26148 31204
rect 26068 31164 26148 31192
rect 14182 31124 14188 31136
rect 13740 31096 14188 31124
rect 14182 31084 14188 31096
rect 14240 31084 14246 31136
rect 15194 31084 15200 31136
rect 15252 31124 15258 31136
rect 15654 31124 15660 31136
rect 15252 31096 15660 31124
rect 15252 31084 15258 31096
rect 15654 31084 15660 31096
rect 15712 31084 15718 31136
rect 16758 31124 16764 31136
rect 16719 31096 16764 31124
rect 16758 31084 16764 31096
rect 16816 31084 16822 31136
rect 18138 31084 18144 31136
rect 18196 31084 18202 31136
rect 18782 31124 18788 31136
rect 18743 31096 18788 31124
rect 18782 31084 18788 31096
rect 18840 31084 18846 31136
rect 19058 31084 19064 31136
rect 19116 31124 19122 31136
rect 23198 31124 23204 31136
rect 19116 31096 23204 31124
rect 19116 31084 19122 31096
rect 23198 31084 23204 31096
rect 23256 31084 23262 31136
rect 23477 31127 23535 31133
rect 23477 31093 23489 31127
rect 23523 31124 23535 31127
rect 23658 31124 23664 31136
rect 23523 31096 23664 31124
rect 23523 31093 23535 31096
rect 23477 31087 23535 31093
rect 23658 31084 23664 31096
rect 23716 31084 23722 31136
rect 24026 31084 24032 31136
rect 24084 31124 24090 31136
rect 24136 31124 24164 31164
rect 26142 31152 26148 31164
rect 26200 31152 26206 31204
rect 29181 31195 29239 31201
rect 29181 31192 29193 31195
rect 26252 31164 29193 31192
rect 24084 31096 24164 31124
rect 24397 31127 24455 31133
rect 24084 31084 24090 31096
rect 24397 31093 24409 31127
rect 24443 31124 24455 31127
rect 24670 31124 24676 31136
rect 24443 31096 24676 31124
rect 24443 31093 24455 31096
rect 24397 31087 24455 31093
rect 24670 31084 24676 31096
rect 24728 31124 24734 31136
rect 25130 31124 25136 31136
rect 24728 31096 25136 31124
rect 24728 31084 24734 31096
rect 25130 31084 25136 31096
rect 25188 31124 25194 31136
rect 25317 31127 25375 31133
rect 25317 31124 25329 31127
rect 25188 31096 25329 31124
rect 25188 31084 25194 31096
rect 25317 31093 25329 31096
rect 25363 31093 25375 31127
rect 25317 31087 25375 31093
rect 25590 31084 25596 31136
rect 25648 31124 25654 31136
rect 26252 31124 26280 31164
rect 29181 31161 29193 31164
rect 29227 31161 29239 31195
rect 29181 31155 29239 31161
rect 29362 31152 29368 31204
rect 29420 31192 29426 31204
rect 30116 31192 30144 31368
rect 29420 31164 30144 31192
rect 29420 31152 29426 31164
rect 25648 31096 26280 31124
rect 25648 31084 25654 31096
rect 26326 31084 26332 31136
rect 26384 31124 26390 31136
rect 27157 31127 27215 31133
rect 27157 31124 27169 31127
rect 26384 31096 27169 31124
rect 26384 31084 26390 31096
rect 27157 31093 27169 31096
rect 27203 31093 27215 31127
rect 27157 31087 27215 31093
rect 1104 31034 30820 31056
rect 1104 30982 5915 31034
rect 5967 30982 5979 31034
rect 6031 30982 6043 31034
rect 6095 30982 6107 31034
rect 6159 30982 6171 31034
rect 6223 30982 15846 31034
rect 15898 30982 15910 31034
rect 15962 30982 15974 31034
rect 16026 30982 16038 31034
rect 16090 30982 16102 31034
rect 16154 30982 25776 31034
rect 25828 30982 25840 31034
rect 25892 30982 25904 31034
rect 25956 30982 25968 31034
rect 26020 30982 26032 31034
rect 26084 30982 30820 31034
rect 31478 31016 31484 31068
rect 31536 31056 31542 31068
rect 31536 31028 31892 31056
rect 31536 31016 31542 31028
rect 1104 30960 30820 30982
rect 11422 30880 11428 30932
rect 11480 30920 11486 30932
rect 25590 30920 25596 30932
rect 11480 30892 25596 30920
rect 11480 30880 11486 30892
rect 25590 30880 25596 30892
rect 25648 30880 25654 30932
rect 26053 30923 26111 30929
rect 26053 30889 26065 30923
rect 26099 30920 26111 30923
rect 26142 30920 26148 30932
rect 26099 30892 26148 30920
rect 26099 30889 26111 30892
rect 26053 30883 26111 30889
rect 26142 30880 26148 30892
rect 26200 30880 26206 30932
rect 28350 30920 28356 30932
rect 28311 30892 28356 30920
rect 28350 30880 28356 30892
rect 28408 30880 28414 30932
rect 30098 30920 30104 30932
rect 30059 30892 30104 30920
rect 30098 30880 30104 30892
rect 30156 30880 30162 30932
rect 1854 30812 1860 30864
rect 1912 30852 1918 30864
rect 1912 30824 17264 30852
rect 1912 30812 1918 30824
rect 9950 30744 9956 30796
rect 10008 30784 10014 30796
rect 17236 30784 17264 30824
rect 17954 30812 17960 30864
rect 18012 30852 18018 30864
rect 20165 30855 20223 30861
rect 20165 30852 20177 30855
rect 18012 30824 20177 30852
rect 18012 30812 18018 30824
rect 20165 30821 20177 30824
rect 20211 30821 20223 30855
rect 20165 30815 20223 30821
rect 21450 30812 21456 30864
rect 21508 30852 21514 30864
rect 23198 30852 23204 30864
rect 21508 30824 23204 30852
rect 21508 30812 21514 30824
rect 23198 30812 23204 30824
rect 23256 30812 23262 30864
rect 24397 30855 24455 30861
rect 24397 30821 24409 30855
rect 24443 30852 24455 30855
rect 25038 30852 25044 30864
rect 24443 30824 25044 30852
rect 24443 30821 24455 30824
rect 24397 30815 24455 30821
rect 25038 30812 25044 30824
rect 25096 30812 25102 30864
rect 28276 30824 28764 30852
rect 28276 30796 28304 30824
rect 10008 30756 15884 30784
rect 17236 30756 18828 30784
rect 10008 30744 10014 30756
rect 1397 30719 1455 30725
rect 1397 30685 1409 30719
rect 1443 30716 1455 30719
rect 1762 30716 1768 30728
rect 1443 30688 1768 30716
rect 1443 30685 1455 30688
rect 1397 30679 1455 30685
rect 1762 30676 1768 30688
rect 1820 30676 1826 30728
rect 2317 30719 2375 30725
rect 2317 30685 2329 30719
rect 2363 30716 2375 30719
rect 4062 30716 4068 30728
rect 2363 30688 4068 30716
rect 2363 30685 2375 30688
rect 2317 30679 2375 30685
rect 4062 30676 4068 30688
rect 4120 30676 4126 30728
rect 9674 30716 9680 30728
rect 9635 30688 9680 30716
rect 9674 30676 9680 30688
rect 9732 30676 9738 30728
rect 9858 30716 9864 30728
rect 9819 30688 9864 30716
rect 9858 30676 9864 30688
rect 9916 30676 9922 30728
rect 11057 30719 11115 30725
rect 11057 30685 11069 30719
rect 11103 30716 11115 30719
rect 11238 30716 11244 30728
rect 11103 30688 11244 30716
rect 11103 30685 11115 30688
rect 11057 30679 11115 30685
rect 11238 30676 11244 30688
rect 11296 30676 11302 30728
rect 15427 30719 15485 30725
rect 15427 30716 15439 30719
rect 15304 30688 15439 30716
rect 10045 30651 10103 30657
rect 10045 30617 10057 30651
rect 10091 30648 10103 30651
rect 13630 30648 13636 30660
rect 10091 30620 13636 30648
rect 10091 30617 10103 30620
rect 10045 30611 10103 30617
rect 13630 30608 13636 30620
rect 13688 30608 13694 30660
rect 1578 30580 1584 30592
rect 1539 30552 1584 30580
rect 1578 30540 1584 30552
rect 1636 30540 1642 30592
rect 2130 30580 2136 30592
rect 2091 30552 2136 30580
rect 2130 30540 2136 30552
rect 2188 30540 2194 30592
rect 11238 30580 11244 30592
rect 11199 30552 11244 30580
rect 11238 30540 11244 30552
rect 11296 30540 11302 30592
rect 15194 30580 15200 30592
rect 15155 30552 15200 30580
rect 15194 30540 15200 30552
rect 15252 30540 15258 30592
rect 15304 30580 15332 30688
rect 15427 30685 15439 30688
rect 15473 30685 15485 30719
rect 15562 30716 15568 30728
rect 15523 30688 15568 30716
rect 15427 30679 15485 30685
rect 15562 30676 15568 30688
rect 15620 30676 15626 30728
rect 15856 30725 15884 30756
rect 15657 30719 15715 30725
rect 15657 30685 15669 30719
rect 15703 30685 15715 30719
rect 15657 30679 15715 30685
rect 15841 30719 15899 30725
rect 15841 30685 15853 30719
rect 15887 30685 15899 30719
rect 18690 30716 18696 30728
rect 18651 30688 18696 30716
rect 15841 30679 15899 30685
rect 15672 30648 15700 30679
rect 18690 30676 18696 30688
rect 18748 30676 18754 30728
rect 18800 30716 18828 30756
rect 18966 30744 18972 30796
rect 19024 30784 19030 30796
rect 19024 30756 20024 30784
rect 19024 30744 19030 30756
rect 19058 30716 19064 30728
rect 18800 30688 19064 30716
rect 19058 30676 19064 30688
rect 19116 30676 19122 30728
rect 19337 30719 19395 30725
rect 19337 30685 19349 30719
rect 19383 30716 19395 30719
rect 19610 30716 19616 30728
rect 19383 30688 19616 30716
rect 19383 30685 19395 30688
rect 19337 30679 19395 30685
rect 19610 30676 19616 30688
rect 19668 30676 19674 30728
rect 19996 30725 20024 30756
rect 22554 30744 22560 30796
rect 22612 30784 22618 30796
rect 24765 30787 24823 30793
rect 22612 30756 24716 30784
rect 22612 30744 22618 30756
rect 19981 30719 20039 30725
rect 19981 30685 19993 30719
rect 20027 30685 20039 30719
rect 19981 30679 20039 30685
rect 23934 30676 23940 30728
rect 23992 30716 23998 30728
rect 24581 30719 24639 30725
rect 24581 30716 24593 30719
rect 23992 30688 24593 30716
rect 23992 30676 23998 30688
rect 24581 30685 24593 30688
rect 24627 30685 24639 30719
rect 24688 30716 24716 30756
rect 24765 30753 24777 30787
rect 24811 30784 24823 30787
rect 25130 30784 25136 30796
rect 24811 30756 25136 30784
rect 24811 30753 24823 30756
rect 24765 30747 24823 30753
rect 25130 30744 25136 30756
rect 25188 30744 25194 30796
rect 25590 30744 25596 30796
rect 25648 30784 25654 30796
rect 26421 30787 26479 30793
rect 26421 30784 26433 30787
rect 25648 30756 26433 30784
rect 25648 30744 25654 30756
rect 26421 30753 26433 30756
rect 26467 30753 26479 30787
rect 26421 30747 26479 30753
rect 28077 30787 28135 30793
rect 28077 30753 28089 30787
rect 28123 30784 28135 30787
rect 28258 30784 28264 30796
rect 28123 30756 28264 30784
rect 28123 30753 28135 30756
rect 28077 30747 28135 30753
rect 28258 30744 28264 30756
rect 28316 30744 28322 30796
rect 24857 30719 24915 30725
rect 24857 30716 24869 30719
rect 24688 30688 24869 30716
rect 24581 30679 24639 30685
rect 24857 30685 24869 30688
rect 24903 30685 24915 30719
rect 24857 30679 24915 30685
rect 24946 30676 24952 30728
rect 25004 30716 25010 30728
rect 25406 30716 25412 30728
rect 25004 30688 25412 30716
rect 25004 30676 25010 30688
rect 25406 30676 25412 30688
rect 25464 30676 25470 30728
rect 26142 30676 26148 30728
rect 26200 30716 26206 30728
rect 26237 30719 26295 30725
rect 26237 30716 26249 30719
rect 26200 30688 26249 30716
rect 26200 30676 26206 30688
rect 26237 30685 26249 30688
rect 26283 30685 26295 30719
rect 26237 30679 26295 30685
rect 26513 30719 26571 30725
rect 26513 30685 26525 30719
rect 26559 30716 26571 30719
rect 27062 30716 27068 30728
rect 26559 30688 27068 30716
rect 26559 30685 26571 30688
rect 26513 30679 26571 30685
rect 27062 30676 27068 30688
rect 27120 30676 27126 30728
rect 28626 30716 28632 30728
rect 28587 30688 28632 30716
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 28736 30725 28764 30824
rect 28718 30719 28776 30725
rect 28718 30685 28730 30719
rect 28764 30685 28776 30719
rect 28718 30679 28776 30685
rect 28834 30719 28892 30725
rect 28834 30685 28846 30719
rect 28880 30716 28892 30719
rect 28997 30719 29055 30725
rect 28880 30688 28948 30716
rect 28880 30685 28892 30688
rect 28834 30679 28892 30685
rect 16206 30648 16212 30660
rect 15672 30620 16212 30648
rect 16206 30608 16212 30620
rect 16264 30608 16270 30660
rect 16301 30651 16359 30657
rect 16301 30617 16313 30651
rect 16347 30648 16359 30651
rect 20622 30648 20628 30660
rect 16347 30620 20628 30648
rect 16347 30617 16359 30620
rect 16301 30611 16359 30617
rect 20622 30608 20628 30620
rect 20680 30608 20686 30660
rect 20714 30608 20720 30660
rect 20772 30648 20778 30660
rect 26326 30648 26332 30660
rect 20772 30620 26332 30648
rect 20772 30608 20778 30620
rect 26326 30608 26332 30620
rect 26384 30608 26390 30660
rect 15470 30580 15476 30592
rect 15304 30552 15476 30580
rect 15470 30540 15476 30552
rect 15528 30540 15534 30592
rect 17586 30580 17592 30592
rect 17547 30552 17592 30580
rect 17586 30540 17592 30552
rect 17644 30540 17650 30592
rect 18506 30580 18512 30592
rect 18467 30552 18512 30580
rect 18506 30540 18512 30552
rect 18564 30540 18570 30592
rect 19518 30580 19524 30592
rect 19479 30552 19524 30580
rect 19518 30540 19524 30552
rect 19576 30540 19582 30592
rect 28718 30540 28724 30592
rect 28776 30580 28782 30592
rect 28920 30580 28948 30688
rect 28997 30685 29009 30719
rect 29043 30716 29055 30719
rect 29086 30716 29092 30728
rect 29043 30688 29092 30716
rect 29043 30685 29055 30688
rect 28997 30679 29055 30685
rect 29086 30676 29092 30688
rect 29144 30676 29150 30728
rect 29362 30676 29368 30728
rect 29420 30716 29426 30728
rect 29917 30719 29975 30725
rect 29917 30716 29929 30719
rect 29420 30688 29929 30716
rect 29420 30676 29426 30688
rect 29917 30685 29929 30688
rect 29963 30685 29975 30719
rect 31864 30716 31892 31028
rect 29917 30679 29975 30685
rect 31772 30688 31892 30716
rect 28776 30552 28948 30580
rect 28776 30540 28782 30552
rect 29086 30540 29092 30592
rect 29144 30580 29150 30592
rect 29380 30580 29408 30676
rect 31772 30660 31800 30688
rect 29546 30608 29552 30660
rect 29604 30648 29610 30660
rect 29733 30651 29791 30657
rect 29733 30648 29745 30651
rect 29604 30620 29745 30648
rect 29604 30608 29610 30620
rect 29733 30617 29745 30620
rect 29779 30648 29791 30651
rect 30374 30648 30380 30660
rect 29779 30620 30380 30648
rect 29779 30617 29791 30620
rect 29733 30611 29791 30617
rect 30374 30608 30380 30620
rect 30432 30608 30438 30660
rect 31754 30608 31760 30660
rect 31812 30608 31818 30660
rect 29144 30552 29408 30580
rect 29144 30540 29150 30552
rect 1104 30490 30820 30512
rect 1104 30438 10880 30490
rect 10932 30438 10944 30490
rect 10996 30438 11008 30490
rect 11060 30438 11072 30490
rect 11124 30438 11136 30490
rect 11188 30438 20811 30490
rect 20863 30438 20875 30490
rect 20927 30438 20939 30490
rect 20991 30438 21003 30490
rect 21055 30438 21067 30490
rect 21119 30438 30820 30490
rect 1104 30416 30820 30438
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 12897 30379 12955 30385
rect 12897 30376 12909 30379
rect 12860 30348 12909 30376
rect 12860 30336 12866 30348
rect 12897 30345 12909 30348
rect 12943 30345 12955 30379
rect 12897 30339 12955 30345
rect 13446 30336 13452 30388
rect 13504 30376 13510 30388
rect 14734 30376 14740 30388
rect 13504 30348 14740 30376
rect 13504 30336 13510 30348
rect 14734 30336 14740 30348
rect 14792 30336 14798 30388
rect 18690 30336 18696 30388
rect 18748 30376 18754 30388
rect 19886 30376 19892 30388
rect 18748 30348 19892 30376
rect 18748 30336 18754 30348
rect 19886 30336 19892 30348
rect 19944 30336 19950 30388
rect 27706 30376 27712 30388
rect 25056 30348 27712 30376
rect 11606 30268 11612 30320
rect 11664 30308 11670 30320
rect 11762 30311 11820 30317
rect 11762 30308 11774 30311
rect 11664 30280 11774 30308
rect 11664 30268 11670 30280
rect 11762 30277 11774 30280
rect 11808 30277 11820 30311
rect 11762 30271 11820 30277
rect 13722 30268 13728 30320
rect 13780 30308 13786 30320
rect 14458 30308 14464 30320
rect 13780 30280 13860 30308
rect 13780 30268 13786 30280
rect 1397 30243 1455 30249
rect 1397 30209 1409 30243
rect 1443 30240 1455 30243
rect 1670 30240 1676 30252
rect 1443 30212 1676 30240
rect 1443 30209 1455 30212
rect 1397 30203 1455 30209
rect 1670 30200 1676 30212
rect 1728 30200 1734 30252
rect 2317 30243 2375 30249
rect 2317 30209 2329 30243
rect 2363 30240 2375 30243
rect 2363 30212 6914 30240
rect 2363 30209 2375 30212
rect 2317 30203 2375 30209
rect 6886 30172 6914 30212
rect 11238 30200 11244 30252
rect 11296 30240 11302 30252
rect 13832 30249 13860 30280
rect 13924 30280 14464 30308
rect 13924 30249 13952 30280
rect 14458 30268 14464 30280
rect 14516 30268 14522 30320
rect 17954 30308 17960 30320
rect 17604 30280 17960 30308
rect 11517 30243 11575 30249
rect 11517 30240 11529 30243
rect 11296 30212 11529 30240
rect 11296 30200 11302 30212
rect 11517 30209 11529 30212
rect 11563 30209 11575 30243
rect 11517 30203 11575 30209
rect 13817 30243 13875 30249
rect 13817 30209 13829 30243
rect 13863 30209 13875 30243
rect 13817 30203 13875 30209
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30209 13967 30243
rect 13909 30203 13967 30209
rect 11422 30172 11428 30184
rect 6886 30144 11428 30172
rect 11422 30132 11428 30144
rect 11480 30132 11486 30184
rect 13078 30132 13084 30184
rect 13136 30172 13142 30184
rect 13924 30172 13952 30203
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 14056 30212 14101 30240
rect 14056 30200 14062 30212
rect 14182 30200 14188 30252
rect 14240 30240 14246 30252
rect 17604 30249 17632 30280
rect 17954 30268 17960 30280
rect 18012 30268 18018 30320
rect 19426 30308 19432 30320
rect 19387 30280 19432 30308
rect 19426 30268 19432 30280
rect 19484 30268 19490 30320
rect 19645 30311 19703 30317
rect 19645 30277 19657 30311
rect 19691 30308 19703 30311
rect 19794 30308 19800 30320
rect 19691 30280 19800 30308
rect 19691 30277 19703 30280
rect 19645 30271 19703 30277
rect 19794 30268 19800 30280
rect 19852 30268 19858 30320
rect 17589 30243 17647 30249
rect 14240 30212 14285 30240
rect 14240 30200 14246 30212
rect 17589 30209 17601 30243
rect 17635 30209 17647 30243
rect 17589 30203 17647 30209
rect 17856 30243 17914 30249
rect 17856 30209 17868 30243
rect 17902 30240 17914 30243
rect 18690 30240 18696 30252
rect 17902 30212 18696 30240
rect 17902 30209 17914 30212
rect 17856 30203 17914 30209
rect 18690 30200 18696 30212
rect 18748 30200 18754 30252
rect 19058 30200 19064 30252
rect 19116 30240 19122 30252
rect 25056 30240 25084 30348
rect 27706 30336 27712 30348
rect 27764 30336 27770 30388
rect 28074 30336 28080 30388
rect 28132 30376 28138 30388
rect 28350 30376 28356 30388
rect 28132 30348 28356 30376
rect 28132 30336 28138 30348
rect 28350 30336 28356 30348
rect 28408 30336 28414 30388
rect 30006 30376 30012 30388
rect 29656 30348 30012 30376
rect 26142 30268 26148 30320
rect 26200 30308 26206 30320
rect 26326 30308 26332 30320
rect 26200 30280 26332 30308
rect 26200 30268 26206 30280
rect 26326 30268 26332 30280
rect 26384 30268 26390 30320
rect 27614 30268 27620 30320
rect 27672 30308 27678 30320
rect 29656 30317 29684 30348
rect 30006 30336 30012 30348
rect 30064 30336 30070 30388
rect 28629 30311 28687 30317
rect 28629 30308 28641 30311
rect 27672 30280 28641 30308
rect 27672 30268 27678 30280
rect 28629 30277 28641 30280
rect 28675 30308 28687 30311
rect 29549 30311 29607 30317
rect 29549 30308 29561 30311
rect 28675 30280 29561 30308
rect 28675 30277 28687 30280
rect 28629 30271 28687 30277
rect 29549 30277 29561 30280
rect 29595 30277 29607 30311
rect 29549 30271 29607 30277
rect 29641 30311 29699 30317
rect 29641 30277 29653 30311
rect 29687 30277 29699 30311
rect 29641 30271 29699 30277
rect 19116 30212 25084 30240
rect 19116 30200 19122 30212
rect 25406 30200 25412 30252
rect 25464 30240 25470 30252
rect 27525 30243 27583 30249
rect 27525 30240 27537 30243
rect 25464 30212 27537 30240
rect 25464 30200 25470 30212
rect 27525 30209 27537 30212
rect 27571 30209 27583 30243
rect 27525 30203 27583 30209
rect 27798 30200 27804 30252
rect 27856 30240 27862 30252
rect 28077 30243 28135 30249
rect 27856 30212 28028 30240
rect 27856 30200 27862 30212
rect 13136 30144 13952 30172
rect 14016 30172 14044 30200
rect 14642 30172 14648 30184
rect 14016 30144 14648 30172
rect 13136 30132 13142 30144
rect 14642 30132 14648 30144
rect 14700 30132 14706 30184
rect 25590 30172 25596 30184
rect 25551 30144 25596 30172
rect 25590 30132 25596 30144
rect 25648 30132 25654 30184
rect 25869 30175 25927 30181
rect 25869 30141 25881 30175
rect 25915 30141 25927 30175
rect 28000 30172 28028 30212
rect 28077 30209 28089 30243
rect 28123 30240 28135 30243
rect 29362 30240 29368 30252
rect 28123 30212 29368 30240
rect 28123 30209 28135 30212
rect 28077 30203 28135 30209
rect 29362 30200 29368 30212
rect 29420 30200 29426 30252
rect 28902 30172 28908 30184
rect 28000 30144 28908 30172
rect 25869 30135 25927 30141
rect 18524 30076 19334 30104
rect 1578 30036 1584 30048
rect 1539 30008 1584 30036
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 1670 29996 1676 30048
rect 1728 30036 1734 30048
rect 2133 30039 2191 30045
rect 2133 30036 2145 30039
rect 1728 30008 2145 30036
rect 1728 29996 1734 30008
rect 2133 30005 2145 30008
rect 2179 30005 2191 30039
rect 2133 29999 2191 30005
rect 13541 30039 13599 30045
rect 13541 30005 13553 30039
rect 13587 30036 13599 30039
rect 13998 30036 14004 30048
rect 13587 30008 14004 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 13998 29996 14004 30008
rect 14056 29996 14062 30048
rect 17770 29996 17776 30048
rect 17828 30036 17834 30048
rect 18524 30036 18552 30076
rect 18966 30036 18972 30048
rect 17828 30008 18552 30036
rect 18927 30008 18972 30036
rect 17828 29996 17834 30008
rect 18966 29996 18972 30008
rect 19024 29996 19030 30048
rect 19306 30036 19334 30076
rect 25130 30064 25136 30116
rect 25188 30104 25194 30116
rect 25884 30104 25912 30135
rect 28902 30132 28908 30144
rect 28960 30132 28966 30184
rect 29546 30172 29552 30184
rect 29507 30144 29552 30172
rect 29546 30132 29552 30144
rect 29604 30132 29610 30184
rect 25188 30076 25912 30104
rect 25188 30064 25194 30076
rect 25608 30048 25636 30076
rect 26786 30064 26792 30116
rect 26844 30104 26850 30116
rect 26844 30076 29132 30104
rect 26844 30064 26850 30076
rect 19613 30039 19671 30045
rect 19613 30036 19625 30039
rect 19306 30008 19625 30036
rect 19613 30005 19625 30008
rect 19659 30005 19671 30039
rect 19794 30036 19800 30048
rect 19755 30008 19800 30036
rect 19613 29999 19671 30005
rect 19794 29996 19800 30008
rect 19852 29996 19858 30048
rect 25590 29996 25596 30048
rect 25648 29996 25654 30048
rect 27709 30039 27767 30045
rect 27709 30005 27721 30039
rect 27755 30036 27767 30039
rect 28074 30036 28080 30048
rect 27755 30008 28080 30036
rect 27755 30005 27767 30008
rect 27709 29999 27767 30005
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 28258 30036 28264 30048
rect 28219 30008 28264 30036
rect 28258 29996 28264 30008
rect 28316 29996 28322 30048
rect 29104 30045 29132 30076
rect 29089 30039 29147 30045
rect 29089 30005 29101 30039
rect 29135 30005 29147 30039
rect 29089 29999 29147 30005
rect 1104 29946 30820 29968
rect 1104 29894 5915 29946
rect 5967 29894 5979 29946
rect 6031 29894 6043 29946
rect 6095 29894 6107 29946
rect 6159 29894 6171 29946
rect 6223 29894 15846 29946
rect 15898 29894 15910 29946
rect 15962 29894 15974 29946
rect 16026 29894 16038 29946
rect 16090 29894 16102 29946
rect 16154 29894 25776 29946
rect 25828 29894 25840 29946
rect 25892 29894 25904 29946
rect 25956 29894 25968 29946
rect 26020 29894 26032 29946
rect 26084 29894 30820 29946
rect 1104 29872 30820 29894
rect 4062 29792 4068 29844
rect 4120 29832 4126 29844
rect 17034 29832 17040 29844
rect 4120 29804 12756 29832
rect 16995 29804 17040 29832
rect 4120 29792 4126 29804
rect 12728 29764 12756 29804
rect 17034 29792 17040 29804
rect 17092 29792 17098 29844
rect 18690 29832 18696 29844
rect 18651 29804 18696 29832
rect 18690 29792 18696 29804
rect 18748 29792 18754 29844
rect 19886 29832 19892 29844
rect 19847 29804 19892 29832
rect 19886 29792 19892 29804
rect 19944 29792 19950 29844
rect 25682 29792 25688 29844
rect 25740 29832 25746 29844
rect 25777 29835 25835 29841
rect 25777 29832 25789 29835
rect 25740 29804 25789 29832
rect 25740 29792 25746 29804
rect 25777 29801 25789 29804
rect 25823 29801 25835 29835
rect 26786 29832 26792 29844
rect 25777 29795 25835 29801
rect 25884 29804 26792 29832
rect 25884 29764 25912 29804
rect 26786 29792 26792 29804
rect 26844 29792 26850 29844
rect 27338 29792 27344 29844
rect 27396 29832 27402 29844
rect 27798 29832 27804 29844
rect 27396 29804 27804 29832
rect 27396 29792 27402 29804
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 30006 29832 30012 29844
rect 27908 29804 28396 29832
rect 29967 29804 30012 29832
rect 6886 29736 12434 29764
rect 12728 29736 25912 29764
rect 1397 29631 1455 29637
rect 1397 29597 1409 29631
rect 1443 29628 1455 29631
rect 2130 29628 2136 29640
rect 1443 29600 2136 29628
rect 1443 29597 1455 29600
rect 1397 29591 1455 29597
rect 2130 29588 2136 29600
rect 2188 29588 2194 29640
rect 2317 29631 2375 29637
rect 2317 29597 2329 29631
rect 2363 29628 2375 29631
rect 6886 29628 6914 29736
rect 12406 29696 12434 29736
rect 25958 29724 25964 29776
rect 26016 29764 26022 29776
rect 27065 29767 27123 29773
rect 27065 29764 27077 29767
rect 26016 29736 27077 29764
rect 26016 29724 26022 29736
rect 27065 29733 27077 29736
rect 27111 29733 27123 29767
rect 27908 29764 27936 29804
rect 28166 29764 28172 29776
rect 27065 29727 27123 29733
rect 27264 29736 27936 29764
rect 28000 29736 28172 29764
rect 20714 29696 20720 29708
rect 12406 29668 20720 29696
rect 20714 29656 20720 29668
rect 20772 29656 20778 29708
rect 22094 29696 22100 29708
rect 21284 29668 22100 29696
rect 12710 29628 12716 29640
rect 2363 29600 6914 29628
rect 12671 29600 12716 29628
rect 2363 29597 2375 29600
rect 2317 29591 2375 29597
rect 12710 29588 12716 29600
rect 12768 29588 12774 29640
rect 12989 29631 13047 29637
rect 12989 29597 13001 29631
rect 13035 29628 13047 29631
rect 13078 29628 13084 29640
rect 13035 29600 13084 29628
rect 13035 29597 13047 29600
rect 12989 29591 13047 29597
rect 13078 29588 13084 29600
rect 13136 29588 13142 29640
rect 14366 29637 14372 29640
rect 14349 29631 14372 29637
rect 14349 29597 14361 29631
rect 14349 29591 14372 29597
rect 14366 29588 14372 29591
rect 14424 29588 14430 29640
rect 14461 29631 14519 29637
rect 14461 29597 14473 29631
rect 14507 29597 14519 29631
rect 14461 29591 14519 29597
rect 14553 29628 14611 29634
rect 14642 29628 14648 29640
rect 14553 29594 14565 29628
rect 14599 29600 14648 29628
rect 14599 29594 14611 29600
rect 14476 29504 14504 29591
rect 14553 29588 14611 29594
rect 14642 29588 14648 29600
rect 14700 29588 14706 29640
rect 14734 29588 14740 29640
rect 14792 29628 14798 29640
rect 15746 29628 15752 29640
rect 14792 29600 14837 29628
rect 15707 29600 15752 29628
rect 14792 29588 14798 29600
rect 15746 29588 15752 29600
rect 15804 29588 15810 29640
rect 18049 29631 18107 29637
rect 18049 29597 18061 29631
rect 18095 29628 18107 29631
rect 18782 29628 18788 29640
rect 18095 29600 18788 29628
rect 18095 29597 18107 29600
rect 18049 29591 18107 29597
rect 18782 29588 18788 29600
rect 18840 29588 18846 29640
rect 19245 29631 19303 29637
rect 19245 29597 19257 29631
rect 19291 29628 19303 29631
rect 19794 29628 19800 29640
rect 19291 29600 19800 29628
rect 19291 29597 19303 29600
rect 19245 29591 19303 29597
rect 19794 29588 19800 29600
rect 19852 29588 19858 29640
rect 21284 29637 21312 29668
rect 22094 29656 22100 29668
rect 22152 29696 22158 29708
rect 22738 29696 22744 29708
rect 22152 29668 22744 29696
rect 22152 29656 22158 29668
rect 22738 29656 22744 29668
rect 22796 29656 22802 29708
rect 25590 29656 25596 29708
rect 25648 29696 25654 29708
rect 26145 29699 26203 29705
rect 26145 29696 26157 29699
rect 25648 29668 26157 29696
rect 25648 29656 25654 29668
rect 26145 29665 26157 29668
rect 26191 29665 26203 29699
rect 26145 29659 26203 29665
rect 21085 29631 21143 29637
rect 21085 29597 21097 29631
rect 21131 29597 21143 29631
rect 21085 29591 21143 29597
rect 21177 29631 21235 29637
rect 21177 29597 21189 29631
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 21269 29631 21327 29637
rect 21269 29597 21281 29631
rect 21315 29597 21327 29631
rect 21269 29591 21327 29597
rect 21453 29631 21511 29637
rect 21453 29597 21465 29631
rect 21499 29628 21511 29631
rect 22830 29628 22836 29640
rect 21499 29600 22836 29628
rect 21499 29597 21511 29600
rect 21453 29591 21511 29597
rect 1578 29492 1584 29504
rect 1539 29464 1584 29492
rect 1578 29452 1584 29464
rect 1636 29452 1642 29504
rect 2130 29492 2136 29504
rect 2091 29464 2136 29492
rect 2130 29452 2136 29464
rect 2188 29452 2194 29504
rect 14093 29495 14151 29501
rect 14093 29461 14105 29495
rect 14139 29492 14151 29495
rect 14182 29492 14188 29504
rect 14139 29464 14188 29492
rect 14139 29461 14151 29464
rect 14093 29455 14151 29461
rect 14182 29452 14188 29464
rect 14240 29452 14246 29504
rect 14458 29452 14464 29504
rect 14516 29452 14522 29504
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20809 29495 20867 29501
rect 20809 29492 20821 29495
rect 20036 29464 20821 29492
rect 20036 29452 20042 29464
rect 20809 29461 20821 29464
rect 20855 29461 20867 29495
rect 21100 29492 21128 29591
rect 21192 29560 21220 29591
rect 22830 29588 22836 29600
rect 22888 29588 22894 29640
rect 25866 29588 25872 29640
rect 25924 29628 25930 29640
rect 25961 29631 26019 29637
rect 25961 29628 25973 29631
rect 25924 29600 25973 29628
rect 25924 29588 25930 29600
rect 25961 29597 25973 29600
rect 26007 29597 26019 29631
rect 25961 29591 26019 29597
rect 26237 29631 26295 29637
rect 26237 29597 26249 29631
rect 26283 29597 26295 29631
rect 26237 29591 26295 29597
rect 26881 29631 26939 29637
rect 26881 29597 26893 29631
rect 26927 29628 26939 29631
rect 27062 29628 27068 29640
rect 26927 29600 27068 29628
rect 26927 29597 26939 29600
rect 26881 29591 26939 29597
rect 21358 29560 21364 29572
rect 21192 29532 21364 29560
rect 21358 29520 21364 29532
rect 21416 29560 21422 29572
rect 22002 29560 22008 29572
rect 21416 29532 22008 29560
rect 21416 29520 21422 29532
rect 22002 29520 22008 29532
rect 22060 29520 22066 29572
rect 23106 29520 23112 29572
rect 23164 29560 23170 29572
rect 26050 29560 26056 29572
rect 23164 29532 26056 29560
rect 23164 29520 23170 29532
rect 26050 29520 26056 29532
rect 26108 29560 26114 29572
rect 26252 29560 26280 29591
rect 27062 29588 27068 29600
rect 27120 29588 27126 29640
rect 26108 29532 26280 29560
rect 26108 29520 26114 29532
rect 27264 29504 27292 29736
rect 27820 29631 27878 29637
rect 27820 29597 27832 29631
rect 27866 29628 27878 29631
rect 28000 29628 28028 29736
rect 28166 29724 28172 29736
rect 28224 29724 28230 29776
rect 28368 29764 28396 29804
rect 30006 29792 30012 29804
rect 30064 29792 30070 29844
rect 28368 29736 29868 29764
rect 28074 29656 28080 29708
rect 28132 29696 28138 29708
rect 28132 29668 28212 29696
rect 28132 29656 28138 29668
rect 27866 29600 28028 29628
rect 28077 29609 28135 29615
rect 27866 29597 27878 29600
rect 27820 29591 27878 29597
rect 28077 29575 28089 29609
rect 28123 29606 28135 29609
rect 28184 29606 28212 29668
rect 28123 29578 28212 29606
rect 28350 29588 28356 29640
rect 28408 29628 28414 29640
rect 29840 29637 29868 29736
rect 28721 29631 28779 29637
rect 28721 29628 28733 29631
rect 28408 29600 28733 29628
rect 28408 29588 28414 29600
rect 28721 29597 28733 29600
rect 28767 29597 28779 29631
rect 28721 29591 28779 29597
rect 29825 29631 29883 29637
rect 29825 29597 29837 29631
rect 29871 29597 29883 29631
rect 29825 29591 29883 29597
rect 28123 29575 28135 29578
rect 27706 29520 27712 29572
rect 27764 29560 27770 29572
rect 28077 29569 28135 29575
rect 27985 29563 28043 29569
rect 27985 29560 27997 29563
rect 27764 29532 27997 29560
rect 27764 29520 27770 29532
rect 27985 29529 27997 29532
rect 28031 29529 28043 29563
rect 27985 29523 28043 29529
rect 21542 29492 21548 29504
rect 21100 29464 21548 29492
rect 20809 29455 20867 29461
rect 21542 29452 21548 29464
rect 21600 29452 21606 29504
rect 25866 29452 25872 29504
rect 25924 29492 25930 29504
rect 26326 29492 26332 29504
rect 25924 29464 26332 29492
rect 25924 29452 25930 29464
rect 26326 29452 26332 29464
rect 26384 29452 26390 29504
rect 27246 29452 27252 29504
rect 27304 29452 27310 29504
rect 27614 29452 27620 29504
rect 27672 29492 27678 29504
rect 28902 29492 28908 29504
rect 27672 29464 27717 29492
rect 28863 29464 28908 29492
rect 27672 29452 27678 29464
rect 28902 29452 28908 29464
rect 28960 29452 28966 29504
rect 1104 29402 30820 29424
rect 1104 29350 10880 29402
rect 10932 29350 10944 29402
rect 10996 29350 11008 29402
rect 11060 29350 11072 29402
rect 11124 29350 11136 29402
rect 11188 29350 20811 29402
rect 20863 29350 20875 29402
rect 20927 29350 20939 29402
rect 20991 29350 21003 29402
rect 21055 29350 21067 29402
rect 21119 29350 30820 29402
rect 1104 29328 30820 29350
rect 15102 29248 15108 29300
rect 15160 29288 15166 29300
rect 15197 29291 15255 29297
rect 15197 29288 15209 29291
rect 15160 29260 15209 29288
rect 15160 29248 15166 29260
rect 15197 29257 15209 29260
rect 15243 29257 15255 29291
rect 15197 29251 15255 29257
rect 16850 29248 16856 29300
rect 16908 29288 16914 29300
rect 18049 29291 18107 29297
rect 18049 29288 18061 29291
rect 16908 29260 18061 29288
rect 16908 29248 16914 29260
rect 18049 29257 18061 29260
rect 18095 29257 18107 29291
rect 18049 29251 18107 29257
rect 21821 29291 21879 29297
rect 21821 29257 21833 29291
rect 21867 29288 21879 29291
rect 21910 29288 21916 29300
rect 21867 29260 21916 29288
rect 21867 29257 21879 29260
rect 21821 29251 21879 29257
rect 21910 29248 21916 29260
rect 21968 29248 21974 29300
rect 22830 29288 22836 29300
rect 22791 29260 22836 29288
rect 22830 29248 22836 29260
rect 22888 29248 22894 29300
rect 23382 29248 23388 29300
rect 23440 29248 23446 29300
rect 25130 29248 25136 29300
rect 25188 29288 25194 29300
rect 25188 29260 27476 29288
rect 25188 29248 25194 29260
rect 13078 29220 13084 29232
rect 12912 29192 13084 29220
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29152 1455 29155
rect 1670 29152 1676 29164
rect 1443 29124 1676 29152
rect 1443 29121 1455 29124
rect 1397 29115 1455 29121
rect 1670 29112 1676 29124
rect 1728 29112 1734 29164
rect 12618 29112 12624 29164
rect 12676 29152 12682 29164
rect 12912 29161 12940 29192
rect 13078 29180 13084 29192
rect 13136 29180 13142 29232
rect 13906 29220 13912 29232
rect 13867 29192 13912 29220
rect 13906 29180 13912 29192
rect 13964 29180 13970 29232
rect 16942 29229 16948 29232
rect 16936 29220 16948 29229
rect 16903 29192 16948 29220
rect 16936 29183 16948 29192
rect 16942 29180 16948 29183
rect 17000 29180 17006 29232
rect 19610 29220 19616 29232
rect 19306 29192 19616 29220
rect 12759 29155 12817 29161
rect 12759 29152 12771 29155
rect 12676 29124 12771 29152
rect 12676 29112 12682 29124
rect 12759 29121 12771 29124
rect 12805 29121 12817 29155
rect 12759 29115 12817 29121
rect 12897 29155 12955 29161
rect 12897 29121 12909 29155
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 12989 29155 13047 29161
rect 12989 29121 13001 29155
rect 13035 29121 13047 29155
rect 12989 29115 13047 29121
rect 13173 29155 13231 29161
rect 13173 29121 13185 29155
rect 13219 29152 13231 29155
rect 13354 29152 13360 29164
rect 13219 29124 13360 29152
rect 13219 29121 13231 29124
rect 13173 29115 13231 29121
rect 13004 29084 13032 29115
rect 13354 29112 13360 29124
rect 13412 29112 13418 29164
rect 13722 29112 13728 29164
rect 13780 29152 13786 29164
rect 15746 29152 15752 29164
rect 13780 29124 15752 29152
rect 13780 29112 13786 29124
rect 15746 29112 15752 29124
rect 15804 29152 15810 29164
rect 19306 29152 19334 29192
rect 19610 29180 19616 29192
rect 19668 29180 19674 29232
rect 19788 29223 19846 29229
rect 19788 29189 19800 29223
rect 19834 29220 19846 29223
rect 19978 29220 19984 29232
rect 19834 29192 19984 29220
rect 19834 29189 19846 29192
rect 19788 29183 19846 29189
rect 19978 29180 19984 29192
rect 20036 29180 20042 29232
rect 20990 29180 20996 29232
rect 21048 29220 21054 29232
rect 21634 29220 21640 29232
rect 21048 29192 21640 29220
rect 21048 29180 21054 29192
rect 21634 29180 21640 29192
rect 21692 29220 21698 29232
rect 21692 29192 22324 29220
rect 21692 29180 21698 29192
rect 19518 29152 19524 29164
rect 15804 29124 19334 29152
rect 19479 29124 19524 29152
rect 15804 29112 15810 29124
rect 19518 29112 19524 29124
rect 19576 29112 19582 29164
rect 21542 29112 21548 29164
rect 21600 29152 21606 29164
rect 22296 29161 22324 29192
rect 22738 29180 22744 29232
rect 22796 29220 22802 29232
rect 23400 29220 23428 29248
rect 22796 29192 23428 29220
rect 22796 29180 22802 29192
rect 22005 29155 22063 29161
rect 22005 29152 22017 29155
rect 21600 29124 22017 29152
rect 21600 29112 21606 29124
rect 22005 29121 22017 29124
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29152 22339 29155
rect 22370 29152 22376 29164
rect 22327 29124 22376 29152
rect 22327 29121 22339 29124
rect 22281 29115 22339 29121
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 22646 29112 22652 29164
rect 22704 29152 22710 29164
rect 23017 29155 23075 29161
rect 23017 29152 23029 29155
rect 22704 29124 23029 29152
rect 22704 29112 22710 29124
rect 23017 29121 23029 29124
rect 23063 29121 23075 29155
rect 23017 29115 23075 29121
rect 23106 29112 23112 29164
rect 23164 29152 23170 29164
rect 23308 29161 23336 29192
rect 25590 29180 25596 29232
rect 25648 29220 25654 29232
rect 27246 29220 27252 29232
rect 25648 29192 27252 29220
rect 25648 29180 25654 29192
rect 27246 29180 27252 29192
rect 27304 29180 27310 29232
rect 23293 29155 23351 29161
rect 23164 29124 23209 29152
rect 23164 29112 23170 29124
rect 23293 29121 23305 29155
rect 23339 29121 23351 29155
rect 23293 29115 23351 29121
rect 23385 29155 23443 29161
rect 23385 29121 23397 29155
rect 23431 29121 23443 29155
rect 23385 29115 23443 29121
rect 14642 29084 14648 29096
rect 13004 29056 14648 29084
rect 14642 29044 14648 29056
rect 14700 29044 14706 29096
rect 16666 29084 16672 29096
rect 16627 29056 16672 29084
rect 16666 29044 16672 29056
rect 16724 29044 16730 29096
rect 22830 29044 22836 29096
rect 22888 29084 22894 29096
rect 23400 29084 23428 29115
rect 26050 29112 26056 29164
rect 26108 29152 26114 29164
rect 27448 29152 27476 29260
rect 27706 29248 27712 29300
rect 27764 29288 27770 29300
rect 28166 29288 28172 29300
rect 27764 29260 28172 29288
rect 27764 29248 27770 29260
rect 28166 29248 28172 29260
rect 28224 29248 28230 29300
rect 28350 29288 28356 29300
rect 28311 29260 28356 29288
rect 28350 29248 28356 29260
rect 28408 29248 28414 29300
rect 30009 29291 30067 29297
rect 30009 29257 30021 29291
rect 30055 29288 30067 29291
rect 30098 29288 30104 29300
rect 30055 29260 30104 29288
rect 30055 29257 30067 29260
rect 30009 29251 30067 29257
rect 30098 29248 30104 29260
rect 30156 29248 30162 29300
rect 28368 29192 28856 29220
rect 28368 29164 28396 29192
rect 27706 29161 27712 29164
rect 27663 29155 27712 29161
rect 26108 29124 26234 29152
rect 27448 29124 27568 29152
rect 26108 29112 26114 29124
rect 22888 29056 23428 29084
rect 22888 29044 22894 29056
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 12342 28976 12348 29028
rect 12400 29016 12406 29028
rect 12529 29019 12587 29025
rect 12529 29016 12541 29019
rect 12400 28988 12541 29016
rect 12400 28976 12406 28988
rect 12529 28985 12541 28988
rect 12575 28985 12587 29019
rect 12529 28979 12587 28985
rect 21818 28976 21824 29028
rect 21876 29016 21882 29028
rect 22097 29019 22155 29025
rect 22097 29016 22109 29019
rect 21876 28988 22109 29016
rect 21876 28976 21882 28988
rect 22097 28985 22109 28988
rect 22143 28985 22155 29019
rect 22097 28979 22155 28985
rect 22189 29019 22247 29025
rect 22189 28985 22201 29019
rect 22235 28985 22247 29019
rect 26206 29016 26234 29124
rect 27540 29096 27568 29124
rect 27663 29121 27675 29155
rect 27709 29121 27712 29155
rect 27663 29115 27712 29121
rect 27706 29112 27712 29115
rect 27764 29112 27770 29164
rect 27801 29155 27859 29161
rect 27801 29121 27813 29155
rect 27847 29121 27859 29155
rect 27801 29115 27859 29121
rect 27893 29155 27951 29161
rect 27893 29121 27905 29155
rect 27939 29152 27951 29155
rect 27982 29152 27988 29164
rect 27939 29124 27988 29152
rect 27939 29121 27951 29124
rect 27893 29115 27951 29121
rect 27246 29044 27252 29096
rect 27304 29084 27310 29096
rect 27433 29087 27491 29093
rect 27433 29084 27445 29087
rect 27304 29056 27445 29084
rect 27304 29044 27310 29056
rect 27433 29053 27445 29056
rect 27479 29053 27491 29087
rect 27433 29047 27491 29053
rect 27522 29044 27528 29096
rect 27580 29044 27586 29096
rect 27816 29016 27844 29115
rect 27982 29112 27988 29124
rect 28040 29112 28046 29164
rect 28350 29112 28356 29164
rect 28408 29112 28414 29164
rect 28828 29161 28856 29192
rect 28609 29155 28667 29161
rect 28609 29121 28621 29155
rect 28655 29152 28667 29155
rect 28721 29155 28779 29161
rect 28655 29121 28672 29152
rect 28609 29115 28672 29121
rect 28721 29121 28733 29155
rect 28767 29121 28779 29155
rect 28721 29115 28779 29121
rect 28813 29155 28871 29161
rect 28813 29121 28825 29155
rect 28859 29121 28871 29155
rect 28813 29115 28871 29121
rect 28997 29155 29055 29161
rect 28997 29121 29009 29155
rect 29043 29152 29055 29155
rect 29454 29152 29460 29164
rect 29043 29124 29460 29152
rect 29043 29121 29055 29124
rect 28997 29115 29055 29121
rect 28644 29028 28672 29115
rect 28736 29084 28764 29115
rect 29454 29112 29460 29124
rect 29512 29112 29518 29164
rect 29825 29155 29883 29161
rect 29825 29121 29837 29155
rect 29871 29152 29883 29155
rect 30006 29152 30012 29164
rect 29871 29124 30012 29152
rect 29871 29121 29883 29124
rect 29825 29115 29883 29121
rect 30006 29112 30012 29124
rect 30064 29112 30070 29164
rect 31386 29084 31392 29096
rect 28736 29056 31392 29084
rect 31386 29044 31392 29056
rect 31444 29044 31450 29096
rect 26206 28988 27844 29016
rect 22189 28979 22247 28985
rect 10594 28908 10600 28960
rect 10652 28948 10658 28960
rect 17310 28948 17316 28960
rect 10652 28920 17316 28948
rect 10652 28908 10658 28920
rect 17310 28908 17316 28920
rect 17368 28908 17374 28960
rect 20901 28951 20959 28957
rect 20901 28917 20913 28951
rect 20947 28948 20959 28951
rect 21174 28948 21180 28960
rect 20947 28920 21180 28948
rect 20947 28917 20959 28920
rect 20901 28911 20959 28917
rect 21174 28908 21180 28920
rect 21232 28908 21238 28960
rect 22002 28908 22008 28960
rect 22060 28948 22066 28960
rect 22204 28948 22232 28979
rect 28626 28976 28632 29028
rect 28684 28976 28690 29028
rect 22060 28920 22232 28948
rect 22060 28908 22066 28920
rect 27614 28908 27620 28960
rect 27672 28948 27678 28960
rect 29454 28948 29460 28960
rect 27672 28920 29460 28948
rect 27672 28908 27678 28920
rect 29454 28908 29460 28920
rect 29512 28908 29518 28960
rect 1104 28858 30820 28880
rect 1104 28806 5915 28858
rect 5967 28806 5979 28858
rect 6031 28806 6043 28858
rect 6095 28806 6107 28858
rect 6159 28806 6171 28858
rect 6223 28806 15846 28858
rect 15898 28806 15910 28858
rect 15962 28806 15974 28858
rect 16026 28806 16038 28858
rect 16090 28806 16102 28858
rect 16154 28806 25776 28858
rect 25828 28806 25840 28858
rect 25892 28806 25904 28858
rect 25956 28806 25968 28858
rect 26020 28806 26032 28858
rect 26084 28806 30820 28858
rect 1104 28784 30820 28806
rect 15565 28747 15623 28753
rect 15565 28713 15577 28747
rect 15611 28744 15623 28747
rect 16666 28744 16672 28756
rect 15611 28716 16672 28744
rect 15611 28713 15623 28716
rect 15565 28707 15623 28713
rect 16666 28704 16672 28716
rect 16724 28704 16730 28756
rect 19610 28704 19616 28756
rect 19668 28744 19674 28756
rect 20346 28744 20352 28756
rect 19668 28716 20352 28744
rect 19668 28704 19674 28716
rect 20346 28704 20352 28716
rect 20404 28704 20410 28756
rect 25130 28744 25136 28756
rect 25091 28716 25136 28744
rect 25130 28704 25136 28716
rect 25188 28704 25194 28756
rect 27614 28704 27620 28756
rect 27672 28744 27678 28756
rect 28810 28744 28816 28756
rect 27672 28716 28816 28744
rect 27672 28704 27678 28716
rect 28810 28704 28816 28716
rect 28868 28704 28874 28756
rect 14458 28636 14464 28688
rect 14516 28636 14522 28688
rect 17310 28636 17316 28688
rect 17368 28676 17374 28688
rect 17368 28648 20208 28676
rect 17368 28636 17374 28648
rect 1397 28543 1455 28549
rect 1397 28509 1409 28543
rect 1443 28540 1455 28543
rect 2130 28540 2136 28552
rect 1443 28512 2136 28540
rect 1443 28509 1455 28512
rect 1397 28503 1455 28509
rect 2130 28500 2136 28512
rect 2188 28500 2194 28552
rect 14467 28549 14495 28636
rect 14642 28608 14648 28620
rect 14568 28580 14648 28608
rect 14568 28549 14596 28580
rect 14642 28568 14648 28580
rect 14700 28568 14706 28620
rect 17586 28608 17592 28620
rect 16132 28580 17592 28608
rect 14349 28543 14407 28549
rect 14349 28540 14361 28543
rect 14292 28512 14361 28540
rect 2222 28432 2228 28484
rect 2280 28472 2286 28484
rect 10778 28472 10784 28484
rect 2280 28444 10784 28472
rect 2280 28432 2286 28444
rect 10778 28432 10784 28444
rect 10836 28432 10842 28484
rect 14292 28472 14320 28512
rect 14349 28509 14361 28512
rect 14395 28509 14407 28543
rect 14349 28503 14407 28509
rect 14442 28543 14500 28549
rect 14442 28509 14454 28543
rect 14488 28509 14500 28543
rect 14442 28503 14500 28509
rect 14558 28543 14616 28549
rect 14558 28509 14570 28543
rect 14604 28509 14616 28543
rect 14734 28540 14740 28552
rect 14695 28512 14740 28540
rect 14558 28503 14616 28509
rect 14734 28500 14740 28512
rect 14792 28500 14798 28552
rect 15381 28543 15439 28549
rect 15381 28509 15393 28543
rect 15427 28540 15439 28543
rect 15470 28540 15476 28552
rect 15427 28512 15476 28540
rect 15427 28509 15439 28512
rect 15381 28503 15439 28509
rect 15470 28500 15476 28512
rect 15528 28500 15534 28552
rect 16132 28549 16160 28580
rect 17586 28568 17592 28580
rect 17644 28568 17650 28620
rect 18601 28611 18659 28617
rect 18601 28577 18613 28611
rect 18647 28608 18659 28611
rect 19337 28611 19395 28617
rect 19337 28608 19349 28611
rect 18647 28580 19349 28608
rect 18647 28577 18659 28580
rect 18601 28571 18659 28577
rect 19337 28577 19349 28580
rect 19383 28577 19395 28611
rect 19337 28571 19395 28577
rect 19521 28611 19579 28617
rect 19521 28577 19533 28611
rect 19567 28608 19579 28611
rect 20070 28608 20076 28620
rect 19567 28580 20076 28608
rect 19567 28577 19579 28580
rect 19521 28571 19579 28577
rect 20070 28568 20076 28580
rect 20128 28568 20134 28620
rect 16117 28543 16175 28549
rect 16117 28509 16129 28543
rect 16163 28509 16175 28543
rect 16117 28503 16175 28509
rect 16853 28543 16911 28549
rect 16853 28509 16865 28543
rect 16899 28540 16911 28543
rect 17034 28540 17040 28552
rect 16899 28512 17040 28540
rect 16899 28509 16911 28512
rect 16853 28503 16911 28509
rect 17034 28500 17040 28512
rect 17092 28500 17098 28552
rect 18322 28500 18328 28552
rect 18380 28540 18386 28552
rect 18509 28543 18567 28549
rect 18509 28540 18521 28543
rect 18380 28512 18521 28540
rect 18380 28500 18386 28512
rect 18509 28509 18521 28512
rect 18555 28509 18567 28543
rect 18509 28503 18567 28509
rect 18693 28543 18751 28549
rect 18693 28509 18705 28543
rect 18739 28509 18751 28543
rect 18693 28503 18751 28509
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28540 19303 28543
rect 19702 28540 19708 28552
rect 19291 28512 19708 28540
rect 19291 28509 19303 28512
rect 19245 28503 19303 28509
rect 16301 28475 16359 28481
rect 14292 28444 15424 28472
rect 15396 28416 15424 28444
rect 16301 28441 16313 28475
rect 16347 28472 16359 28475
rect 16482 28472 16488 28484
rect 16347 28444 16488 28472
rect 16347 28441 16359 28444
rect 16301 28435 16359 28441
rect 16482 28432 16488 28444
rect 16540 28432 16546 28484
rect 18708 28472 18736 28503
rect 19702 28500 19708 28512
rect 19760 28500 19766 28552
rect 19610 28472 19616 28484
rect 18708 28444 19616 28472
rect 19610 28432 19616 28444
rect 19668 28432 19674 28484
rect 20070 28472 20076 28484
rect 20031 28444 20076 28472
rect 20070 28432 20076 28444
rect 20128 28432 20134 28484
rect 20180 28472 20208 28648
rect 20530 28636 20536 28688
rect 20588 28676 20594 28688
rect 20588 28648 25544 28676
rect 20588 28636 20594 28648
rect 22649 28611 22707 28617
rect 22649 28608 22661 28611
rect 21192 28580 22661 28608
rect 21192 28552 21220 28580
rect 22649 28577 22661 28580
rect 22695 28577 22707 28611
rect 22649 28571 22707 28577
rect 22848 28580 24624 28608
rect 20990 28540 20996 28552
rect 20951 28512 20996 28540
rect 20990 28500 20996 28512
rect 21048 28500 21054 28552
rect 21174 28540 21180 28552
rect 21135 28512 21180 28540
rect 21174 28500 21180 28512
rect 21232 28500 21238 28552
rect 21729 28543 21787 28549
rect 21729 28509 21741 28543
rect 21775 28540 21787 28543
rect 21818 28540 21824 28552
rect 21775 28512 21824 28540
rect 21775 28509 21787 28512
rect 21729 28503 21787 28509
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 22002 28540 22008 28552
rect 21963 28512 22008 28540
rect 22002 28500 22008 28512
rect 22060 28500 22066 28552
rect 22848 28472 22876 28580
rect 24596 28549 24624 28580
rect 22925 28543 22983 28549
rect 22925 28509 22937 28543
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 24581 28543 24639 28549
rect 24581 28509 24593 28543
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 24949 28543 25007 28549
rect 24949 28509 24961 28543
rect 24995 28540 25007 28543
rect 25130 28540 25136 28552
rect 24995 28512 25136 28540
rect 24995 28509 25007 28512
rect 24949 28503 25007 28509
rect 20180 28444 22876 28472
rect 1578 28404 1584 28416
rect 1539 28376 1584 28404
rect 1578 28364 1584 28376
rect 1636 28364 1642 28416
rect 14093 28407 14151 28413
rect 14093 28373 14105 28407
rect 14139 28404 14151 28407
rect 15286 28404 15292 28416
rect 14139 28376 15292 28404
rect 14139 28373 14151 28376
rect 14093 28367 14151 28373
rect 15286 28364 15292 28376
rect 15344 28364 15350 28416
rect 15378 28364 15384 28416
rect 15436 28364 15442 28416
rect 16942 28404 16948 28416
rect 16903 28376 16948 28404
rect 16942 28364 16948 28376
rect 17000 28364 17006 28416
rect 19518 28404 19524 28416
rect 19479 28376 19524 28404
rect 19518 28364 19524 28376
rect 19576 28364 19582 28416
rect 20162 28404 20168 28416
rect 20123 28376 20168 28404
rect 20162 28364 20168 28376
rect 20220 28364 20226 28416
rect 20993 28407 21051 28413
rect 20993 28373 21005 28407
rect 21039 28404 21051 28407
rect 21266 28404 21272 28416
rect 21039 28376 21272 28404
rect 21039 28373 21051 28376
rect 20993 28367 21051 28373
rect 21266 28364 21272 28376
rect 21324 28364 21330 28416
rect 21542 28364 21548 28416
rect 21600 28404 21606 28416
rect 22940 28404 22968 28503
rect 25130 28500 25136 28512
rect 25188 28500 25194 28552
rect 24762 28472 24768 28484
rect 24723 28444 24768 28472
rect 24762 28432 24768 28444
rect 24820 28432 24826 28484
rect 24857 28475 24915 28481
rect 24857 28441 24869 28475
rect 24903 28472 24915 28475
rect 25038 28472 25044 28484
rect 24903 28444 25044 28472
rect 24903 28441 24915 28444
rect 24857 28435 24915 28441
rect 25038 28432 25044 28444
rect 25096 28432 25102 28484
rect 25516 28472 25544 28648
rect 29638 28636 29644 28688
rect 29696 28676 29702 28688
rect 30098 28676 30104 28688
rect 29696 28648 30104 28676
rect 29696 28636 29702 28648
rect 30098 28636 30104 28648
rect 30156 28636 30162 28688
rect 28445 28611 28503 28617
rect 28445 28577 28457 28611
rect 28491 28608 28503 28611
rect 28626 28608 28632 28620
rect 28491 28580 28632 28608
rect 28491 28577 28503 28580
rect 28445 28571 28503 28577
rect 28626 28568 28632 28580
rect 28684 28568 28690 28620
rect 29086 28568 29092 28620
rect 29144 28568 29150 28620
rect 27433 28543 27491 28549
rect 27433 28509 27445 28543
rect 27479 28540 27491 28543
rect 27614 28540 27620 28552
rect 27479 28512 27620 28540
rect 27479 28509 27491 28512
rect 27433 28503 27491 28509
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 27709 28543 27767 28549
rect 27709 28509 27721 28543
rect 27755 28540 27767 28543
rect 27982 28540 27988 28552
rect 27755 28512 27988 28540
rect 27755 28509 27767 28512
rect 27709 28503 27767 28509
rect 27982 28500 27988 28512
rect 28040 28500 28046 28552
rect 28074 28500 28080 28552
rect 28132 28540 28138 28552
rect 28169 28543 28227 28549
rect 28169 28540 28181 28543
rect 28132 28512 28181 28540
rect 28132 28500 28138 28512
rect 28169 28509 28181 28512
rect 28215 28509 28227 28543
rect 28169 28503 28227 28509
rect 26786 28472 26792 28484
rect 25516 28444 26792 28472
rect 26786 28432 26792 28444
rect 26844 28472 26850 28484
rect 26844 28444 27660 28472
rect 26844 28432 26850 28444
rect 27246 28404 27252 28416
rect 21600 28376 22968 28404
rect 27207 28376 27252 28404
rect 21600 28364 21606 28376
rect 27246 28364 27252 28376
rect 27304 28364 27310 28416
rect 27632 28413 27660 28444
rect 27617 28407 27675 28413
rect 27617 28373 27629 28407
rect 27663 28373 27675 28407
rect 27617 28367 27675 28373
rect 27982 28364 27988 28416
rect 28040 28404 28046 28416
rect 28442 28404 28448 28416
rect 28040 28376 28448 28404
rect 28040 28364 28046 28376
rect 28442 28364 28448 28376
rect 28500 28364 28506 28416
rect 28994 28364 29000 28416
rect 29052 28404 29058 28416
rect 29104 28404 29132 28568
rect 29638 28500 29644 28552
rect 29696 28540 29702 28552
rect 29825 28543 29883 28549
rect 29825 28540 29837 28543
rect 29696 28512 29837 28540
rect 29696 28500 29702 28512
rect 29825 28509 29837 28512
rect 29871 28509 29883 28543
rect 29825 28503 29883 28509
rect 30006 28404 30012 28416
rect 29052 28376 29132 28404
rect 29967 28376 30012 28404
rect 29052 28364 29058 28376
rect 30006 28364 30012 28376
rect 30064 28364 30070 28416
rect 1104 28314 30820 28336
rect 1104 28262 10880 28314
rect 10932 28262 10944 28314
rect 10996 28262 11008 28314
rect 11060 28262 11072 28314
rect 11124 28262 11136 28314
rect 11188 28262 20811 28314
rect 20863 28262 20875 28314
rect 20927 28262 20939 28314
rect 20991 28262 21003 28314
rect 21055 28262 21067 28314
rect 21119 28262 30820 28314
rect 1104 28240 30820 28262
rect 13814 28160 13820 28212
rect 13872 28200 13878 28212
rect 14461 28203 14519 28209
rect 14461 28200 14473 28203
rect 13872 28172 14473 28200
rect 13872 28160 13878 28172
rect 14461 28169 14473 28172
rect 14507 28169 14519 28203
rect 14461 28163 14519 28169
rect 15838 28160 15844 28212
rect 15896 28200 15902 28212
rect 20530 28200 20536 28212
rect 15896 28172 20536 28200
rect 15896 28160 15902 28172
rect 20530 28160 20536 28172
rect 20588 28160 20594 28212
rect 23198 28160 23204 28212
rect 23256 28200 23262 28212
rect 23566 28200 23572 28212
rect 23256 28172 23572 28200
rect 23256 28160 23262 28172
rect 23566 28160 23572 28172
rect 23624 28160 23630 28212
rect 24026 28200 24032 28212
rect 23987 28172 24032 28200
rect 24026 28160 24032 28172
rect 24084 28160 24090 28212
rect 25041 28203 25099 28209
rect 25041 28169 25053 28203
rect 25087 28200 25099 28203
rect 25590 28200 25596 28212
rect 25087 28172 25596 28200
rect 25087 28169 25099 28172
rect 25041 28163 25099 28169
rect 25590 28160 25596 28172
rect 25648 28160 25654 28212
rect 28442 28160 28448 28212
rect 28500 28200 28506 28212
rect 28626 28200 28632 28212
rect 28500 28172 28632 28200
rect 28500 28160 28506 28172
rect 28626 28160 28632 28172
rect 28684 28200 28690 28212
rect 29362 28200 29368 28212
rect 28684 28172 29224 28200
rect 29323 28172 29368 28200
rect 28684 28160 28690 28172
rect 13173 28135 13231 28141
rect 13173 28101 13185 28135
rect 13219 28132 13231 28135
rect 13538 28132 13544 28144
rect 13219 28104 13544 28132
rect 13219 28101 13231 28104
rect 13173 28095 13231 28101
rect 13538 28092 13544 28104
rect 13596 28092 13602 28144
rect 15933 28135 15991 28141
rect 15933 28101 15945 28135
rect 15979 28132 15991 28135
rect 16482 28132 16488 28144
rect 15979 28104 16488 28132
rect 15979 28101 15991 28104
rect 15933 28095 15991 28101
rect 16482 28092 16488 28104
rect 16540 28092 16546 28144
rect 20162 28132 20168 28144
rect 18432 28104 20168 28132
rect 15654 28024 15660 28076
rect 15712 28064 15718 28076
rect 18432 28073 18460 28104
rect 20162 28092 20168 28104
rect 20220 28092 20226 28144
rect 23106 28092 23112 28144
rect 23164 28132 23170 28144
rect 24673 28135 24731 28141
rect 24673 28132 24685 28135
rect 23164 28104 24685 28132
rect 23164 28092 23170 28104
rect 24673 28101 24685 28104
rect 24719 28101 24731 28135
rect 24673 28095 24731 28101
rect 24765 28135 24823 28141
rect 24765 28101 24777 28135
rect 24811 28132 24823 28135
rect 26786 28132 26792 28144
rect 24811 28104 26792 28132
rect 24811 28101 24823 28104
rect 24765 28095 24823 28101
rect 26786 28092 26792 28104
rect 26844 28092 26850 28144
rect 27246 28092 27252 28144
rect 27304 28132 27310 28144
rect 27304 28104 28948 28132
rect 27304 28092 27310 28104
rect 16025 28067 16083 28073
rect 16025 28064 16037 28067
rect 15712 28036 16037 28064
rect 15712 28024 15718 28036
rect 16025 28033 16037 28036
rect 16071 28033 16083 28067
rect 16025 28027 16083 28033
rect 18417 28067 18475 28073
rect 18417 28033 18429 28067
rect 18463 28033 18475 28067
rect 18417 28027 18475 28033
rect 18684 28067 18742 28073
rect 18684 28033 18696 28067
rect 18730 28064 18742 28067
rect 19518 28064 19524 28076
rect 18730 28036 19524 28064
rect 18730 28033 18742 28036
rect 18684 28027 18742 28033
rect 19518 28024 19524 28036
rect 19576 28024 19582 28076
rect 21913 28067 21971 28073
rect 21913 28033 21925 28067
rect 21959 28064 21971 28067
rect 22002 28064 22008 28076
rect 21959 28036 22008 28064
rect 21959 28033 21971 28036
rect 21913 28027 21971 28033
rect 22002 28024 22008 28036
rect 22060 28024 22066 28076
rect 22462 28024 22468 28076
rect 22520 28064 22526 28076
rect 22649 28067 22707 28073
rect 22649 28064 22661 28067
rect 22520 28036 22661 28064
rect 22520 28024 22526 28036
rect 22649 28033 22661 28036
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 22916 28067 22974 28073
rect 22916 28033 22928 28067
rect 22962 28064 22974 28067
rect 23198 28064 23204 28076
rect 22962 28036 23204 28064
rect 22962 28033 22974 28036
rect 22916 28027 22974 28033
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 23842 28024 23848 28076
rect 23900 28064 23906 28076
rect 24489 28067 24547 28073
rect 24489 28064 24501 28067
rect 23900 28036 24501 28064
rect 23900 28024 23906 28036
rect 24489 28033 24501 28036
rect 24535 28033 24547 28067
rect 24489 28027 24547 28033
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28064 24915 28067
rect 25130 28064 25136 28076
rect 24903 28036 25136 28064
rect 24903 28033 24915 28036
rect 24857 28027 24915 28033
rect 25130 28024 25136 28036
rect 25188 28024 25194 28076
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28033 27583 28067
rect 27525 28027 27583 28033
rect 15746 27956 15752 28008
rect 15804 27996 15810 28008
rect 15841 27999 15899 28005
rect 15841 27996 15853 27999
rect 15804 27968 15853 27996
rect 15804 27956 15810 27968
rect 15841 27965 15853 27968
rect 15887 27965 15899 27999
rect 27540 27996 27568 28027
rect 28442 28024 28448 28076
rect 28500 28064 28506 28076
rect 28537 28067 28595 28073
rect 28537 28064 28549 28067
rect 28500 28036 28549 28064
rect 28500 28024 28506 28036
rect 28537 28033 28549 28036
rect 28583 28033 28595 28067
rect 28537 28027 28595 28033
rect 28629 28067 28687 28073
rect 28629 28033 28641 28067
rect 28675 28033 28687 28067
rect 28629 28027 28687 28033
rect 28721 28067 28779 28073
rect 28721 28033 28733 28067
rect 28767 28064 28779 28067
rect 28810 28064 28816 28076
rect 28767 28036 28816 28064
rect 28767 28033 28779 28036
rect 28721 28027 28779 28033
rect 28261 27999 28319 28005
rect 28261 27996 28273 27999
rect 27540 27968 28273 27996
rect 15841 27959 15899 27965
rect 28261 27965 28273 27968
rect 28307 27965 28319 27999
rect 28261 27959 28319 27965
rect 15470 27928 15476 27940
rect 15431 27900 15476 27928
rect 15470 27888 15476 27900
rect 15528 27888 15534 27940
rect 27706 27928 27712 27940
rect 27667 27900 27712 27928
rect 27706 27888 27712 27900
rect 27764 27888 27770 27940
rect 18322 27820 18328 27872
rect 18380 27860 18386 27872
rect 19426 27860 19432 27872
rect 18380 27832 19432 27860
rect 18380 27820 18386 27832
rect 19426 27820 19432 27832
rect 19484 27860 19490 27872
rect 19797 27863 19855 27869
rect 19797 27860 19809 27863
rect 19484 27832 19809 27860
rect 19484 27820 19490 27832
rect 19797 27829 19809 27832
rect 19843 27829 19855 27863
rect 19797 27823 19855 27829
rect 22097 27863 22155 27869
rect 22097 27829 22109 27863
rect 22143 27860 22155 27863
rect 23566 27860 23572 27872
rect 22143 27832 23572 27860
rect 22143 27829 22155 27832
rect 22097 27823 22155 27829
rect 23566 27820 23572 27832
rect 23624 27820 23630 27872
rect 28644 27860 28672 28027
rect 28810 28024 28816 28036
rect 28868 28024 28874 28076
rect 28920 28073 28948 28104
rect 28905 28067 28963 28073
rect 28905 28033 28917 28067
rect 28951 28033 28963 28067
rect 28905 28027 28963 28033
rect 29196 27928 29224 28172
rect 29362 28160 29368 28172
rect 29420 28160 29426 28212
rect 29454 28160 29460 28212
rect 29512 28200 29518 28212
rect 29512 28172 29960 28200
rect 29512 28160 29518 28172
rect 29288 28104 29776 28132
rect 29288 27996 29316 28104
rect 29748 28073 29776 28104
rect 29641 28067 29699 28073
rect 29641 28064 29653 28067
rect 29472 28036 29653 28064
rect 29362 27996 29368 28008
rect 29288 27968 29368 27996
rect 29362 27956 29368 27968
rect 29420 27956 29426 28008
rect 29472 27928 29500 28036
rect 29641 28033 29653 28036
rect 29687 28033 29699 28067
rect 29641 28027 29699 28033
rect 29733 28067 29791 28073
rect 29733 28033 29745 28067
rect 29779 28033 29791 28067
rect 29733 28027 29791 28033
rect 29825 28067 29883 28073
rect 29825 28033 29837 28067
rect 29871 28033 29883 28067
rect 29932 28064 29960 28172
rect 30009 28067 30067 28073
rect 30009 28064 30021 28067
rect 29932 28036 30021 28064
rect 29825 28027 29883 28033
rect 30009 28033 30021 28036
rect 30055 28033 30067 28067
rect 30009 28027 30067 28033
rect 29546 27956 29552 28008
rect 29604 27996 29610 28008
rect 29840 27996 29868 28027
rect 29604 27968 29868 27996
rect 29604 27956 29610 27968
rect 29196 27900 29500 27928
rect 31478 27860 31484 27872
rect 28644 27832 31484 27860
rect 31478 27820 31484 27832
rect 31536 27820 31542 27872
rect 1104 27770 30820 27792
rect 1104 27718 5915 27770
rect 5967 27718 5979 27770
rect 6031 27718 6043 27770
rect 6095 27718 6107 27770
rect 6159 27718 6171 27770
rect 6223 27718 15846 27770
rect 15898 27718 15910 27770
rect 15962 27718 15974 27770
rect 16026 27718 16038 27770
rect 16090 27718 16102 27770
rect 16154 27718 25776 27770
rect 25828 27718 25840 27770
rect 25892 27718 25904 27770
rect 25956 27718 25968 27770
rect 26020 27718 26032 27770
rect 26084 27718 30820 27770
rect 1104 27696 30820 27718
rect 15378 27616 15384 27668
rect 15436 27656 15442 27668
rect 16393 27659 16451 27665
rect 16393 27656 16405 27659
rect 15436 27628 16405 27656
rect 15436 27616 15442 27628
rect 16393 27625 16405 27628
rect 16439 27625 16451 27659
rect 21542 27656 21548 27668
rect 21503 27628 21548 27656
rect 16393 27619 16451 27625
rect 21542 27616 21548 27628
rect 21600 27616 21606 27668
rect 26694 27656 26700 27668
rect 26528 27628 26700 27656
rect 14553 27591 14611 27597
rect 14553 27557 14565 27591
rect 14599 27557 14611 27591
rect 14553 27551 14611 27557
rect 17037 27591 17095 27597
rect 17037 27557 17049 27591
rect 17083 27557 17095 27591
rect 17037 27551 17095 27557
rect 25317 27591 25375 27597
rect 25317 27557 25329 27591
rect 25363 27588 25375 27591
rect 25406 27588 25412 27600
rect 25363 27560 25412 27588
rect 25363 27557 25375 27560
rect 25317 27551 25375 27557
rect 14568 27520 14596 27551
rect 15013 27523 15071 27529
rect 15013 27520 15025 27523
rect 14568 27492 15025 27520
rect 15013 27489 15025 27492
rect 15059 27489 15071 27523
rect 15013 27483 15071 27489
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 12066 27452 12072 27464
rect 12027 27424 12072 27452
rect 12066 27412 12072 27424
rect 12124 27412 12130 27464
rect 12342 27461 12348 27464
rect 12336 27452 12348 27461
rect 12303 27424 12348 27452
rect 12336 27415 12348 27424
rect 12342 27412 12348 27415
rect 12400 27412 12406 27464
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27452 14427 27455
rect 17052 27452 17080 27551
rect 25406 27548 25412 27560
rect 25464 27548 25470 27600
rect 25774 27548 25780 27600
rect 25832 27588 25838 27600
rect 26528 27588 26556 27628
rect 26694 27616 26700 27628
rect 26752 27616 26758 27668
rect 28074 27588 28080 27600
rect 25832 27560 26556 27588
rect 27540 27560 28080 27588
rect 25832 27548 25838 27560
rect 21545 27523 21603 27529
rect 21545 27489 21557 27523
rect 21591 27520 21603 27523
rect 21818 27520 21824 27532
rect 21591 27492 21824 27520
rect 21591 27489 21603 27492
rect 21545 27483 21603 27489
rect 21818 27480 21824 27492
rect 21876 27480 21882 27532
rect 25148 27492 26096 27520
rect 25148 27464 25176 27492
rect 21634 27452 21640 27464
rect 14415 27424 17080 27452
rect 21595 27424 21640 27452
rect 14415 27421 14427 27424
rect 14369 27415 14427 27421
rect 21634 27412 21640 27424
rect 21692 27412 21698 27464
rect 24578 27412 24584 27464
rect 24636 27452 24642 27464
rect 24765 27455 24823 27461
rect 24765 27452 24777 27455
rect 24636 27424 24777 27452
rect 24636 27412 24642 27424
rect 24765 27421 24777 27424
rect 24811 27421 24823 27455
rect 25130 27452 25136 27464
rect 25043 27424 25136 27452
rect 24765 27415 24823 27421
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25406 27412 25412 27464
rect 25464 27452 25470 27464
rect 25774 27452 25780 27464
rect 25464 27424 25780 27452
rect 25464 27412 25470 27424
rect 25774 27412 25780 27424
rect 25832 27412 25838 27464
rect 26068 27461 26096 27492
rect 26510 27480 26516 27532
rect 26568 27520 26574 27532
rect 26694 27520 26700 27532
rect 26568 27492 26700 27520
rect 26568 27480 26574 27492
rect 26694 27480 26700 27492
rect 26752 27480 26758 27532
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27452 26111 27455
rect 26142 27452 26148 27464
rect 26099 27424 26148 27452
rect 26099 27421 26111 27424
rect 26053 27415 26111 27421
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 27430 27452 27436 27464
rect 27391 27424 27436 27452
rect 27430 27412 27436 27424
rect 27488 27412 27494 27464
rect 27540 27452 27568 27560
rect 28074 27548 28080 27560
rect 28132 27548 28138 27600
rect 29454 27548 29460 27600
rect 29512 27588 29518 27600
rect 30101 27591 30159 27597
rect 30101 27588 30113 27591
rect 29512 27560 30113 27588
rect 29512 27548 29518 27560
rect 30101 27557 30113 27560
rect 30147 27557 30159 27591
rect 30101 27551 30159 27557
rect 31478 27548 31484 27600
rect 31536 27588 31542 27600
rect 31754 27588 31760 27600
rect 31536 27560 31760 27588
rect 31536 27548 31542 27560
rect 31754 27548 31760 27560
rect 31812 27548 31818 27600
rect 27706 27520 27712 27532
rect 27667 27492 27712 27520
rect 27706 27480 27712 27492
rect 27764 27480 27770 27532
rect 27801 27523 27859 27529
rect 27801 27489 27813 27523
rect 27847 27520 27859 27523
rect 28258 27520 28264 27532
rect 27847 27492 28264 27520
rect 27847 27489 27859 27492
rect 27801 27483 27859 27489
rect 28258 27480 28264 27492
rect 28316 27480 28322 27532
rect 27617 27455 27675 27461
rect 27617 27452 27629 27455
rect 27540 27424 27629 27452
rect 27617 27421 27629 27424
rect 27663 27421 27675 27455
rect 27617 27415 27675 27421
rect 27996 27455 28054 27461
rect 27996 27421 28008 27455
rect 28042 27421 28054 27455
rect 27996 27415 28054 27421
rect 15286 27393 15292 27396
rect 15280 27384 15292 27393
rect 15247 27356 15292 27384
rect 15280 27347 15292 27356
rect 15286 27344 15292 27347
rect 15344 27344 15350 27396
rect 15746 27344 15752 27396
rect 15804 27384 15810 27396
rect 16942 27384 16948 27396
rect 15804 27356 16948 27384
rect 15804 27344 15810 27356
rect 16942 27344 16948 27356
rect 17000 27384 17006 27396
rect 17313 27387 17371 27393
rect 17313 27384 17325 27387
rect 17000 27356 17325 27384
rect 17000 27344 17006 27356
rect 17313 27353 17325 27356
rect 17359 27353 17371 27387
rect 17586 27384 17592 27396
rect 17547 27356 17592 27384
rect 17313 27347 17371 27353
rect 17586 27344 17592 27356
rect 17644 27344 17650 27396
rect 21361 27387 21419 27393
rect 21361 27353 21373 27387
rect 21407 27384 21419 27387
rect 21450 27384 21456 27396
rect 21407 27356 21456 27384
rect 21407 27353 21419 27356
rect 21361 27347 21419 27353
rect 21450 27344 21456 27356
rect 21508 27384 21514 27396
rect 21910 27384 21916 27396
rect 21508 27356 21916 27384
rect 21508 27344 21514 27356
rect 21910 27344 21916 27356
rect 21968 27344 21974 27396
rect 24670 27344 24676 27396
rect 24728 27384 24734 27396
rect 24949 27387 25007 27393
rect 24949 27384 24961 27387
rect 24728 27356 24961 27384
rect 24728 27344 24734 27356
rect 24949 27353 24961 27356
rect 24995 27353 25007 27387
rect 24949 27347 25007 27353
rect 25041 27387 25099 27393
rect 25041 27353 25053 27387
rect 25087 27384 25099 27387
rect 26510 27384 26516 27396
rect 25087 27356 26516 27384
rect 25087 27353 25099 27356
rect 25041 27347 25099 27353
rect 26510 27344 26516 27356
rect 26568 27344 26574 27396
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 12802 27276 12808 27328
rect 12860 27316 12866 27328
rect 13449 27319 13507 27325
rect 13449 27316 13461 27319
rect 12860 27288 13461 27316
rect 12860 27276 12866 27288
rect 13449 27285 13461 27288
rect 13495 27285 13507 27319
rect 13449 27279 13507 27285
rect 16482 27276 16488 27328
rect 16540 27316 16546 27328
rect 17497 27319 17555 27325
rect 17497 27316 17509 27319
rect 16540 27288 17509 27316
rect 16540 27276 16546 27288
rect 17497 27285 17509 27288
rect 17543 27285 17555 27319
rect 17497 27279 17555 27285
rect 21821 27319 21879 27325
rect 21821 27285 21833 27319
rect 21867 27316 21879 27319
rect 22002 27316 22008 27328
rect 21867 27288 22008 27316
rect 21867 27285 21879 27288
rect 21821 27279 21879 27285
rect 22002 27276 22008 27288
rect 22060 27276 22066 27328
rect 22370 27276 22376 27328
rect 22428 27316 22434 27328
rect 22554 27316 22560 27328
rect 22428 27288 22560 27316
rect 22428 27276 22434 27288
rect 22554 27276 22560 27288
rect 22612 27276 22618 27328
rect 24210 27276 24216 27328
rect 24268 27316 24274 27328
rect 24578 27316 24584 27328
rect 24268 27288 24584 27316
rect 24268 27276 24274 27288
rect 24578 27276 24584 27288
rect 24636 27276 24642 27328
rect 27522 27276 27528 27328
rect 27580 27316 27586 27328
rect 28000 27316 28028 27415
rect 28442 27412 28448 27464
rect 28500 27452 28506 27464
rect 28721 27455 28779 27461
rect 28721 27452 28733 27455
rect 28500 27424 28733 27452
rect 28500 27412 28506 27424
rect 28721 27421 28733 27424
rect 28767 27421 28779 27455
rect 28721 27415 28779 27421
rect 28902 27412 28908 27464
rect 28960 27452 28966 27464
rect 29917 27455 29975 27461
rect 29917 27452 29929 27455
rect 28960 27424 29929 27452
rect 28960 27412 28966 27424
rect 29917 27421 29929 27424
rect 29963 27421 29975 27455
rect 29917 27415 29975 27421
rect 31018 27412 31024 27464
rect 31076 27452 31082 27464
rect 31754 27452 31760 27464
rect 31076 27424 31760 27452
rect 31076 27412 31082 27424
rect 31754 27412 31760 27424
rect 31812 27412 31818 27464
rect 28920 27384 28948 27412
rect 28092 27356 28948 27384
rect 28092 27328 28120 27356
rect 29362 27344 29368 27396
rect 29420 27384 29426 27396
rect 29733 27387 29791 27393
rect 29733 27384 29745 27387
rect 29420 27356 29745 27384
rect 29420 27344 29426 27356
rect 29733 27353 29745 27356
rect 29779 27353 29791 27387
rect 29733 27347 29791 27353
rect 27580 27288 28028 27316
rect 27580 27276 27586 27288
rect 28074 27276 28080 27328
rect 28132 27276 28138 27328
rect 28169 27319 28227 27325
rect 28169 27285 28181 27319
rect 28215 27316 28227 27319
rect 28442 27316 28448 27328
rect 28215 27288 28448 27316
rect 28215 27285 28227 27288
rect 28169 27279 28227 27285
rect 28442 27276 28448 27288
rect 28500 27276 28506 27328
rect 28902 27316 28908 27328
rect 28863 27288 28908 27316
rect 28902 27276 28908 27288
rect 28960 27276 28966 27328
rect 1104 27226 30820 27248
rect 1104 27174 10880 27226
rect 10932 27174 10944 27226
rect 10996 27174 11008 27226
rect 11060 27174 11072 27226
rect 11124 27174 11136 27226
rect 11188 27174 20811 27226
rect 20863 27174 20875 27226
rect 20927 27174 20939 27226
rect 20991 27174 21003 27226
rect 21055 27174 21067 27226
rect 21119 27174 30820 27226
rect 1104 27152 30820 27174
rect 2133 27115 2191 27121
rect 2133 27081 2145 27115
rect 2179 27081 2191 27115
rect 2133 27075 2191 27081
rect 1397 26979 1455 26985
rect 1397 26945 1409 26979
rect 1443 26976 1455 26979
rect 2148 26976 2176 27075
rect 2314 27072 2320 27124
rect 2372 27112 2378 27124
rect 2372 27084 6914 27112
rect 2372 27072 2378 27084
rect 6886 27044 6914 27084
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 12529 27115 12587 27121
rect 12529 27112 12541 27115
rect 12124 27084 12541 27112
rect 12124 27072 12130 27084
rect 12529 27081 12541 27084
rect 12575 27081 12587 27115
rect 15657 27115 15715 27121
rect 12529 27075 12587 27081
rect 13464 27084 15424 27112
rect 13464 27044 13492 27084
rect 6886 27016 13492 27044
rect 13541 27047 13599 27053
rect 13541 27013 13553 27047
rect 13587 27044 13599 27047
rect 15010 27044 15016 27056
rect 13587 27016 15016 27044
rect 13587 27013 13599 27016
rect 13541 27007 13599 27013
rect 15010 27004 15016 27016
rect 15068 27004 15074 27056
rect 1443 26948 2176 26976
rect 2317 26979 2375 26985
rect 1443 26945 1455 26948
rect 1397 26939 1455 26945
rect 2317 26945 2329 26979
rect 2363 26976 2375 26979
rect 12345 26979 12403 26985
rect 2363 26948 6914 26976
rect 2363 26945 2375 26948
rect 2317 26939 2375 26945
rect 6886 26908 6914 26948
rect 12345 26945 12357 26979
rect 12391 26976 12403 26979
rect 12526 26976 12532 26988
rect 12391 26948 12532 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 12526 26936 12532 26948
rect 12584 26936 12590 26988
rect 14461 26979 14519 26985
rect 14461 26945 14473 26979
rect 14507 26976 14519 26979
rect 15179 26979 15237 26985
rect 15179 26976 15191 26979
rect 14507 26948 15191 26976
rect 14507 26945 14519 26948
rect 14461 26939 14519 26945
rect 15179 26945 15191 26948
rect 15225 26945 15237 26979
rect 15396 26976 15424 27084
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16482 27112 16488 27124
rect 15703 27084 16488 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16482 27072 16488 27084
rect 16540 27072 16546 27124
rect 22278 27072 22284 27124
rect 22336 27112 22342 27124
rect 22554 27112 22560 27124
rect 22336 27084 22560 27112
rect 22336 27072 22342 27084
rect 22554 27072 22560 27084
rect 22612 27072 22618 27124
rect 23198 27112 23204 27124
rect 23159 27084 23204 27112
rect 23198 27072 23204 27084
rect 23256 27072 23262 27124
rect 24946 27112 24952 27124
rect 24907 27084 24952 27112
rect 24946 27072 24952 27084
rect 25004 27072 25010 27124
rect 25409 27115 25467 27121
rect 25409 27081 25421 27115
rect 25455 27112 25467 27115
rect 26234 27112 26240 27124
rect 25455 27084 26240 27112
rect 25455 27081 25467 27084
rect 25409 27075 25467 27081
rect 26234 27072 26240 27084
rect 26292 27072 26298 27124
rect 27338 27072 27344 27124
rect 27396 27112 27402 27124
rect 27525 27115 27583 27121
rect 27525 27112 27537 27115
rect 27396 27084 27537 27112
rect 27396 27072 27402 27084
rect 27525 27081 27537 27084
rect 27571 27112 27583 27115
rect 27985 27115 28043 27121
rect 27985 27112 27997 27115
rect 27571 27084 27997 27112
rect 27571 27081 27583 27084
rect 27525 27075 27583 27081
rect 27985 27081 27997 27084
rect 28031 27081 28043 27115
rect 27985 27075 28043 27081
rect 28721 27115 28779 27121
rect 28721 27081 28733 27115
rect 28767 27112 28779 27115
rect 29178 27112 29184 27124
rect 28767 27084 29184 27112
rect 28767 27081 28779 27084
rect 28721 27075 28779 27081
rect 29178 27072 29184 27084
rect 29236 27072 29242 27124
rect 29454 27072 29460 27124
rect 29512 27112 29518 27124
rect 29917 27115 29975 27121
rect 29917 27112 29929 27115
rect 29512 27084 29929 27112
rect 29512 27072 29518 27084
rect 29917 27081 29929 27084
rect 29963 27112 29975 27115
rect 30834 27112 30840 27124
rect 29963 27084 30840 27112
rect 29963 27081 29975 27084
rect 29917 27075 29975 27081
rect 30834 27072 30840 27084
rect 30892 27072 30898 27124
rect 15473 27047 15531 27053
rect 15473 27013 15485 27047
rect 15519 27044 15531 27047
rect 15746 27044 15752 27056
rect 15519 27016 15752 27044
rect 15519 27013 15531 27016
rect 15473 27007 15531 27013
rect 15746 27004 15752 27016
rect 15804 27004 15810 27056
rect 18874 27044 18880 27056
rect 18835 27016 18880 27044
rect 18874 27004 18880 27016
rect 18932 27004 18938 27056
rect 24302 27004 24308 27056
rect 24360 27044 24366 27056
rect 24581 27047 24639 27053
rect 24581 27044 24593 27047
rect 24360 27016 24593 27044
rect 24360 27004 24366 27016
rect 24581 27013 24593 27016
rect 24627 27013 24639 27047
rect 24581 27007 24639 27013
rect 24673 27047 24731 27053
rect 24673 27013 24685 27047
rect 24719 27044 24731 27047
rect 24719 27016 25452 27044
rect 24719 27013 24731 27016
rect 24673 27007 24731 27013
rect 25424 26988 25452 27016
rect 25590 27004 25596 27056
rect 25648 27044 25654 27056
rect 25866 27044 25872 27056
rect 25648 27016 25872 27044
rect 25648 27004 25654 27016
rect 25866 27004 25872 27016
rect 25924 27044 25930 27056
rect 26053 27047 26111 27053
rect 26053 27044 26065 27047
rect 25924 27016 26065 27044
rect 25924 27004 25930 27016
rect 26053 27013 26065 27016
rect 26099 27013 26111 27047
rect 26053 27007 26111 27013
rect 27246 27004 27252 27056
rect 27304 27044 27310 27056
rect 27430 27044 27436 27056
rect 27304 27016 27436 27044
rect 27304 27004 27310 27016
rect 27430 27004 27436 27016
rect 27488 27004 27494 27056
rect 28074 27004 28080 27056
rect 28132 27044 28138 27056
rect 28537 27047 28595 27053
rect 28537 27044 28549 27047
rect 28132 27016 28549 27044
rect 28132 27004 28138 27016
rect 28537 27013 28549 27016
rect 28583 27013 28595 27047
rect 28537 27007 28595 27013
rect 22278 26976 22284 26988
rect 15396 26948 22094 26976
rect 22239 26948 22284 26976
rect 15179 26939 15237 26945
rect 6886 26880 15700 26908
rect 15672 26840 15700 26880
rect 15746 26868 15752 26920
rect 15804 26908 15810 26920
rect 17586 26908 17592 26920
rect 15804 26880 17592 26908
rect 15804 26868 15810 26880
rect 17586 26868 17592 26880
rect 17644 26868 17650 26920
rect 22066 26908 22094 26948
rect 22278 26936 22284 26948
rect 22336 26936 22342 26988
rect 23382 26976 23388 26988
rect 23343 26948 23388 26976
rect 23382 26936 23388 26948
rect 23440 26936 23446 26988
rect 23661 26979 23719 26985
rect 23661 26945 23673 26979
rect 23707 26976 23719 26979
rect 24026 26976 24032 26988
rect 23707 26948 24032 26976
rect 23707 26945 23719 26948
rect 23661 26939 23719 26945
rect 24026 26936 24032 26948
rect 24084 26936 24090 26988
rect 24394 26976 24400 26988
rect 24355 26948 24400 26976
rect 24394 26936 24400 26948
rect 24452 26936 24458 26988
rect 24765 26979 24823 26985
rect 24765 26945 24777 26979
rect 24811 26976 24823 26979
rect 25130 26976 25136 26988
rect 24811 26948 25136 26976
rect 24811 26945 24823 26948
rect 24765 26939 24823 26945
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 25406 26936 25412 26988
rect 25464 26936 25470 26988
rect 26329 26979 26387 26985
rect 26329 26945 26341 26979
rect 26375 26976 26387 26979
rect 27338 26976 27344 26988
rect 26375 26948 27344 26976
rect 26375 26945 26387 26948
rect 26329 26939 26387 26945
rect 27338 26936 27344 26948
rect 27396 26976 27402 26988
rect 27617 26979 27675 26985
rect 27617 26976 27629 26979
rect 27396 26948 27629 26976
rect 27396 26936 27402 26948
rect 27617 26945 27629 26948
rect 27663 26945 27675 26979
rect 28353 26979 28411 26985
rect 28353 26976 28365 26979
rect 27617 26939 27675 26945
rect 28000 26948 28365 26976
rect 22066 26880 26188 26908
rect 22462 26840 22468 26852
rect 15672 26812 22094 26840
rect 22423 26812 22468 26840
rect 1578 26772 1584 26784
rect 1539 26744 1584 26772
rect 1578 26732 1584 26744
rect 1636 26732 1642 26784
rect 13630 26772 13636 26784
rect 13591 26744 13636 26772
rect 13630 26732 13636 26744
rect 13688 26732 13694 26784
rect 14645 26775 14703 26781
rect 14645 26741 14657 26775
rect 14691 26772 14703 26775
rect 15654 26772 15660 26784
rect 14691 26744 15660 26772
rect 14691 26741 14703 26744
rect 14645 26735 14703 26741
rect 15654 26732 15660 26744
rect 15712 26732 15718 26784
rect 20162 26772 20168 26784
rect 20123 26744 20168 26772
rect 20162 26732 20168 26744
rect 20220 26732 20226 26784
rect 22066 26772 22094 26812
rect 22462 26800 22468 26812
rect 22520 26800 22526 26852
rect 25777 26843 25835 26849
rect 25777 26840 25789 26843
rect 22572 26812 25789 26840
rect 22572 26772 22600 26812
rect 25777 26809 25789 26812
rect 25823 26809 25835 26843
rect 25777 26803 25835 26809
rect 25866 26800 25872 26852
rect 25924 26800 25930 26852
rect 26050 26800 26056 26852
rect 26108 26800 26114 26852
rect 26160 26840 26188 26880
rect 26878 26868 26884 26920
rect 26936 26908 26942 26920
rect 27154 26908 27160 26920
rect 26936 26880 27160 26908
rect 26936 26868 26942 26880
rect 27154 26868 27160 26880
rect 27212 26868 27218 26920
rect 27430 26908 27436 26920
rect 27391 26880 27436 26908
rect 27430 26868 27436 26880
rect 27488 26868 27494 26920
rect 27065 26843 27123 26849
rect 27065 26840 27077 26843
rect 26160 26812 27077 26840
rect 27065 26809 27077 26812
rect 27111 26809 27123 26843
rect 27065 26803 27123 26809
rect 28000 26840 28028 26948
rect 28353 26945 28365 26948
rect 28399 26945 28411 26979
rect 28353 26939 28411 26945
rect 29089 26979 29147 26985
rect 29089 26945 29101 26979
rect 29135 26976 29147 26979
rect 29454 26976 29460 26988
rect 29135 26948 29460 26976
rect 29135 26945 29147 26948
rect 29089 26939 29147 26945
rect 29454 26936 29460 26948
rect 29512 26936 29518 26988
rect 29825 26911 29883 26917
rect 29825 26908 29837 26911
rect 28644 26880 29837 26908
rect 28644 26840 28672 26880
rect 29825 26877 29837 26880
rect 29871 26877 29883 26911
rect 30006 26908 30012 26920
rect 29967 26880 30012 26908
rect 29825 26871 29883 26877
rect 30006 26868 30012 26880
rect 30064 26868 30070 26920
rect 30558 26868 30564 26920
rect 30616 26908 30622 26920
rect 30926 26908 30932 26920
rect 30616 26880 30932 26908
rect 30616 26868 30622 26880
rect 30926 26868 30932 26880
rect 30984 26868 30990 26920
rect 28000 26812 28672 26840
rect 22066 26744 22600 26772
rect 23569 26775 23627 26781
rect 23569 26741 23581 26775
rect 23615 26772 23627 26775
rect 23658 26772 23664 26784
rect 23615 26744 23664 26772
rect 23615 26741 23627 26744
rect 23569 26735 23627 26741
rect 23658 26732 23664 26744
rect 23716 26732 23722 26784
rect 24854 26732 24860 26784
rect 24912 26772 24918 26784
rect 25884 26772 25912 26800
rect 24912 26744 25912 26772
rect 26068 26772 26096 26800
rect 26234 26772 26240 26784
rect 26068 26744 26240 26772
rect 24912 26732 24918 26744
rect 26234 26732 26240 26744
rect 26292 26732 26298 26784
rect 26878 26732 26884 26784
rect 26936 26772 26942 26784
rect 28000 26772 28028 26812
rect 29178 26800 29184 26852
rect 29236 26840 29242 26852
rect 30374 26840 30380 26852
rect 29236 26812 30380 26840
rect 29236 26800 29242 26812
rect 30374 26800 30380 26812
rect 30432 26800 30438 26852
rect 29454 26772 29460 26784
rect 26936 26744 28028 26772
rect 29415 26744 29460 26772
rect 26936 26732 26942 26744
rect 29454 26732 29460 26744
rect 29512 26732 29518 26784
rect 1104 26682 30820 26704
rect 1104 26630 5915 26682
rect 5967 26630 5979 26682
rect 6031 26630 6043 26682
rect 6095 26630 6107 26682
rect 6159 26630 6171 26682
rect 6223 26630 15846 26682
rect 15898 26630 15910 26682
rect 15962 26630 15974 26682
rect 16026 26630 16038 26682
rect 16090 26630 16102 26682
rect 16154 26630 25776 26682
rect 25828 26630 25840 26682
rect 25892 26630 25904 26682
rect 25956 26630 25968 26682
rect 26020 26630 26032 26682
rect 26084 26630 30820 26682
rect 1104 26608 30820 26630
rect 15562 26528 15568 26580
rect 15620 26568 15626 26580
rect 17037 26571 17095 26577
rect 17037 26568 17049 26571
rect 15620 26540 17049 26568
rect 15620 26528 15626 26540
rect 17037 26537 17049 26540
rect 17083 26537 17095 26571
rect 17037 26531 17095 26537
rect 18046 26528 18052 26580
rect 18104 26568 18110 26580
rect 29454 26568 29460 26580
rect 18104 26540 29460 26568
rect 18104 26528 18110 26540
rect 29454 26528 29460 26540
rect 29512 26528 29518 26580
rect 29914 26528 29920 26580
rect 29972 26568 29978 26580
rect 30101 26571 30159 26577
rect 30101 26568 30113 26571
rect 29972 26540 30113 26568
rect 29972 26528 29978 26540
rect 30101 26537 30113 26540
rect 30147 26537 30159 26571
rect 30101 26531 30159 26537
rect 2133 26503 2191 26509
rect 2133 26469 2145 26503
rect 2179 26469 2191 26503
rect 2133 26463 2191 26469
rect 25869 26503 25927 26509
rect 25869 26469 25881 26503
rect 25915 26500 25927 26503
rect 27430 26500 27436 26512
rect 25915 26472 27436 26500
rect 25915 26469 25927 26472
rect 25869 26463 25927 26469
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26364 1455 26367
rect 2148 26364 2176 26463
rect 27430 26460 27436 26472
rect 27488 26460 27494 26512
rect 28074 26500 28080 26512
rect 28035 26472 28080 26500
rect 28074 26460 28080 26472
rect 28132 26460 28138 26512
rect 28902 26500 28908 26512
rect 28863 26472 28908 26500
rect 28902 26460 28908 26472
rect 28960 26460 28966 26512
rect 31386 26500 31392 26512
rect 29656 26472 31392 26500
rect 15654 26432 15660 26444
rect 15615 26404 15660 26432
rect 15654 26392 15660 26404
rect 15712 26392 15718 26444
rect 29656 26432 29684 26472
rect 31386 26460 31392 26472
rect 31444 26460 31450 26512
rect 28736 26404 29684 26432
rect 2314 26364 2320 26376
rect 1443 26336 2176 26364
rect 2275 26336 2320 26364
rect 1443 26333 1455 26336
rect 1397 26327 1455 26333
rect 2314 26324 2320 26336
rect 2372 26324 2378 26376
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26364 13231 26367
rect 13814 26364 13820 26376
rect 13219 26336 13820 26364
rect 13219 26333 13231 26336
rect 13173 26327 13231 26333
rect 13814 26324 13820 26336
rect 13872 26324 13878 26376
rect 15194 26324 15200 26376
rect 15252 26364 15258 26376
rect 15913 26367 15971 26373
rect 15913 26364 15925 26367
rect 15252 26336 15925 26364
rect 15252 26324 15258 26336
rect 15913 26333 15925 26336
rect 15959 26333 15971 26367
rect 15913 26327 15971 26333
rect 22922 26324 22928 26376
rect 22980 26364 22986 26376
rect 25317 26367 25375 26373
rect 25317 26364 25329 26367
rect 22980 26336 25329 26364
rect 22980 26324 22986 26336
rect 25317 26333 25329 26336
rect 25363 26333 25375 26367
rect 25317 26327 25375 26333
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26364 25743 26367
rect 26142 26364 26148 26376
rect 25731 26336 26148 26364
rect 25731 26333 25743 26336
rect 25685 26327 25743 26333
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 26234 26324 26240 26376
rect 26292 26364 26298 26376
rect 27706 26364 27712 26376
rect 26292 26336 27712 26364
rect 26292 26324 26298 26336
rect 27706 26324 27712 26336
rect 27764 26364 27770 26376
rect 28736 26373 28764 26404
rect 28261 26367 28319 26373
rect 28261 26364 28273 26367
rect 27764 26336 28273 26364
rect 27764 26324 27770 26336
rect 28261 26333 28273 26336
rect 28307 26333 28319 26367
rect 28261 26327 28319 26333
rect 28721 26367 28779 26373
rect 28721 26333 28733 26367
rect 28767 26333 28779 26367
rect 28721 26327 28779 26333
rect 29733 26367 29791 26373
rect 29733 26333 29745 26367
rect 29779 26364 29791 26367
rect 30374 26364 30380 26376
rect 29779 26336 30380 26364
rect 29779 26333 29791 26336
rect 29733 26327 29791 26333
rect 30374 26324 30380 26336
rect 30432 26324 30438 26376
rect 25498 26296 25504 26308
rect 25459 26268 25504 26296
rect 25498 26256 25504 26268
rect 25556 26256 25562 26308
rect 25593 26299 25651 26305
rect 25593 26265 25605 26299
rect 25639 26296 25651 26299
rect 27430 26296 27436 26308
rect 25639 26268 27436 26296
rect 25639 26265 25651 26268
rect 25593 26259 25651 26265
rect 27430 26256 27436 26268
rect 27488 26256 27494 26308
rect 28074 26256 28080 26308
rect 28132 26296 28138 26308
rect 29917 26299 29975 26305
rect 29917 26296 29929 26299
rect 28132 26268 29929 26296
rect 28132 26256 28138 26268
rect 29917 26265 29929 26268
rect 29963 26265 29975 26299
rect 29917 26259 29975 26265
rect 1578 26228 1584 26240
rect 1539 26200 1584 26228
rect 1578 26188 1584 26200
rect 1636 26188 1642 26240
rect 12986 26188 12992 26240
rect 13044 26228 13050 26240
rect 13265 26231 13323 26237
rect 13265 26228 13277 26231
rect 13044 26200 13277 26228
rect 13044 26188 13050 26200
rect 13265 26197 13277 26200
rect 13311 26197 13323 26231
rect 13265 26191 13323 26197
rect 1104 26138 30820 26160
rect 1104 26086 10880 26138
rect 10932 26086 10944 26138
rect 10996 26086 11008 26138
rect 11060 26086 11072 26138
rect 11124 26086 11136 26138
rect 11188 26086 20811 26138
rect 20863 26086 20875 26138
rect 20927 26086 20939 26138
rect 20991 26086 21003 26138
rect 21055 26086 21067 26138
rect 21119 26086 30820 26138
rect 1104 26064 30820 26086
rect 12989 26027 13047 26033
rect 12989 25993 13001 26027
rect 13035 26024 13047 26027
rect 13262 26024 13268 26036
rect 13035 25996 13268 26024
rect 13035 25993 13047 25996
rect 12989 25987 13047 25993
rect 13262 25984 13268 25996
rect 13320 26024 13326 26036
rect 13630 26024 13636 26036
rect 13320 25996 13636 26024
rect 13320 25984 13326 25996
rect 13630 25984 13636 25996
rect 13688 25984 13694 26036
rect 22370 25984 22376 26036
rect 22428 26024 22434 26036
rect 22922 26024 22928 26036
rect 22428 25996 22928 26024
rect 22428 25984 22434 25996
rect 22922 25984 22928 25996
rect 22980 25984 22986 26036
rect 23842 25984 23848 26036
rect 23900 26024 23906 26036
rect 24118 26024 24124 26036
rect 23900 25996 24124 26024
rect 23900 25984 23906 25996
rect 24118 25984 24124 25996
rect 24176 25984 24182 26036
rect 26694 25984 26700 26036
rect 26752 26024 26758 26036
rect 28169 26027 28227 26033
rect 28169 26024 28181 26027
rect 26752 25996 28181 26024
rect 26752 25984 26758 25996
rect 28169 25993 28181 25996
rect 28215 25993 28227 26027
rect 28626 26024 28632 26036
rect 28587 25996 28632 26024
rect 28169 25987 28227 25993
rect 28626 25984 28632 25996
rect 28684 25984 28690 26036
rect 29086 26024 29092 26036
rect 29047 25996 29092 26024
rect 29086 25984 29092 25996
rect 29144 26024 29150 26036
rect 29917 26027 29975 26033
rect 29917 26024 29929 26027
rect 29144 25996 29929 26024
rect 29144 25984 29150 25996
rect 29917 25993 29929 25996
rect 29963 25993 29975 26027
rect 29917 25987 29975 25993
rect 18046 25956 18052 25968
rect 6886 25928 18052 25956
rect 1397 25891 1455 25897
rect 1397 25857 1409 25891
rect 1443 25888 1455 25891
rect 2317 25891 2375 25897
rect 1443 25860 2176 25888
rect 1443 25857 1455 25860
rect 1397 25851 1455 25857
rect 2148 25761 2176 25860
rect 2317 25857 2329 25891
rect 2363 25888 2375 25891
rect 6886 25888 6914 25928
rect 18046 25916 18052 25928
rect 18104 25916 18110 25968
rect 18601 25959 18659 25965
rect 18601 25925 18613 25959
rect 18647 25956 18659 25959
rect 20162 25956 20168 25968
rect 18647 25928 20168 25956
rect 18647 25925 18659 25928
rect 18601 25919 18659 25925
rect 20162 25916 20168 25928
rect 20220 25916 20226 25968
rect 22646 25956 22652 25968
rect 22480 25928 22652 25956
rect 13078 25888 13084 25900
rect 2363 25860 6914 25888
rect 13039 25860 13084 25888
rect 2363 25857 2375 25860
rect 2317 25851 2375 25857
rect 13078 25848 13084 25860
rect 13136 25848 13142 25900
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25857 17923 25891
rect 19334 25888 19340 25900
rect 19295 25860 19340 25888
rect 17865 25851 17923 25857
rect 12986 25820 12992 25832
rect 12947 25792 12992 25820
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 17880 25820 17908 25851
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 22370 25848 22376 25900
rect 22428 25888 22434 25900
rect 22480 25897 22508 25928
rect 22646 25916 22652 25928
rect 22704 25916 22710 25968
rect 27338 25916 27344 25968
rect 27396 25956 27402 25968
rect 29454 25956 29460 25968
rect 27396 25928 29460 25956
rect 27396 25916 27402 25928
rect 29454 25916 29460 25928
rect 29512 25956 29518 25968
rect 30006 25956 30012 25968
rect 29512 25928 30012 25956
rect 29512 25916 29518 25928
rect 30006 25916 30012 25928
rect 30064 25916 30070 25968
rect 22465 25891 22523 25897
rect 22465 25888 22477 25891
rect 22428 25860 22477 25888
rect 22428 25848 22434 25860
rect 22465 25857 22477 25860
rect 22511 25857 22523 25891
rect 22465 25851 22523 25857
rect 22557 25891 22615 25897
rect 22557 25857 22569 25891
rect 22603 25857 22615 25891
rect 22738 25888 22744 25900
rect 22699 25860 22744 25888
rect 22557 25851 22615 25857
rect 18506 25820 18512 25832
rect 17880 25792 18512 25820
rect 18506 25780 18512 25792
rect 18564 25820 18570 25832
rect 18785 25823 18843 25829
rect 18785 25820 18797 25823
rect 18564 25792 18797 25820
rect 18564 25780 18570 25792
rect 18785 25789 18797 25792
rect 18831 25789 18843 25823
rect 22572 25820 22600 25851
rect 22738 25848 22744 25860
rect 22796 25848 22802 25900
rect 22833 25891 22891 25897
rect 22833 25857 22845 25891
rect 22879 25888 22891 25891
rect 24118 25888 24124 25900
rect 22879 25860 24124 25888
rect 22879 25857 22891 25860
rect 22833 25851 22891 25857
rect 24118 25848 24124 25860
rect 24176 25848 24182 25900
rect 27798 25888 27804 25900
rect 27759 25860 27804 25888
rect 27798 25848 27804 25860
rect 27856 25848 27862 25900
rect 27985 25891 28043 25897
rect 27985 25857 27997 25891
rect 28031 25888 28043 25891
rect 28074 25888 28080 25900
rect 28031 25860 28080 25888
rect 28031 25857 28043 25860
rect 27985 25851 28043 25857
rect 28074 25848 28080 25860
rect 28132 25848 28138 25900
rect 28442 25888 28448 25900
rect 28403 25860 28448 25888
rect 28442 25848 28448 25860
rect 28500 25848 28506 25900
rect 24026 25820 24032 25832
rect 22572 25792 24032 25820
rect 18785 25783 18843 25789
rect 24026 25780 24032 25792
rect 24084 25780 24090 25832
rect 29362 25780 29368 25832
rect 29420 25820 29426 25832
rect 29917 25823 29975 25829
rect 29917 25820 29929 25823
rect 29420 25792 29929 25820
rect 29420 25780 29426 25792
rect 29917 25789 29929 25792
rect 29963 25789 29975 25823
rect 29917 25783 29975 25789
rect 2133 25755 2191 25761
rect 2133 25721 2145 25755
rect 2179 25721 2191 25755
rect 12526 25752 12532 25764
rect 12487 25724 12532 25752
rect 2133 25715 2191 25721
rect 12526 25712 12532 25724
rect 12584 25712 12590 25764
rect 24394 25712 24400 25764
rect 24452 25752 24458 25764
rect 29457 25755 29515 25761
rect 29457 25752 29469 25755
rect 24452 25724 29469 25752
rect 24452 25712 24458 25724
rect 29457 25721 29469 25724
rect 29503 25721 29515 25755
rect 29932 25752 29960 25783
rect 30558 25752 30564 25764
rect 29932 25724 30564 25752
rect 29457 25715 29515 25721
rect 30558 25712 30564 25724
rect 30616 25712 30622 25764
rect 1578 25684 1584 25696
rect 1539 25656 1584 25684
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 17862 25644 17868 25696
rect 17920 25684 17926 25696
rect 17957 25687 18015 25693
rect 17957 25684 17969 25687
rect 17920 25656 17969 25684
rect 17920 25644 17926 25656
rect 17957 25653 17969 25656
rect 18003 25653 18015 25687
rect 17957 25647 18015 25653
rect 19521 25687 19579 25693
rect 19521 25653 19533 25687
rect 19567 25684 19579 25687
rect 19610 25684 19616 25696
rect 19567 25656 19616 25684
rect 19567 25653 19579 25656
rect 19521 25647 19579 25653
rect 19610 25644 19616 25656
rect 19668 25644 19674 25696
rect 21450 25644 21456 25696
rect 21508 25684 21514 25696
rect 22281 25687 22339 25693
rect 22281 25684 22293 25687
rect 21508 25656 22293 25684
rect 21508 25644 21514 25656
rect 22281 25653 22293 25656
rect 22327 25653 22339 25687
rect 22281 25647 22339 25653
rect 1104 25594 30820 25616
rect 1104 25542 5915 25594
rect 5967 25542 5979 25594
rect 6031 25542 6043 25594
rect 6095 25542 6107 25594
rect 6159 25542 6171 25594
rect 6223 25542 15846 25594
rect 15898 25542 15910 25594
rect 15962 25542 15974 25594
rect 16026 25542 16038 25594
rect 16090 25542 16102 25594
rect 16154 25542 25776 25594
rect 25828 25542 25840 25594
rect 25892 25542 25904 25594
rect 25956 25542 25968 25594
rect 26020 25542 26032 25594
rect 26084 25542 30820 25594
rect 1104 25520 30820 25542
rect 1670 25480 1676 25492
rect 1631 25452 1676 25480
rect 1670 25440 1676 25452
rect 1728 25440 1734 25492
rect 2314 25440 2320 25492
rect 2372 25480 2378 25492
rect 24394 25480 24400 25492
rect 2372 25452 24400 25480
rect 2372 25440 2378 25452
rect 24394 25440 24400 25452
rect 24452 25440 24458 25492
rect 24489 25483 24547 25489
rect 24489 25449 24501 25483
rect 24535 25480 24547 25483
rect 25498 25480 25504 25492
rect 24535 25452 25504 25480
rect 24535 25449 24547 25452
rect 24489 25443 24547 25449
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 27338 25440 27344 25492
rect 27396 25480 27402 25492
rect 27433 25483 27491 25489
rect 27433 25480 27445 25483
rect 27396 25452 27445 25480
rect 27396 25440 27402 25452
rect 27433 25449 27445 25452
rect 27479 25449 27491 25483
rect 27433 25443 27491 25449
rect 28166 25440 28172 25492
rect 28224 25480 28230 25492
rect 28353 25483 28411 25489
rect 28353 25480 28365 25483
rect 28224 25452 28365 25480
rect 28224 25440 28230 25452
rect 28353 25449 28365 25452
rect 28399 25449 28411 25483
rect 30006 25480 30012 25492
rect 29967 25452 30012 25480
rect 28353 25443 28411 25449
rect 30006 25440 30012 25452
rect 30064 25440 30070 25492
rect 16850 25372 16856 25424
rect 16908 25412 16914 25424
rect 17405 25415 17463 25421
rect 17405 25412 17417 25415
rect 16908 25384 17417 25412
rect 16908 25372 16914 25384
rect 17405 25381 17417 25384
rect 17451 25381 17463 25415
rect 17405 25375 17463 25381
rect 20993 25415 21051 25421
rect 20993 25381 21005 25415
rect 21039 25412 21051 25415
rect 21818 25412 21824 25424
rect 21039 25384 21824 25412
rect 21039 25381 21051 25384
rect 20993 25375 21051 25381
rect 21818 25372 21824 25384
rect 21876 25372 21882 25424
rect 27614 25372 27620 25424
rect 27672 25412 27678 25424
rect 28813 25415 28871 25421
rect 28813 25412 28825 25415
rect 27672 25384 28825 25412
rect 27672 25372 27678 25384
rect 17957 25347 18015 25353
rect 17957 25313 17969 25347
rect 18003 25344 18015 25347
rect 18322 25344 18328 25356
rect 18003 25316 18328 25344
rect 18003 25313 18015 25316
rect 17957 25307 18015 25313
rect 18322 25304 18328 25316
rect 18380 25304 18386 25356
rect 19610 25344 19616 25356
rect 19571 25316 19616 25344
rect 19610 25304 19616 25316
rect 19668 25304 19674 25356
rect 22922 25344 22928 25356
rect 22480 25316 22928 25344
rect 1854 25276 1860 25288
rect 1815 25248 1860 25276
rect 1854 25236 1860 25248
rect 1912 25236 1918 25288
rect 16390 25276 16396 25288
rect 16351 25248 16396 25276
rect 16390 25236 16396 25248
rect 16448 25236 16454 25288
rect 18506 25276 18512 25288
rect 18467 25248 18512 25276
rect 18506 25236 18512 25248
rect 18564 25236 18570 25288
rect 22370 25276 22376 25288
rect 22331 25248 22376 25276
rect 22370 25236 22376 25248
rect 22428 25236 22434 25288
rect 22480 25285 22508 25316
rect 22922 25304 22928 25316
rect 22980 25304 22986 25356
rect 24394 25304 24400 25356
rect 24452 25344 24458 25356
rect 24949 25347 25007 25353
rect 24949 25344 24961 25347
rect 24452 25316 24961 25344
rect 24452 25304 24458 25316
rect 24949 25313 24961 25316
rect 24995 25313 25007 25347
rect 24949 25307 25007 25313
rect 26326 25304 26332 25356
rect 26384 25344 26390 25356
rect 27338 25344 27344 25356
rect 26384 25316 27344 25344
rect 26384 25304 26390 25316
rect 27338 25304 27344 25316
rect 27396 25304 27402 25356
rect 22465 25279 22523 25285
rect 22465 25245 22477 25279
rect 22511 25245 22523 25279
rect 22646 25276 22652 25288
rect 22607 25248 22652 25276
rect 22465 25239 22523 25245
rect 17678 25208 17684 25220
rect 17639 25180 17684 25208
rect 17678 25168 17684 25180
rect 17736 25168 17742 25220
rect 17862 25208 17868 25220
rect 17823 25180 17868 25208
rect 17862 25168 17868 25180
rect 17920 25168 17926 25220
rect 19880 25211 19938 25217
rect 19880 25177 19892 25211
rect 19926 25208 19938 25211
rect 20622 25208 20628 25220
rect 19926 25180 20628 25208
rect 19926 25177 19938 25180
rect 19880 25171 19938 25177
rect 20622 25168 20628 25180
rect 20680 25168 20686 25220
rect 16574 25140 16580 25152
rect 16535 25112 16580 25140
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 18046 25100 18052 25152
rect 18104 25140 18110 25152
rect 18601 25143 18659 25149
rect 18601 25140 18613 25143
rect 18104 25112 18613 25140
rect 18104 25100 18110 25112
rect 18601 25109 18613 25112
rect 18647 25109 18659 25143
rect 18601 25103 18659 25109
rect 21266 25100 21272 25152
rect 21324 25140 21330 25152
rect 22189 25143 22247 25149
rect 22189 25140 22201 25143
rect 21324 25112 22201 25140
rect 21324 25100 21330 25112
rect 22189 25109 22201 25112
rect 22235 25109 22247 25143
rect 22189 25103 22247 25109
rect 22370 25100 22376 25152
rect 22428 25140 22434 25152
rect 22480 25140 22508 25239
rect 22646 25236 22652 25248
rect 22704 25236 22710 25288
rect 22738 25236 22744 25288
rect 22796 25276 22802 25288
rect 22796 25248 22841 25276
rect 22796 25236 22802 25248
rect 23934 25236 23940 25288
rect 23992 25276 23998 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 23992 25248 24685 25276
rect 23992 25236 23998 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24854 25276 24860 25288
rect 24815 25248 24860 25276
rect 24673 25239 24731 25245
rect 24688 25208 24716 25239
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25276 25559 25279
rect 26513 25279 26571 25285
rect 26513 25276 26525 25279
rect 25547 25248 26525 25276
rect 25547 25245 25559 25248
rect 25501 25239 25559 25245
rect 26513 25245 26525 25248
rect 26559 25276 26571 25279
rect 26694 25276 26700 25288
rect 26559 25248 26700 25276
rect 26559 25245 26571 25248
rect 26513 25239 26571 25245
rect 26694 25236 26700 25248
rect 26752 25276 26758 25288
rect 28074 25276 28080 25288
rect 26752 25248 28080 25276
rect 26752 25236 26758 25248
rect 28074 25236 28080 25248
rect 28132 25276 28138 25288
rect 28169 25279 28227 25285
rect 28169 25276 28181 25279
rect 28132 25248 28181 25276
rect 28132 25236 28138 25248
rect 28169 25245 28181 25248
rect 28215 25245 28227 25279
rect 28169 25239 28227 25245
rect 25685 25211 25743 25217
rect 25685 25208 25697 25211
rect 24688 25180 25697 25208
rect 25685 25177 25697 25180
rect 25731 25177 25743 25211
rect 25685 25171 25743 25177
rect 27341 25211 27399 25217
rect 27341 25177 27353 25211
rect 27387 25208 27399 25211
rect 27614 25208 27620 25220
rect 27387 25180 27620 25208
rect 27387 25177 27399 25180
rect 27341 25171 27399 25177
rect 27614 25168 27620 25180
rect 27672 25168 27678 25220
rect 27985 25211 28043 25217
rect 27985 25177 27997 25211
rect 28031 25208 28043 25211
rect 28276 25208 28304 25384
rect 28813 25381 28825 25384
rect 28859 25381 28871 25415
rect 28813 25375 28871 25381
rect 28994 25372 29000 25424
rect 29052 25412 29058 25424
rect 29362 25412 29368 25424
rect 29052 25384 29368 25412
rect 29052 25372 29058 25384
rect 29362 25372 29368 25384
rect 29420 25372 29426 25424
rect 28994 25276 29000 25288
rect 28955 25248 29000 25276
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 29825 25279 29883 25285
rect 29825 25245 29837 25279
rect 29871 25276 29883 25279
rect 30834 25276 30840 25288
rect 29871 25248 30840 25276
rect 29871 25245 29883 25248
rect 29825 25239 29883 25245
rect 30834 25236 30840 25248
rect 30892 25236 30898 25288
rect 28031 25180 28304 25208
rect 28031 25177 28043 25180
rect 27985 25171 28043 25177
rect 22428 25112 22508 25140
rect 22428 25100 22434 25112
rect 26326 25100 26332 25152
rect 26384 25140 26390 25152
rect 26697 25143 26755 25149
rect 26697 25140 26709 25143
rect 26384 25112 26709 25140
rect 26384 25100 26390 25112
rect 26697 25109 26709 25112
rect 26743 25140 26755 25143
rect 27522 25140 27528 25152
rect 26743 25112 27528 25140
rect 26743 25109 26755 25112
rect 26697 25103 26755 25109
rect 27522 25100 27528 25112
rect 27580 25100 27586 25152
rect 1104 25050 30820 25072
rect 1104 24998 10880 25050
rect 10932 24998 10944 25050
rect 10996 24998 11008 25050
rect 11060 24998 11072 25050
rect 11124 24998 11136 25050
rect 11188 24998 20811 25050
rect 20863 24998 20875 25050
rect 20927 24998 20939 25050
rect 20991 24998 21003 25050
rect 21055 24998 21067 25050
rect 21119 24998 30820 25050
rect 1104 24976 30820 24998
rect 13262 24936 13268 24948
rect 13223 24908 13268 24936
rect 13262 24896 13268 24908
rect 13320 24896 13326 24948
rect 20622 24936 20628 24948
rect 14476 24908 19334 24936
rect 20583 24908 20628 24936
rect 1854 24828 1860 24880
rect 1912 24868 1918 24880
rect 1912 24840 9674 24868
rect 1912 24828 1918 24840
rect 1397 24803 1455 24809
rect 1397 24769 1409 24803
rect 1443 24800 1455 24803
rect 2314 24800 2320 24812
rect 1443 24772 2176 24800
rect 2275 24772 2320 24800
rect 1443 24769 1455 24772
rect 1397 24763 1455 24769
rect 1578 24664 1584 24676
rect 1539 24636 1584 24664
rect 1578 24624 1584 24636
rect 1636 24624 1642 24676
rect 2148 24673 2176 24772
rect 2314 24760 2320 24772
rect 2372 24760 2378 24812
rect 9646 24800 9674 24840
rect 12986 24828 12992 24880
rect 13044 24868 13050 24880
rect 13081 24871 13139 24877
rect 13081 24868 13093 24871
rect 13044 24840 13093 24868
rect 13044 24828 13050 24840
rect 13081 24837 13093 24840
rect 13127 24837 13139 24871
rect 14476 24868 14504 24908
rect 18598 24868 18604 24880
rect 13081 24831 13139 24837
rect 13188 24840 14504 24868
rect 17420 24840 18604 24868
rect 13188 24800 13216 24840
rect 9646 24772 13216 24800
rect 13998 24760 14004 24812
rect 14056 24800 14062 24812
rect 14165 24803 14223 24809
rect 14165 24800 14177 24803
rect 14056 24772 14177 24800
rect 14056 24760 14062 24772
rect 14165 24769 14177 24772
rect 14211 24769 14223 24803
rect 14165 24763 14223 24769
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24769 17187 24803
rect 17129 24763 17187 24769
rect 17221 24806 17279 24812
rect 17221 24772 17233 24806
rect 17267 24772 17279 24806
rect 17221 24766 17279 24772
rect 17334 24803 17392 24809
rect 17334 24769 17346 24803
rect 17380 24800 17392 24803
rect 17420 24800 17448 24840
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 19306 24868 19334 24908
rect 20622 24896 20628 24908
rect 20680 24896 20686 24948
rect 21836 24908 23612 24936
rect 21836 24868 21864 24908
rect 19306 24840 21864 24868
rect 17380 24772 17448 24800
rect 17380 24769 17392 24772
rect 13078 24692 13084 24744
rect 13136 24732 13142 24744
rect 13357 24735 13415 24741
rect 13357 24732 13369 24735
rect 13136 24704 13369 24732
rect 13136 24692 13142 24704
rect 13357 24701 13369 24704
rect 13403 24732 13415 24735
rect 13446 24732 13452 24744
rect 13403 24704 13452 24732
rect 13403 24701 13415 24704
rect 13357 24695 13415 24701
rect 13446 24692 13452 24704
rect 13504 24692 13510 24744
rect 13906 24732 13912 24744
rect 13867 24704 13912 24732
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 2133 24667 2191 24673
rect 2133 24633 2145 24667
rect 2179 24633 2191 24667
rect 2133 24627 2191 24633
rect 15289 24667 15347 24673
rect 15289 24633 15301 24667
rect 15335 24664 15347 24667
rect 15378 24664 15384 24676
rect 15335 24636 15384 24664
rect 15335 24633 15347 24636
rect 15289 24627 15347 24633
rect 15378 24624 15384 24636
rect 15436 24624 15442 24676
rect 12805 24599 12863 24605
rect 12805 24565 12817 24599
rect 12851 24596 12863 24599
rect 14090 24596 14096 24608
rect 12851 24568 14096 24596
rect 12851 24565 12863 24568
rect 12805 24559 12863 24565
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 16853 24599 16911 24605
rect 16853 24565 16865 24599
rect 16899 24596 16911 24599
rect 16942 24596 16948 24608
rect 16899 24568 16948 24596
rect 16899 24565 16911 24568
rect 16853 24559 16911 24565
rect 16942 24556 16948 24568
rect 17000 24556 17006 24608
rect 17144 24596 17172 24763
rect 17236 24732 17264 24766
rect 17334 24763 17392 24769
rect 17494 24760 17500 24812
rect 17552 24800 17558 24812
rect 17957 24803 18015 24809
rect 17552 24772 17597 24800
rect 17552 24760 17558 24772
rect 17957 24769 17969 24803
rect 18003 24800 18015 24803
rect 18046 24800 18052 24812
rect 18003 24772 18052 24800
rect 18003 24769 18015 24772
rect 17957 24763 18015 24769
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18224 24803 18282 24809
rect 18224 24769 18236 24803
rect 18270 24800 18282 24803
rect 19242 24800 19248 24812
rect 18270 24772 19248 24800
rect 18270 24769 18282 24772
rect 18224 24763 18282 24769
rect 19242 24760 19248 24772
rect 19300 24760 19306 24812
rect 20901 24803 20959 24809
rect 20901 24769 20913 24803
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 20993 24803 21051 24809
rect 20993 24769 21005 24803
rect 21039 24769 21051 24803
rect 20993 24763 21051 24769
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21266 24800 21272 24812
rect 21227 24772 21272 24800
rect 21085 24763 21143 24769
rect 17862 24732 17868 24744
rect 17236 24704 17868 24732
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 18138 24596 18144 24608
rect 17144 24568 18144 24596
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 19337 24599 19395 24605
rect 19337 24565 19349 24599
rect 19383 24596 19395 24599
rect 19518 24596 19524 24608
rect 19383 24568 19524 24596
rect 19383 24565 19395 24568
rect 19337 24559 19395 24565
rect 19518 24556 19524 24568
rect 19576 24556 19582 24608
rect 20916 24596 20944 24763
rect 21008 24664 21036 24763
rect 21100 24732 21128 24763
rect 21266 24760 21272 24772
rect 21324 24760 21330 24812
rect 22094 24800 22100 24812
rect 21560 24772 22100 24800
rect 21560 24732 21588 24772
rect 22094 24760 22100 24772
rect 22152 24760 22158 24812
rect 22922 24760 22928 24812
rect 22980 24800 22986 24812
rect 23109 24803 23167 24809
rect 23109 24800 23121 24803
rect 22980 24772 23121 24800
rect 22980 24760 22986 24772
rect 23109 24769 23121 24772
rect 23155 24769 23167 24803
rect 23290 24800 23296 24812
rect 23251 24772 23296 24800
rect 23109 24763 23167 24769
rect 23290 24760 23296 24772
rect 23348 24760 23354 24812
rect 21818 24732 21824 24744
rect 21100 24704 21588 24732
rect 21779 24704 21824 24732
rect 21818 24692 21824 24704
rect 21876 24692 21882 24744
rect 22002 24692 22008 24744
rect 22060 24732 22066 24744
rect 22060 24692 22094 24732
rect 22646 24692 22652 24744
rect 22704 24732 22710 24744
rect 23385 24735 23443 24741
rect 23385 24732 23397 24735
rect 22704 24704 23397 24732
rect 22704 24692 22710 24704
rect 23385 24701 23397 24704
rect 23431 24701 23443 24735
rect 23385 24695 23443 24701
rect 23477 24735 23535 24741
rect 23477 24701 23489 24735
rect 23523 24701 23535 24735
rect 23477 24695 23535 24701
rect 21358 24664 21364 24676
rect 21008 24636 21364 24664
rect 21358 24624 21364 24636
rect 21416 24624 21422 24676
rect 22066 24664 22094 24692
rect 23492 24664 23520 24695
rect 22066 24636 23520 24664
rect 23584 24664 23612 24908
rect 23934 24896 23940 24948
rect 23992 24936 23998 24948
rect 26605 24939 26663 24945
rect 23992 24908 24716 24936
rect 23992 24896 23998 24908
rect 24688 24868 24716 24908
rect 26605 24905 26617 24939
rect 26651 24936 26663 24939
rect 26694 24936 26700 24948
rect 26651 24908 26700 24936
rect 26651 24905 26663 24908
rect 26605 24899 26663 24905
rect 26694 24896 26700 24908
rect 26752 24896 26758 24948
rect 28261 24939 28319 24945
rect 28261 24905 28273 24939
rect 28307 24936 28319 24939
rect 28902 24936 28908 24948
rect 28307 24908 28908 24936
rect 28307 24905 28319 24908
rect 28261 24899 28319 24905
rect 24688 24840 24808 24868
rect 23661 24803 23719 24809
rect 23661 24769 23673 24803
rect 23707 24769 23719 24803
rect 24302 24800 24308 24812
rect 24263 24772 24308 24800
rect 23661 24763 23719 24769
rect 23676 24732 23704 24763
rect 24302 24760 24308 24772
rect 24360 24760 24366 24812
rect 24780 24809 24808 24840
rect 27798 24828 27804 24880
rect 27856 24868 27862 24880
rect 28077 24871 28135 24877
rect 28077 24868 28089 24871
rect 27856 24840 28089 24868
rect 27856 24828 27862 24840
rect 28077 24837 28089 24840
rect 28123 24837 28135 24871
rect 28077 24831 28135 24837
rect 24489 24803 24547 24809
rect 24489 24769 24501 24803
rect 24535 24769 24547 24803
rect 24489 24763 24547 24769
rect 24765 24803 24823 24809
rect 24765 24769 24777 24803
rect 24811 24769 24823 24803
rect 24765 24763 24823 24769
rect 24394 24732 24400 24744
rect 23676 24704 24400 24732
rect 24394 24692 24400 24704
rect 24452 24692 24458 24744
rect 24504 24732 24532 24763
rect 26234 24760 26240 24812
rect 26292 24800 26298 24812
rect 26789 24803 26847 24809
rect 26789 24800 26801 24803
rect 26292 24772 26801 24800
rect 26292 24760 26298 24772
rect 26789 24769 26801 24772
rect 26835 24769 26847 24803
rect 26789 24763 26847 24769
rect 27433 24803 27491 24809
rect 27433 24769 27445 24803
rect 27479 24800 27491 24803
rect 28276 24800 28304 24899
rect 28902 24896 28908 24908
rect 28960 24896 28966 24948
rect 29086 24896 29092 24948
rect 29144 24936 29150 24948
rect 29917 24939 29975 24945
rect 29917 24936 29929 24939
rect 29144 24908 29929 24936
rect 29144 24896 29150 24908
rect 29917 24905 29929 24908
rect 29963 24905 29975 24939
rect 29917 24899 29975 24905
rect 27479 24772 28304 24800
rect 27479 24769 27491 24772
rect 27433 24763 27491 24769
rect 24578 24732 24584 24744
rect 24504 24704 24584 24732
rect 24578 24692 24584 24704
rect 24636 24692 24642 24744
rect 25314 24732 25320 24744
rect 25275 24704 25320 24732
rect 25314 24692 25320 24704
rect 25372 24692 25378 24744
rect 26804 24732 26832 24763
rect 29454 24760 29460 24812
rect 29512 24800 29518 24812
rect 30009 24803 30067 24809
rect 30009 24800 30021 24803
rect 29512 24772 30021 24800
rect 29512 24760 29518 24772
rect 30009 24769 30021 24772
rect 30055 24769 30067 24803
rect 30009 24763 30067 24769
rect 27614 24732 27620 24744
rect 26804 24704 27620 24732
rect 27614 24692 27620 24704
rect 27672 24692 27678 24744
rect 28353 24735 28411 24741
rect 28353 24701 28365 24735
rect 28399 24732 28411 24735
rect 29086 24732 29092 24744
rect 28399 24704 29092 24732
rect 28399 24701 28411 24704
rect 28353 24695 28411 24701
rect 29086 24692 29092 24704
rect 29144 24692 29150 24744
rect 29917 24735 29975 24741
rect 29917 24701 29929 24735
rect 29963 24732 29975 24735
rect 30374 24732 30380 24744
rect 29963 24704 30380 24732
rect 29963 24701 29975 24704
rect 29917 24695 29975 24701
rect 30374 24692 30380 24704
rect 30432 24692 30438 24744
rect 27801 24667 27859 24673
rect 27801 24664 27813 24667
rect 23584 24636 27813 24664
rect 27801 24633 27813 24636
rect 27847 24633 27859 24667
rect 27801 24627 27859 24633
rect 21266 24596 21272 24608
rect 20916 24568 21272 24596
rect 21266 24556 21272 24568
rect 21324 24596 21330 24608
rect 22051 24599 22109 24605
rect 22051 24596 22063 24599
rect 21324 24568 22063 24596
rect 21324 24556 21330 24568
rect 22051 24565 22063 24568
rect 22097 24565 22109 24599
rect 22051 24559 22109 24565
rect 22738 24556 22744 24608
rect 22796 24596 22802 24608
rect 23845 24599 23903 24605
rect 23845 24596 23857 24599
rect 22796 24568 23857 24596
rect 22796 24556 22802 24568
rect 23845 24565 23857 24568
rect 23891 24565 23903 24599
rect 23845 24559 23903 24565
rect 24673 24599 24731 24605
rect 24673 24565 24685 24599
rect 24719 24596 24731 24599
rect 24854 24596 24860 24608
rect 24719 24568 24860 24596
rect 24719 24565 24731 24568
rect 24673 24559 24731 24565
rect 24854 24556 24860 24568
rect 24912 24596 24918 24608
rect 25547 24599 25605 24605
rect 25547 24596 25559 24599
rect 24912 24568 25559 24596
rect 24912 24556 24918 24568
rect 25547 24565 25559 24568
rect 25593 24565 25605 24599
rect 25547 24559 25605 24565
rect 27338 24556 27344 24608
rect 27396 24596 27402 24608
rect 27982 24596 27988 24608
rect 27396 24568 27988 24596
rect 27396 24556 27402 24568
rect 27982 24556 27988 24568
rect 28040 24556 28046 24608
rect 28258 24556 28264 24608
rect 28316 24596 28322 24608
rect 28718 24596 28724 24608
rect 28316 24568 28724 24596
rect 28316 24556 28322 24568
rect 28718 24556 28724 24568
rect 28776 24556 28782 24608
rect 29454 24596 29460 24608
rect 29415 24568 29460 24596
rect 29454 24556 29460 24568
rect 29512 24556 29518 24608
rect 1104 24506 30820 24528
rect 1104 24454 5915 24506
rect 5967 24454 5979 24506
rect 6031 24454 6043 24506
rect 6095 24454 6107 24506
rect 6159 24454 6171 24506
rect 6223 24454 15846 24506
rect 15898 24454 15910 24506
rect 15962 24454 15974 24506
rect 16026 24454 16038 24506
rect 16090 24454 16102 24506
rect 16154 24454 25776 24506
rect 25828 24454 25840 24506
rect 25892 24454 25904 24506
rect 25956 24454 25968 24506
rect 26020 24454 26032 24506
rect 26084 24454 30820 24506
rect 1104 24432 30820 24454
rect 13906 24352 13912 24404
rect 13964 24392 13970 24404
rect 14277 24395 14335 24401
rect 14277 24392 14289 24395
rect 13964 24364 14289 24392
rect 13964 24352 13970 24364
rect 14277 24361 14289 24364
rect 14323 24361 14335 24395
rect 14277 24355 14335 24361
rect 14384 24364 17448 24392
rect 2133 24327 2191 24333
rect 2133 24293 2145 24327
rect 2179 24293 2191 24327
rect 2133 24287 2191 24293
rect 12897 24327 12955 24333
rect 12897 24293 12909 24327
rect 12943 24324 12955 24327
rect 13170 24324 13176 24336
rect 12943 24296 13176 24324
rect 12943 24293 12955 24296
rect 12897 24287 12955 24293
rect 1397 24191 1455 24197
rect 1397 24157 1409 24191
rect 1443 24188 1455 24191
rect 2148 24188 2176 24287
rect 13170 24284 13176 24296
rect 13228 24284 13234 24336
rect 14384 24256 14412 24364
rect 17420 24324 17448 24364
rect 17678 24352 17684 24404
rect 17736 24392 17742 24404
rect 17865 24395 17923 24401
rect 17865 24392 17877 24395
rect 17736 24364 17877 24392
rect 17736 24352 17742 24364
rect 17865 24361 17877 24364
rect 17911 24361 17923 24395
rect 19242 24392 19248 24404
rect 19203 24364 19248 24392
rect 17865 24355 17923 24361
rect 19242 24352 19248 24364
rect 19300 24352 19306 24404
rect 22278 24352 22284 24404
rect 22336 24392 22342 24404
rect 23293 24395 23351 24401
rect 23293 24392 23305 24395
rect 22336 24364 23305 24392
rect 22336 24352 22342 24364
rect 23293 24361 23305 24364
rect 23339 24361 23351 24395
rect 23293 24355 23351 24361
rect 24118 24352 24124 24404
rect 24176 24392 24182 24404
rect 24397 24395 24455 24401
rect 24397 24392 24409 24395
rect 24176 24364 24409 24392
rect 24176 24352 24182 24364
rect 24397 24361 24409 24364
rect 24443 24361 24455 24395
rect 24397 24355 24455 24361
rect 24596 24364 24808 24392
rect 24596 24324 24624 24364
rect 17420 24296 24624 24324
rect 24780 24324 24808 24364
rect 27338 24352 27344 24404
rect 27396 24392 27402 24404
rect 27522 24392 27528 24404
rect 27396 24364 27528 24392
rect 27396 24352 27402 24364
rect 27522 24352 27528 24364
rect 27580 24352 27586 24404
rect 27798 24352 27804 24404
rect 27856 24392 27862 24404
rect 28169 24395 28227 24401
rect 28169 24392 28181 24395
rect 27856 24364 28181 24392
rect 27856 24352 27862 24364
rect 28169 24361 28181 24364
rect 28215 24361 28227 24395
rect 28169 24355 28227 24361
rect 28626 24352 28632 24404
rect 28684 24392 28690 24404
rect 28813 24395 28871 24401
rect 28813 24392 28825 24395
rect 28684 24364 28825 24392
rect 28684 24352 28690 24364
rect 28813 24361 28825 24364
rect 28859 24361 28871 24395
rect 28813 24355 28871 24361
rect 28994 24352 29000 24404
rect 29052 24392 29058 24404
rect 29178 24392 29184 24404
rect 29052 24364 29184 24392
rect 29052 24352 29058 24364
rect 29178 24352 29184 24364
rect 29236 24352 29242 24404
rect 29454 24324 29460 24336
rect 24780 24296 29460 24324
rect 29454 24284 29460 24296
rect 29512 24284 29518 24336
rect 18966 24256 18972 24268
rect 12406 24228 14412 24256
rect 18524 24228 18972 24256
rect 1443 24160 2176 24188
rect 2317 24191 2375 24197
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 2317 24157 2329 24191
rect 2363 24188 2375 24191
rect 12406 24188 12434 24228
rect 18524 24200 18552 24228
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 22094 24256 22100 24268
rect 21284 24228 22100 24256
rect 2363 24160 12434 24188
rect 2363 24157 2375 24160
rect 2317 24151 2375 24157
rect 12986 24148 12992 24200
rect 13044 24188 13050 24200
rect 13173 24191 13231 24197
rect 13173 24188 13185 24191
rect 13044 24160 13185 24188
rect 13044 24148 13050 24160
rect 13173 24157 13185 24160
rect 13219 24157 13231 24191
rect 13446 24188 13452 24200
rect 13407 24160 13452 24188
rect 13173 24151 13231 24157
rect 13446 24148 13452 24160
rect 13504 24148 13510 24200
rect 14090 24188 14096 24200
rect 14051 24160 14096 24188
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24188 16543 24191
rect 16574 24188 16580 24200
rect 16531 24160 16580 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 18506 24188 18512 24200
rect 18419 24160 18512 24188
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 18647 24160 19441 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 19429 24157 19441 24160
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19518 24148 19524 24200
rect 19576 24188 19582 24200
rect 19705 24191 19763 24197
rect 19576 24160 19621 24188
rect 19576 24148 19582 24160
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 13262 24080 13268 24132
rect 13320 24120 13326 24132
rect 13357 24123 13415 24129
rect 13357 24120 13369 24123
rect 13320 24092 13369 24120
rect 13320 24080 13326 24092
rect 13357 24089 13369 24092
rect 13403 24089 13415 24123
rect 13357 24083 13415 24089
rect 16752 24123 16810 24129
rect 16752 24089 16764 24123
rect 16798 24120 16810 24123
rect 16942 24120 16948 24132
rect 16798 24092 16948 24120
rect 16798 24089 16810 24092
rect 16752 24083 16810 24089
rect 16942 24080 16948 24092
rect 17000 24080 17006 24132
rect 19610 24080 19616 24132
rect 19668 24120 19674 24132
rect 19720 24120 19748 24151
rect 19794 24148 19800 24200
rect 19852 24188 19858 24200
rect 21082 24188 21088 24200
rect 19852 24160 19897 24188
rect 21043 24160 21088 24188
rect 19852 24148 19858 24160
rect 21082 24148 21088 24160
rect 21140 24148 21146 24200
rect 21284 24197 21312 24228
rect 22094 24216 22100 24228
rect 22152 24216 22158 24268
rect 23842 24216 23848 24268
rect 23900 24256 23906 24268
rect 23900 24228 25544 24256
rect 23900 24216 23906 24228
rect 21177 24191 21235 24197
rect 21177 24157 21189 24191
rect 21223 24157 21235 24191
rect 21177 24151 21235 24157
rect 21269 24191 21327 24197
rect 21269 24157 21281 24191
rect 21315 24157 21327 24191
rect 21450 24188 21456 24200
rect 21411 24160 21456 24188
rect 21269 24151 21327 24157
rect 19668 24092 19748 24120
rect 21192 24120 21220 24151
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 22922 24148 22928 24200
rect 22980 24188 22986 24200
rect 22980 24160 23520 24188
rect 22980 24148 22986 24160
rect 21358 24120 21364 24132
rect 21192 24092 21364 24120
rect 19668 24080 19674 24092
rect 21358 24080 21364 24092
rect 21416 24080 21422 24132
rect 22002 24120 22008 24132
rect 21963 24092 22008 24120
rect 22002 24080 22008 24092
rect 22060 24080 22066 24132
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 20714 24012 20720 24064
rect 20772 24052 20778 24064
rect 20809 24055 20867 24061
rect 20809 24052 20821 24055
rect 20772 24024 20821 24052
rect 20772 24012 20778 24024
rect 20809 24021 20821 24024
rect 20855 24021 20867 24055
rect 20809 24015 20867 24021
rect 22186 24012 22192 24064
rect 22244 24052 22250 24064
rect 22738 24052 22744 24064
rect 22244 24024 22744 24052
rect 22244 24012 22250 24024
rect 22738 24012 22744 24024
rect 22796 24012 22802 24064
rect 23492 24052 23520 24160
rect 23934 24148 23940 24200
rect 23992 24188 23998 24200
rect 24653 24191 24711 24197
rect 24653 24188 24665 24191
rect 23992 24185 24348 24188
rect 23992 24182 24532 24185
rect 24596 24182 24665 24188
rect 23992 24160 24665 24182
rect 23992 24148 23998 24160
rect 24320 24157 24624 24160
rect 24504 24154 24624 24157
rect 24653 24157 24665 24160
rect 24699 24157 24711 24191
rect 24653 24151 24711 24157
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 24857 24191 24915 24197
rect 24857 24157 24869 24191
rect 24903 24157 24915 24191
rect 24857 24151 24915 24157
rect 25041 24191 25099 24197
rect 25041 24157 25053 24191
rect 25087 24188 25099 24191
rect 25406 24188 25412 24200
rect 25087 24160 25412 24188
rect 25087 24157 25099 24160
rect 25041 24151 25099 24157
rect 23566 24080 23572 24132
rect 23624 24120 23630 24132
rect 24780 24120 24808 24151
rect 23624 24092 24808 24120
rect 23624 24080 23630 24092
rect 24872 24052 24900 24151
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 25516 24120 25544 24228
rect 25593 24191 25651 24197
rect 25593 24157 25605 24191
rect 25639 24188 25651 24191
rect 26694 24188 26700 24200
rect 25639 24160 26700 24188
rect 25639 24157 25651 24160
rect 25593 24151 25651 24157
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 28350 24188 28356 24200
rect 28311 24160 28356 24188
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 28902 24148 28908 24200
rect 28960 24188 28966 24200
rect 28997 24191 29055 24197
rect 28997 24188 29009 24191
rect 28960 24160 29009 24188
rect 28960 24148 28966 24160
rect 28997 24157 29009 24160
rect 29043 24157 29055 24191
rect 28997 24151 29055 24157
rect 29914 24120 29920 24132
rect 25516 24092 26740 24120
rect 29875 24092 29920 24120
rect 26712 24064 26740 24092
rect 29914 24080 29920 24092
rect 29972 24080 29978 24132
rect 23492 24024 24900 24052
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 25685 24055 25743 24061
rect 25685 24052 25697 24055
rect 25004 24024 25697 24052
rect 25004 24012 25010 24024
rect 25685 24021 25697 24024
rect 25731 24021 25743 24055
rect 25685 24015 25743 24021
rect 26694 24012 26700 24064
rect 26752 24012 26758 24064
rect 27798 24012 27804 24064
rect 27856 24052 27862 24064
rect 30009 24055 30067 24061
rect 30009 24052 30021 24055
rect 27856 24024 30021 24052
rect 27856 24012 27862 24024
rect 30009 24021 30021 24024
rect 30055 24021 30067 24055
rect 30009 24015 30067 24021
rect 1104 23962 30820 23984
rect 1104 23910 10880 23962
rect 10932 23910 10944 23962
rect 10996 23910 11008 23962
rect 11060 23910 11072 23962
rect 11124 23910 11136 23962
rect 11188 23910 20811 23962
rect 20863 23910 20875 23962
rect 20927 23910 20939 23962
rect 20991 23910 21003 23962
rect 21055 23910 21067 23962
rect 21119 23910 30820 23962
rect 1104 23888 30820 23910
rect 10778 23808 10784 23860
rect 10836 23848 10842 23860
rect 14274 23848 14280 23860
rect 10836 23820 14280 23848
rect 10836 23808 10842 23820
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 17405 23851 17463 23857
rect 17405 23817 17417 23851
rect 17451 23848 17463 23851
rect 17494 23848 17500 23860
rect 17451 23820 17500 23848
rect 17451 23817 17463 23820
rect 17405 23811 17463 23817
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 17773 23851 17831 23857
rect 17773 23817 17785 23851
rect 17819 23848 17831 23851
rect 18138 23848 18144 23860
rect 17819 23820 18144 23848
rect 17819 23817 17831 23820
rect 17773 23811 17831 23817
rect 18138 23808 18144 23820
rect 18196 23808 18202 23860
rect 21177 23851 21235 23857
rect 21177 23817 21189 23851
rect 21223 23848 21235 23851
rect 22646 23848 22652 23860
rect 21223 23820 22652 23848
rect 21223 23817 21235 23820
rect 21177 23811 21235 23817
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 22741 23851 22799 23857
rect 22741 23817 22753 23851
rect 22787 23848 22799 23851
rect 22830 23848 22836 23860
rect 22787 23820 22836 23848
rect 22787 23817 22799 23820
rect 22741 23811 22799 23817
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 23106 23808 23112 23860
rect 23164 23848 23170 23860
rect 23385 23851 23443 23857
rect 23385 23848 23397 23851
rect 23164 23820 23397 23848
rect 23164 23808 23170 23820
rect 23385 23817 23397 23820
rect 23431 23817 23443 23851
rect 23385 23811 23443 23817
rect 24397 23851 24455 23857
rect 24397 23817 24409 23851
rect 24443 23848 24455 23851
rect 24670 23848 24676 23860
rect 24443 23820 24676 23848
rect 24443 23817 24455 23820
rect 24397 23811 24455 23817
rect 24670 23808 24676 23820
rect 24728 23808 24734 23860
rect 25406 23848 25412 23860
rect 25367 23820 25412 23848
rect 25406 23808 25412 23820
rect 25464 23808 25470 23860
rect 21192 23752 25360 23780
rect 21192 23724 21220 23752
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23712 1455 23715
rect 2317 23715 2375 23721
rect 1443 23684 2176 23712
rect 1443 23681 1455 23684
rect 1397 23675 1455 23681
rect 2148 23585 2176 23684
rect 2317 23681 2329 23715
rect 2363 23712 2375 23715
rect 12986 23712 12992 23724
rect 2363 23684 12992 23712
rect 2363 23681 2375 23684
rect 2317 23675 2375 23681
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13170 23712 13176 23724
rect 13131 23684 13176 23712
rect 13170 23672 13176 23684
rect 13228 23672 13234 23724
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23712 17647 23715
rect 17678 23712 17684 23724
rect 17635 23684 17684 23712
rect 17635 23681 17647 23684
rect 17589 23675 17647 23681
rect 17678 23672 17684 23684
rect 17736 23672 17742 23724
rect 17865 23715 17923 23721
rect 17865 23681 17877 23715
rect 17911 23712 17923 23715
rect 18506 23712 18512 23724
rect 17911 23684 18512 23712
rect 17911 23681 17923 23684
rect 17865 23675 17923 23681
rect 18506 23672 18512 23684
rect 18564 23672 18570 23724
rect 19150 23672 19156 23724
rect 19208 23712 19214 23724
rect 19521 23715 19579 23721
rect 19521 23712 19533 23715
rect 19208 23684 19533 23712
rect 19208 23672 19214 23684
rect 19521 23681 19533 23684
rect 19567 23681 19579 23715
rect 19521 23675 19579 23681
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21174 23712 21180 23724
rect 21131 23684 21180 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21174 23672 21180 23684
rect 21232 23672 21238 23724
rect 21266 23672 21272 23724
rect 21324 23712 21330 23724
rect 21324 23684 21369 23712
rect 21324 23672 21330 23684
rect 21910 23672 21916 23724
rect 21968 23712 21974 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21968 23684 22017 23712
rect 21968 23672 21974 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22186 23712 22192 23724
rect 22147 23684 22192 23712
rect 22005 23675 22063 23681
rect 22186 23672 22192 23684
rect 22244 23672 22250 23724
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23712 22615 23715
rect 22738 23712 22744 23724
rect 22603 23684 22744 23712
rect 22603 23681 22615 23684
rect 22557 23675 22615 23681
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 23569 23715 23627 23721
rect 23569 23681 23581 23715
rect 23615 23712 23627 23715
rect 24578 23712 24584 23724
rect 23615 23684 24584 23712
rect 23615 23681 23627 23684
rect 23569 23675 23627 23681
rect 24578 23672 24584 23684
rect 24636 23712 24642 23724
rect 24946 23712 24952 23724
rect 24636 23684 24952 23712
rect 24636 23672 24642 23684
rect 24946 23672 24952 23684
rect 25004 23672 25010 23724
rect 25332 23721 25360 23752
rect 27614 23740 27620 23792
rect 27672 23780 27678 23792
rect 27801 23783 27859 23789
rect 27801 23780 27813 23783
rect 27672 23752 27813 23780
rect 27672 23740 27678 23752
rect 27801 23749 27813 23752
rect 27847 23749 27859 23783
rect 27801 23743 27859 23749
rect 28442 23740 28448 23792
rect 28500 23780 28506 23792
rect 29917 23783 29975 23789
rect 29917 23780 29929 23783
rect 28500 23752 29929 23780
rect 28500 23740 28506 23752
rect 29917 23749 29929 23752
rect 29963 23749 29975 23783
rect 29917 23743 29975 23749
rect 25317 23715 25375 23721
rect 25317 23681 25329 23715
rect 25363 23681 25375 23715
rect 28626 23712 28632 23724
rect 28587 23684 28632 23712
rect 25317 23675 25375 23681
rect 28626 23672 28632 23684
rect 28684 23672 28690 23724
rect 29178 23712 29184 23724
rect 29139 23684 29184 23712
rect 29178 23672 29184 23684
rect 29236 23672 29242 23724
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 22152 23616 22293 23644
rect 22152 23604 22158 23616
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 22281 23607 22339 23613
rect 22373 23647 22431 23653
rect 22373 23613 22385 23647
rect 22419 23644 22431 23647
rect 23845 23647 23903 23653
rect 22419 23616 23060 23644
rect 22419 23613 22431 23616
rect 22373 23607 22431 23613
rect 2133 23579 2191 23585
rect 2133 23545 2145 23579
rect 2179 23545 2191 23579
rect 2133 23539 2191 23545
rect 17862 23536 17868 23588
rect 17920 23576 17926 23588
rect 21910 23576 21916 23588
rect 17920 23548 21916 23576
rect 17920 23536 17926 23548
rect 21910 23536 21916 23548
rect 21968 23536 21974 23588
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 13357 23511 13415 23517
rect 13357 23477 13369 23511
rect 13403 23508 13415 23511
rect 14090 23508 14096 23520
rect 13403 23480 14096 23508
rect 13403 23477 13415 23480
rect 13357 23471 13415 23477
rect 14090 23468 14096 23480
rect 14148 23468 14154 23520
rect 19702 23508 19708 23520
rect 19663 23480 19708 23508
rect 19702 23468 19708 23480
rect 19760 23468 19766 23520
rect 23032 23508 23060 23616
rect 23845 23613 23857 23647
rect 23891 23644 23903 23647
rect 24118 23644 24124 23656
rect 23891 23616 24124 23644
rect 23891 23613 23903 23616
rect 23845 23607 23903 23613
rect 24118 23604 24124 23616
rect 24176 23604 24182 23656
rect 24857 23647 24915 23653
rect 24857 23613 24869 23647
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 23106 23536 23112 23588
rect 23164 23576 23170 23588
rect 24872 23576 24900 23607
rect 25406 23604 25412 23656
rect 25464 23644 25470 23656
rect 27798 23644 27804 23656
rect 25464 23616 27804 23644
rect 25464 23604 25470 23616
rect 27798 23604 27804 23616
rect 27856 23644 27862 23656
rect 30101 23647 30159 23653
rect 30101 23644 30113 23647
rect 27856 23616 30113 23644
rect 27856 23604 27862 23616
rect 30101 23613 30113 23616
rect 30147 23613 30159 23647
rect 30101 23607 30159 23613
rect 27982 23576 27988 23588
rect 23164 23548 24900 23576
rect 27943 23548 27988 23576
rect 23164 23536 23170 23548
rect 27982 23536 27988 23548
rect 28040 23536 28046 23588
rect 28445 23579 28503 23585
rect 28445 23545 28457 23579
rect 28491 23576 28503 23579
rect 28994 23576 29000 23588
rect 28491 23548 29000 23576
rect 28491 23545 28503 23548
rect 28445 23539 28503 23545
rect 28994 23536 29000 23548
rect 29052 23536 29058 23588
rect 23566 23508 23572 23520
rect 23032 23480 23572 23508
rect 23566 23468 23572 23480
rect 23624 23468 23630 23520
rect 23753 23511 23811 23517
rect 23753 23477 23765 23511
rect 23799 23508 23811 23511
rect 24670 23508 24676 23520
rect 23799 23480 24676 23508
rect 23799 23477 23811 23480
rect 23753 23471 23811 23477
rect 24670 23468 24676 23480
rect 24728 23508 24734 23520
rect 24765 23511 24823 23517
rect 24765 23508 24777 23511
rect 24728 23480 24777 23508
rect 24728 23468 24734 23480
rect 24765 23477 24777 23480
rect 24811 23508 24823 23511
rect 24854 23508 24860 23520
rect 24811 23480 24860 23508
rect 24811 23477 24823 23480
rect 24765 23471 24823 23477
rect 24854 23468 24860 23480
rect 24912 23468 24918 23520
rect 28718 23468 28724 23520
rect 28776 23508 28782 23520
rect 29273 23511 29331 23517
rect 29273 23508 29285 23511
rect 28776 23480 29285 23508
rect 28776 23468 28782 23480
rect 29273 23477 29285 23480
rect 29319 23477 29331 23511
rect 29273 23471 29331 23477
rect 1104 23418 30820 23440
rect 1104 23366 5915 23418
rect 5967 23366 5979 23418
rect 6031 23366 6043 23418
rect 6095 23366 6107 23418
rect 6159 23366 6171 23418
rect 6223 23366 15846 23418
rect 15898 23366 15910 23418
rect 15962 23366 15974 23418
rect 16026 23366 16038 23418
rect 16090 23366 16102 23418
rect 16154 23366 25776 23418
rect 25828 23366 25840 23418
rect 25892 23366 25904 23418
rect 25956 23366 25968 23418
rect 26020 23366 26032 23418
rect 26084 23366 30820 23418
rect 1104 23344 30820 23366
rect 12986 23264 12992 23316
rect 13044 23304 13050 23316
rect 22646 23304 22652 23316
rect 13044 23276 22652 23304
rect 13044 23264 13050 23276
rect 22646 23264 22652 23276
rect 22704 23264 22710 23316
rect 23290 23304 23296 23316
rect 23251 23276 23296 23304
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 24397 23307 24455 23313
rect 24397 23273 24409 23307
rect 24443 23304 24455 23307
rect 24762 23304 24768 23316
rect 24443 23276 24768 23304
rect 24443 23273 24455 23276
rect 24397 23267 24455 23273
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 24854 23264 24860 23316
rect 24912 23304 24918 23316
rect 25314 23304 25320 23316
rect 24912 23276 25320 23304
rect 24912 23264 24918 23276
rect 25314 23264 25320 23276
rect 25372 23264 25378 23316
rect 28905 23307 28963 23313
rect 28905 23304 28917 23307
rect 26528 23276 28917 23304
rect 2133 23239 2191 23245
rect 2133 23205 2145 23239
rect 2179 23205 2191 23239
rect 15470 23236 15476 23248
rect 15431 23208 15476 23236
rect 2133 23199 2191 23205
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23100 1455 23103
rect 2148 23100 2176 23199
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 26421 23239 26479 23245
rect 26421 23236 26433 23239
rect 20824 23208 26433 23236
rect 14090 23168 14096 23180
rect 14051 23140 14096 23168
rect 14090 23128 14096 23140
rect 14148 23128 14154 23180
rect 19702 23128 19708 23180
rect 19760 23168 19766 23180
rect 19797 23171 19855 23177
rect 19797 23168 19809 23171
rect 19760 23140 19809 23168
rect 19760 23128 19766 23140
rect 19797 23137 19809 23140
rect 19843 23137 19855 23171
rect 19797 23131 19855 23137
rect 2314 23100 2320 23112
rect 1443 23072 2176 23100
rect 2275 23072 2320 23100
rect 1443 23069 1455 23072
rect 1397 23063 1455 23069
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 14349 23103 14407 23109
rect 14349 23100 14361 23103
rect 14240 23072 14361 23100
rect 14240 23060 14246 23072
rect 14349 23069 14361 23072
rect 14395 23069 14407 23103
rect 14349 23063 14407 23069
rect 17126 23060 17132 23112
rect 17184 23100 17190 23112
rect 20824 23100 20852 23208
rect 26421 23205 26433 23208
rect 26467 23205 26479 23239
rect 26421 23199 26479 23205
rect 21174 23128 21180 23180
rect 21232 23168 21238 23180
rect 21913 23171 21971 23177
rect 21913 23168 21925 23171
rect 21232 23140 21925 23168
rect 21232 23128 21238 23140
rect 21913 23137 21925 23140
rect 21959 23137 21971 23171
rect 21913 23131 21971 23137
rect 17184 23072 20852 23100
rect 17184 23060 17190 23072
rect 21542 23060 21548 23112
rect 21600 23100 21606 23112
rect 21637 23103 21695 23109
rect 21637 23100 21649 23103
rect 21600 23072 21649 23100
rect 21600 23060 21606 23072
rect 21637 23069 21649 23072
rect 21683 23069 21695 23103
rect 21928 23100 21956 23131
rect 22830 23128 22836 23180
rect 22888 23168 22894 23180
rect 24857 23171 24915 23177
rect 24857 23168 24869 23171
rect 22888 23140 24869 23168
rect 22888 23128 22894 23140
rect 24857 23137 24869 23140
rect 24903 23137 24915 23171
rect 26528 23168 26556 23276
rect 28905 23273 28917 23276
rect 28951 23273 28963 23307
rect 28905 23267 28963 23273
rect 29362 23264 29368 23316
rect 29420 23304 29426 23316
rect 29917 23307 29975 23313
rect 29917 23304 29929 23307
rect 29420 23276 29929 23304
rect 29420 23264 29426 23276
rect 29917 23273 29929 23276
rect 29963 23273 29975 23307
rect 29917 23267 29975 23273
rect 28077 23239 28135 23245
rect 28077 23205 28089 23239
rect 28123 23205 28135 23239
rect 28077 23199 28135 23205
rect 24857 23131 24915 23137
rect 26068 23140 26556 23168
rect 22370 23100 22376 23112
rect 21928 23072 22376 23100
rect 21637 23063 21695 23069
rect 20064 23035 20122 23041
rect 20064 23001 20076 23035
rect 20110 23032 20122 23035
rect 20714 23032 20720 23044
rect 20110 23004 20720 23032
rect 20110 23001 20122 23004
rect 20064 22995 20122 23001
rect 20714 22992 20720 23004
rect 20772 22992 20778 23044
rect 21652 23032 21680 23063
rect 22370 23060 22376 23072
rect 22428 23060 22434 23112
rect 22922 23100 22928 23112
rect 22883 23072 22928 23100
rect 22922 23060 22928 23072
rect 22980 23060 22986 23112
rect 23109 23103 23167 23109
rect 23109 23069 23121 23103
rect 23155 23069 23167 23103
rect 23109 23063 23167 23069
rect 23124 23032 23152 23063
rect 23842 23060 23848 23112
rect 23900 23100 23906 23112
rect 24578 23100 24584 23112
rect 23900 23072 24584 23100
rect 23900 23060 23906 23072
rect 24578 23060 24584 23072
rect 24636 23060 24642 23112
rect 24670 23060 24676 23112
rect 24728 23100 24734 23112
rect 24765 23103 24823 23109
rect 24765 23100 24777 23103
rect 24728 23072 24777 23100
rect 24728 23060 24734 23072
rect 24765 23069 24777 23072
rect 24811 23069 24823 23103
rect 24765 23063 24823 23069
rect 25406 23060 25412 23112
rect 25464 23100 25470 23112
rect 26068 23100 26096 23140
rect 27614 23128 27620 23180
rect 27672 23128 27678 23180
rect 28092 23168 28120 23199
rect 29362 23168 29368 23180
rect 28092 23140 29368 23168
rect 29362 23128 29368 23140
rect 29420 23168 29426 23180
rect 29420 23140 29776 23168
rect 29420 23128 29426 23140
rect 25464 23072 26096 23100
rect 25464 23060 25470 23072
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26697 23103 26755 23109
rect 26697 23100 26709 23103
rect 26200 23072 26709 23100
rect 26200 23060 26206 23072
rect 26697 23069 26709 23072
rect 26743 23069 26755 23103
rect 27632 23100 27660 23128
rect 28261 23103 28319 23109
rect 28261 23100 28273 23103
rect 27632 23072 28273 23100
rect 26697 23063 26755 23069
rect 28261 23069 28273 23072
rect 28307 23069 28319 23103
rect 28261 23063 28319 23069
rect 28721 23103 28779 23109
rect 28721 23069 28733 23103
rect 28767 23100 28779 23103
rect 28902 23100 28908 23112
rect 28767 23072 28908 23100
rect 28767 23069 28779 23072
rect 28721 23063 28779 23069
rect 28902 23060 28908 23072
rect 28960 23060 28966 23112
rect 29748 23109 29776 23140
rect 29733 23103 29791 23109
rect 29733 23069 29745 23103
rect 29779 23069 29791 23103
rect 29733 23063 29791 23069
rect 21192 23004 23152 23032
rect 1578 22964 1584 22976
rect 1539 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 21192 22973 21220 23004
rect 24946 22992 24952 23044
rect 25004 23032 25010 23044
rect 25130 23032 25136 23044
rect 25004 23004 25136 23032
rect 25004 22992 25010 23004
rect 25130 22992 25136 23004
rect 25188 22992 25194 23044
rect 26973 23035 27031 23041
rect 26973 23001 26985 23035
rect 27019 23032 27031 23035
rect 27614 23032 27620 23044
rect 27019 23004 27620 23032
rect 27019 23001 27031 23004
rect 26973 22995 27031 23001
rect 27614 22992 27620 23004
rect 27672 22992 27678 23044
rect 28994 22992 29000 23044
rect 29052 23032 29058 23044
rect 29549 23035 29607 23041
rect 29549 23032 29561 23035
rect 29052 23004 29561 23032
rect 29052 22992 29058 23004
rect 29549 23001 29561 23004
rect 29595 23001 29607 23035
rect 29549 22995 29607 23001
rect 21177 22967 21235 22973
rect 21177 22933 21189 22967
rect 21223 22933 21235 22967
rect 21177 22927 21235 22933
rect 23014 22924 23020 22976
rect 23072 22964 23078 22976
rect 23566 22964 23572 22976
rect 23072 22936 23572 22964
rect 23072 22924 23078 22936
rect 23566 22924 23572 22936
rect 23624 22924 23630 22976
rect 24762 22924 24768 22976
rect 24820 22964 24826 22976
rect 25314 22964 25320 22976
rect 24820 22936 25320 22964
rect 24820 22924 24826 22936
rect 25314 22924 25320 22936
rect 25372 22924 25378 22976
rect 26694 22924 26700 22976
rect 26752 22964 26758 22976
rect 26881 22967 26939 22973
rect 26881 22964 26893 22967
rect 26752 22936 26893 22964
rect 26752 22924 26758 22936
rect 26881 22933 26893 22936
rect 26927 22933 26939 22967
rect 26881 22927 26939 22933
rect 29086 22924 29092 22976
rect 29144 22964 29150 22976
rect 29270 22964 29276 22976
rect 29144 22936 29276 22964
rect 29144 22924 29150 22936
rect 29270 22924 29276 22936
rect 29328 22924 29334 22976
rect 1104 22874 30820 22896
rect 1104 22822 10880 22874
rect 10932 22822 10944 22874
rect 10996 22822 11008 22874
rect 11060 22822 11072 22874
rect 11124 22822 11136 22874
rect 11188 22822 20811 22874
rect 20863 22822 20875 22874
rect 20927 22822 20939 22874
rect 20991 22822 21003 22874
rect 21055 22822 21067 22874
rect 21119 22822 30820 22874
rect 1104 22800 30820 22822
rect 2314 22720 2320 22772
rect 2372 22760 2378 22772
rect 17126 22760 17132 22772
rect 2372 22732 17132 22760
rect 2372 22720 2378 22732
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17957 22763 18015 22769
rect 17957 22729 17969 22763
rect 18003 22760 18015 22763
rect 18138 22760 18144 22772
rect 18003 22732 18144 22760
rect 18003 22729 18015 22732
rect 17957 22723 18015 22729
rect 18138 22720 18144 22732
rect 18196 22720 18202 22772
rect 20993 22763 21051 22769
rect 20993 22729 21005 22763
rect 21039 22729 21051 22763
rect 20993 22723 21051 22729
rect 21821 22763 21879 22769
rect 21821 22729 21833 22763
rect 21867 22760 21879 22763
rect 22186 22760 22192 22772
rect 21867 22732 22192 22760
rect 21867 22729 21879 22732
rect 21821 22723 21879 22729
rect 21008 22692 21036 22723
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 22646 22720 22652 22772
rect 22704 22760 22710 22772
rect 28243 22763 28301 22769
rect 28243 22760 28255 22763
rect 22704 22732 28255 22760
rect 22704 22720 22710 22732
rect 28243 22729 28255 22732
rect 28289 22729 28301 22763
rect 29822 22760 29828 22772
rect 29783 22732 29828 22760
rect 28243 22723 28301 22729
rect 29822 22720 29828 22732
rect 29880 22720 29886 22772
rect 22094 22692 22100 22704
rect 21008 22664 22100 22692
rect 22094 22652 22100 22664
rect 22152 22652 22158 22704
rect 22370 22692 22376 22704
rect 22204 22664 22376 22692
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22624 1455 22627
rect 2317 22627 2375 22633
rect 1443 22596 2176 22624
rect 1443 22593 1455 22596
rect 1397 22587 1455 22593
rect 2148 22497 2176 22596
rect 2317 22593 2329 22627
rect 2363 22624 2375 22627
rect 17862 22624 17868 22636
rect 2363 22596 6914 22624
rect 17823 22596 17868 22624
rect 2363 22593 2375 22596
rect 2317 22587 2375 22593
rect 2133 22491 2191 22497
rect 2133 22457 2145 22491
rect 2179 22457 2191 22491
rect 6886 22488 6914 22596
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 20993 22627 21051 22633
rect 20993 22593 21005 22627
rect 21039 22624 21051 22627
rect 21174 22624 21180 22636
rect 21039 22596 21180 22624
rect 21039 22593 21051 22596
rect 20993 22587 21051 22593
rect 21174 22584 21180 22596
rect 21232 22584 21238 22636
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22624 21327 22627
rect 21634 22624 21640 22636
rect 21315 22596 21640 22624
rect 21315 22593 21327 22596
rect 21269 22587 21327 22593
rect 21634 22584 21640 22596
rect 21692 22624 21698 22636
rect 22204 22633 22232 22664
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 26694 22652 26700 22704
rect 26752 22692 26758 22704
rect 27341 22695 27399 22701
rect 27341 22692 27353 22695
rect 26752 22664 27353 22692
rect 26752 22652 26758 22664
rect 27341 22661 27353 22664
rect 27387 22661 27399 22695
rect 27341 22655 27399 22661
rect 27525 22695 27583 22701
rect 27525 22661 27537 22695
rect 27571 22661 27583 22695
rect 27525 22655 27583 22661
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21692 22596 22017 22624
rect 21692 22584 21698 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 22281 22627 22339 22633
rect 22281 22593 22293 22627
rect 22327 22624 22339 22627
rect 22922 22624 22928 22636
rect 22327 22596 22928 22624
rect 22327 22593 22339 22596
rect 22281 22587 22339 22593
rect 12406 22528 21312 22556
rect 12406 22488 12434 22528
rect 6886 22460 12434 22488
rect 21085 22491 21143 22497
rect 2133 22451 2191 22457
rect 21085 22457 21097 22491
rect 21131 22457 21143 22491
rect 21284 22488 21312 22528
rect 21358 22516 21364 22568
rect 21416 22556 21422 22568
rect 22296 22556 22324 22587
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 23198 22584 23204 22636
rect 23256 22624 23262 22636
rect 23385 22627 23443 22633
rect 23385 22624 23397 22627
rect 23256 22596 23397 22624
rect 23256 22584 23262 22596
rect 23385 22593 23397 22596
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 23474 22584 23480 22636
rect 23532 22624 23538 22636
rect 23569 22627 23627 22633
rect 23569 22624 23581 22627
rect 23532 22596 23581 22624
rect 23532 22584 23538 22596
rect 23569 22593 23581 22596
rect 23615 22624 23627 22627
rect 23934 22624 23940 22636
rect 23615 22596 23940 22624
rect 23615 22593 23627 22596
rect 23569 22587 23627 22593
rect 23934 22584 23940 22596
rect 23992 22584 23998 22636
rect 24302 22584 24308 22636
rect 24360 22624 24366 22636
rect 25406 22624 25412 22636
rect 24360 22596 25268 22624
rect 25367 22596 25412 22624
rect 24360 22584 24366 22596
rect 21416 22528 22324 22556
rect 23661 22559 23719 22565
rect 21416 22516 21422 22528
rect 23661 22525 23673 22559
rect 23707 22556 23719 22559
rect 25130 22556 25136 22568
rect 23707 22528 25136 22556
rect 23707 22525 23719 22528
rect 23661 22519 23719 22525
rect 25130 22516 25136 22528
rect 25188 22516 25194 22568
rect 25240 22556 25268 22596
rect 25406 22584 25412 22596
rect 25464 22584 25470 22636
rect 25685 22627 25743 22633
rect 25685 22593 25697 22627
rect 25731 22624 25743 22627
rect 26234 22624 26240 22636
rect 25731 22596 26240 22624
rect 25731 22593 25743 22596
rect 25685 22587 25743 22593
rect 26234 22584 26240 22596
rect 26292 22584 26298 22636
rect 27540 22556 27568 22655
rect 27614 22652 27620 22704
rect 27672 22692 27678 22704
rect 28721 22695 28779 22701
rect 27672 22664 27717 22692
rect 27672 22652 27678 22664
rect 28721 22661 28733 22695
rect 28767 22692 28779 22695
rect 28767 22664 29316 22692
rect 28767 22661 28779 22664
rect 28721 22655 28779 22661
rect 28537 22627 28595 22633
rect 28537 22593 28549 22627
rect 28583 22624 28595 22627
rect 28994 22624 29000 22636
rect 28583 22596 29000 22624
rect 28583 22593 28595 22596
rect 28537 22587 28595 22593
rect 28994 22584 29000 22596
rect 29052 22584 29058 22636
rect 25240 22528 27568 22556
rect 28626 22516 28632 22568
rect 28684 22556 28690 22568
rect 28813 22559 28871 22565
rect 28813 22556 28825 22559
rect 28684 22528 28825 22556
rect 28684 22516 28690 22528
rect 28813 22525 28825 22528
rect 28859 22525 28871 22559
rect 29288 22556 29316 22664
rect 29362 22652 29368 22704
rect 29420 22692 29426 22704
rect 29641 22695 29699 22701
rect 29641 22692 29653 22695
rect 29420 22664 29653 22692
rect 29420 22652 29426 22664
rect 29641 22661 29653 22664
rect 29687 22661 29699 22695
rect 29641 22655 29699 22661
rect 29454 22624 29460 22636
rect 29415 22596 29460 22624
rect 29454 22584 29460 22596
rect 29512 22584 29518 22636
rect 31478 22556 31484 22568
rect 29288 22528 31484 22556
rect 28813 22519 28871 22525
rect 31478 22516 31484 22528
rect 31536 22516 31542 22568
rect 21284 22460 21404 22488
rect 21085 22451 21143 22457
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 21100 22420 21128 22451
rect 21266 22420 21272 22432
rect 21100 22392 21272 22420
rect 21266 22380 21272 22392
rect 21324 22380 21330 22432
rect 21376 22420 21404 22460
rect 22370 22448 22376 22500
rect 22428 22488 22434 22500
rect 23201 22491 23259 22497
rect 23201 22488 23213 22491
rect 22428 22460 23213 22488
rect 22428 22448 22434 22460
rect 23201 22457 23213 22460
rect 23247 22457 23259 22491
rect 27065 22491 27123 22497
rect 27065 22488 27077 22491
rect 23201 22451 23259 22457
rect 23308 22460 27077 22488
rect 23308 22420 23336 22460
rect 27065 22457 27077 22460
rect 27111 22457 27123 22491
rect 27065 22451 27123 22457
rect 21376 22392 23336 22420
rect 25225 22423 25283 22429
rect 25225 22389 25237 22423
rect 25271 22420 25283 22423
rect 25314 22420 25320 22432
rect 25271 22392 25320 22420
rect 25271 22389 25283 22392
rect 25225 22383 25283 22389
rect 25314 22380 25320 22392
rect 25372 22380 25378 22432
rect 25590 22420 25596 22432
rect 25551 22392 25596 22420
rect 25590 22380 25596 22392
rect 25648 22380 25654 22432
rect 26694 22380 26700 22432
rect 26752 22420 26758 22432
rect 28718 22420 28724 22432
rect 26752 22392 28724 22420
rect 26752 22380 26758 22392
rect 28718 22380 28724 22392
rect 28776 22380 28782 22432
rect 1104 22330 30820 22352
rect 1104 22278 5915 22330
rect 5967 22278 5979 22330
rect 6031 22278 6043 22330
rect 6095 22278 6107 22330
rect 6159 22278 6171 22330
rect 6223 22278 15846 22330
rect 15898 22278 15910 22330
rect 15962 22278 15974 22330
rect 16026 22278 16038 22330
rect 16090 22278 16102 22330
rect 16154 22278 25776 22330
rect 25828 22278 25840 22330
rect 25892 22278 25904 22330
rect 25956 22278 25968 22330
rect 26020 22278 26032 22330
rect 26084 22278 30820 22330
rect 1104 22256 30820 22278
rect 22094 22176 22100 22228
rect 22152 22216 22158 22228
rect 22554 22216 22560 22228
rect 22152 22188 22560 22216
rect 22152 22176 22158 22188
rect 22554 22176 22560 22188
rect 22612 22176 22618 22228
rect 26234 22176 26240 22228
rect 26292 22216 26298 22228
rect 26421 22219 26479 22225
rect 26421 22216 26433 22219
rect 26292 22188 26433 22216
rect 26292 22176 26298 22188
rect 26421 22185 26433 22188
rect 26467 22185 26479 22219
rect 26421 22179 26479 22185
rect 26786 22176 26792 22228
rect 26844 22216 26850 22228
rect 26844 22188 27476 22216
rect 26844 22176 26850 22188
rect 27448 22160 27476 22188
rect 27522 22176 27528 22228
rect 27580 22176 27586 22228
rect 28442 22176 28448 22228
rect 28500 22216 28506 22228
rect 28902 22216 28908 22228
rect 28500 22188 28908 22216
rect 28500 22176 28506 22188
rect 28902 22176 28908 22188
rect 28960 22176 28966 22228
rect 30009 22219 30067 22225
rect 30009 22216 30021 22219
rect 29012 22188 30021 22216
rect 27430 22108 27436 22160
rect 27488 22108 27494 22160
rect 22066 22052 25176 22080
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 1903 21984 6914 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 6886 21944 6914 21984
rect 18506 21972 18512 22024
rect 18564 22012 18570 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 18564 21984 19257 22012
rect 18564 21972 18570 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19245 21975 19303 21981
rect 22066 21944 22094 22052
rect 22278 21972 22284 22024
rect 22336 22012 22342 22024
rect 22465 22015 22523 22021
rect 22465 22012 22477 22015
rect 22336 21984 22477 22012
rect 22336 21972 22342 21984
rect 22465 21981 22477 21984
rect 22511 21981 22523 22015
rect 25041 22015 25099 22021
rect 25041 22012 25053 22015
rect 22465 21975 22523 21981
rect 22572 21984 25053 22012
rect 6886 21916 22094 21944
rect 22572 21888 22600 21984
rect 25041 21981 25053 21984
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 22738 21904 22744 21956
rect 22796 21944 22802 21956
rect 23106 21944 23112 21956
rect 22796 21916 23112 21944
rect 22796 21904 22802 21916
rect 23106 21904 23112 21916
rect 23164 21904 23170 21956
rect 25148 21944 25176 22052
rect 26234 22040 26240 22092
rect 26292 22080 26298 22092
rect 27157 22083 27215 22089
rect 27157 22080 27169 22083
rect 26292 22052 27169 22080
rect 26292 22040 26298 22052
rect 27157 22049 27169 22052
rect 27203 22049 27215 22083
rect 27157 22043 27215 22049
rect 27341 22083 27399 22089
rect 27341 22049 27353 22083
rect 27387 22080 27399 22083
rect 27540 22080 27568 22176
rect 27706 22080 27712 22092
rect 27387 22052 27712 22080
rect 27387 22049 27399 22052
rect 27341 22043 27399 22049
rect 27706 22040 27712 22052
rect 27764 22080 27770 22092
rect 28626 22080 28632 22092
rect 27764 22052 28632 22080
rect 27764 22040 27770 22052
rect 28626 22040 28632 22052
rect 28684 22080 28690 22092
rect 28721 22083 28779 22089
rect 28721 22080 28733 22083
rect 28684 22052 28733 22080
rect 28684 22040 28690 22052
rect 28721 22049 28733 22052
rect 28767 22049 28779 22083
rect 28721 22043 28779 22049
rect 25314 22021 25320 22024
rect 25308 21975 25320 22021
rect 25372 22012 25378 22024
rect 28151 22015 28209 22021
rect 28151 22012 28163 22015
rect 25372 21984 25408 22012
rect 25516 21984 28163 22012
rect 25314 21972 25320 21975
rect 25372 21972 25378 21984
rect 25516 21944 25544 21984
rect 28151 21981 28163 21984
rect 28197 21981 28209 22015
rect 28151 21975 28209 21981
rect 28258 21972 28264 22024
rect 28316 22012 28322 22024
rect 29012 22012 29040 22188
rect 30009 22185 30021 22188
rect 30055 22185 30067 22219
rect 30009 22179 30067 22185
rect 30282 22040 30288 22092
rect 30340 22040 30346 22092
rect 28316 21984 29040 22012
rect 28316 21972 28322 21984
rect 29362 21972 29368 22024
rect 29420 22012 29426 22024
rect 29825 22015 29883 22021
rect 29825 22012 29837 22015
rect 29420 21984 29837 22012
rect 29420 21972 29426 21984
rect 29825 21981 29837 21984
rect 29871 22012 29883 22015
rect 29914 22012 29920 22024
rect 29871 21984 29920 22012
rect 29871 21981 29883 21984
rect 29825 21975 29883 21981
rect 29914 21972 29920 21984
rect 29972 21972 29978 22024
rect 25148 21916 25544 21944
rect 25590 21904 25596 21956
rect 25648 21944 25654 21956
rect 26142 21944 26148 21956
rect 25648 21916 26148 21944
rect 25648 21904 25654 21916
rect 26142 21904 26148 21916
rect 26200 21904 26206 21956
rect 27246 21944 27252 21956
rect 27207 21916 27252 21944
rect 27246 21904 27252 21916
rect 27304 21904 27310 21956
rect 27798 21944 27804 21956
rect 27759 21916 27804 21944
rect 27798 21904 27804 21916
rect 27856 21904 27862 21956
rect 28442 21944 28448 21956
rect 28403 21916 28448 21944
rect 28442 21904 28448 21916
rect 28500 21944 28506 21956
rect 28810 21944 28816 21956
rect 28500 21916 28816 21944
rect 28500 21904 28506 21916
rect 28810 21904 28816 21916
rect 28868 21904 28874 21956
rect 29638 21944 29644 21956
rect 29599 21916 29644 21944
rect 29638 21904 29644 21916
rect 29696 21904 29702 21956
rect 30006 21904 30012 21956
rect 30064 21944 30070 21956
rect 30300 21944 30328 22040
rect 30064 21916 30328 21944
rect 30064 21904 30070 21916
rect 1394 21836 1400 21888
rect 1452 21876 1458 21888
rect 1673 21879 1731 21885
rect 1673 21876 1685 21879
rect 1452 21848 1685 21876
rect 1452 21836 1458 21848
rect 1673 21845 1685 21848
rect 1719 21845 1731 21879
rect 1673 21839 1731 21845
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 19889 21879 19947 21885
rect 19889 21876 19901 21879
rect 19300 21848 19901 21876
rect 19300 21836 19306 21848
rect 19889 21845 19901 21848
rect 19935 21845 19947 21879
rect 22554 21876 22560 21888
rect 22515 21848 22560 21876
rect 19889 21839 19947 21845
rect 22554 21836 22560 21848
rect 22612 21836 22618 21888
rect 24394 21836 24400 21888
rect 24452 21876 24458 21888
rect 26771 21879 26829 21885
rect 26771 21876 26783 21879
rect 24452 21848 26783 21876
rect 24452 21836 24458 21848
rect 26771 21845 26783 21848
rect 26817 21845 26829 21879
rect 27816 21876 27844 21904
rect 28629 21879 28687 21885
rect 28629 21876 28641 21879
rect 27816 21848 28641 21876
rect 26771 21839 26829 21845
rect 28629 21845 28641 21848
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 29178 21836 29184 21888
rect 29236 21876 29242 21888
rect 30558 21876 30564 21888
rect 29236 21848 30564 21876
rect 29236 21836 29242 21848
rect 30558 21836 30564 21848
rect 30616 21836 30622 21888
rect 1104 21786 30820 21808
rect 1104 21734 10880 21786
rect 10932 21734 10944 21786
rect 10996 21734 11008 21786
rect 11060 21734 11072 21786
rect 11124 21734 11136 21786
rect 11188 21734 20811 21786
rect 20863 21734 20875 21786
rect 20927 21734 20939 21786
rect 20991 21734 21003 21786
rect 21055 21734 21067 21786
rect 21119 21734 30820 21786
rect 1104 21712 30820 21734
rect 17862 21632 17868 21684
rect 17920 21672 17926 21684
rect 18693 21675 18751 21681
rect 18693 21672 18705 21675
rect 17920 21644 18705 21672
rect 17920 21632 17926 21644
rect 18693 21641 18705 21644
rect 18739 21641 18751 21675
rect 18693 21635 18751 21641
rect 23290 21632 23296 21684
rect 23348 21672 23354 21684
rect 24029 21675 24087 21681
rect 24029 21672 24041 21675
rect 23348 21644 24041 21672
rect 23348 21632 23354 21644
rect 24029 21641 24041 21644
rect 24075 21641 24087 21675
rect 24029 21635 24087 21641
rect 24762 21632 24768 21684
rect 24820 21632 24826 21684
rect 25225 21675 25283 21681
rect 25225 21641 25237 21675
rect 25271 21672 25283 21675
rect 25406 21672 25412 21684
rect 25271 21644 25412 21672
rect 25271 21641 25283 21644
rect 25225 21635 25283 21641
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 26050 21632 26056 21684
rect 26108 21672 26114 21684
rect 26234 21672 26240 21684
rect 26108 21644 26240 21672
rect 26108 21632 26114 21644
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 27617 21675 27675 21681
rect 27617 21641 27629 21675
rect 27663 21672 27675 21675
rect 27706 21672 27712 21684
rect 27663 21644 27712 21672
rect 27663 21641 27675 21644
rect 27617 21635 27675 21641
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 28994 21632 29000 21684
rect 29052 21672 29058 21684
rect 29089 21675 29147 21681
rect 29089 21672 29101 21675
rect 29052 21644 29101 21672
rect 29052 21632 29058 21644
rect 29089 21641 29101 21644
rect 29135 21641 29147 21675
rect 29089 21635 29147 21641
rect 30101 21675 30159 21681
rect 30101 21641 30113 21675
rect 30147 21672 30159 21675
rect 30190 21672 30196 21684
rect 30147 21644 30196 21672
rect 30147 21641 30159 21644
rect 30101 21635 30159 21641
rect 30190 21632 30196 21644
rect 30248 21632 30254 21684
rect 24578 21604 24584 21616
rect 24228 21576 24584 21604
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21496 1458 21548
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21536 2375 21539
rect 16666 21536 16672 21548
rect 2363 21508 6914 21536
rect 16627 21508 16672 21536
rect 2363 21505 2375 21508
rect 2317 21499 2375 21505
rect 1578 21400 1584 21412
rect 1539 21372 1584 21400
rect 1578 21360 1584 21372
rect 1636 21360 1642 21412
rect 6886 21400 6914 21508
rect 16666 21496 16672 21508
rect 16724 21496 16730 21548
rect 17865 21539 17923 21545
rect 17865 21505 17877 21539
rect 17911 21536 17923 21539
rect 18414 21536 18420 21548
rect 17911 21508 18420 21536
rect 17911 21505 17923 21508
rect 17865 21499 17923 21505
rect 18414 21496 18420 21508
rect 18472 21496 18478 21548
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21536 18567 21539
rect 18598 21536 18604 21548
rect 18555 21508 18604 21536
rect 18555 21505 18567 21508
rect 18509 21499 18567 21505
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21505 18843 21539
rect 19242 21536 19248 21548
rect 19203 21508 19248 21536
rect 18785 21499 18843 21505
rect 18138 21428 18144 21480
rect 18196 21468 18202 21480
rect 18800 21468 18828 21499
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21536 19487 21539
rect 19610 21536 19616 21548
rect 19475 21508 19616 21536
rect 19475 21505 19487 21508
rect 19429 21499 19487 21505
rect 19610 21496 19616 21508
rect 19668 21536 19674 21548
rect 22370 21536 22376 21548
rect 19668 21508 22376 21536
rect 19668 21496 19674 21508
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 24228 21545 24256 21576
rect 24578 21564 24584 21576
rect 24636 21564 24642 21616
rect 24213 21539 24271 21545
rect 24213 21505 24225 21539
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 24489 21539 24547 21545
rect 24489 21505 24501 21539
rect 24535 21536 24547 21539
rect 24673 21539 24731 21545
rect 24535 21508 24624 21536
rect 24535 21505 24547 21508
rect 24489 21499 24547 21505
rect 18196 21440 18828 21468
rect 24596 21468 24624 21508
rect 24673 21505 24685 21539
rect 24719 21536 24731 21539
rect 24780 21536 24808 21632
rect 25590 21564 25596 21616
rect 25648 21604 25654 21616
rect 25958 21604 25964 21616
rect 25648 21576 25964 21604
rect 25648 21564 25654 21576
rect 25958 21564 25964 21576
rect 26016 21564 26022 21616
rect 27338 21564 27344 21616
rect 27396 21604 27402 21616
rect 27525 21607 27583 21613
rect 27525 21604 27537 21607
rect 27396 21576 27537 21604
rect 27396 21564 27402 21576
rect 27525 21573 27537 21576
rect 27571 21604 27583 21607
rect 27571 21576 28212 21604
rect 27571 21573 27583 21576
rect 27525 21567 27583 21573
rect 28184 21548 28212 21576
rect 28626 21564 28632 21616
rect 28684 21604 28690 21616
rect 29733 21607 29791 21613
rect 29733 21604 29745 21607
rect 28684 21576 29745 21604
rect 28684 21564 28690 21576
rect 29733 21573 29745 21576
rect 29779 21573 29791 21607
rect 29914 21604 29920 21616
rect 29875 21576 29920 21604
rect 29733 21567 29791 21573
rect 29914 21564 29920 21576
rect 29972 21564 29978 21616
rect 24719 21508 24808 21536
rect 24719 21505 24731 21508
rect 24673 21499 24731 21505
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 25406 21536 25412 21548
rect 25188 21508 25412 21536
rect 25188 21496 25194 21508
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21536 25927 21539
rect 26786 21536 26792 21548
rect 25915 21508 26792 21536
rect 25915 21505 25927 21508
rect 25869 21499 25927 21505
rect 24854 21468 24860 21480
rect 24596 21440 24860 21468
rect 18196 21428 18202 21440
rect 24854 21428 24860 21440
rect 24912 21468 24918 21480
rect 25700 21468 25728 21499
rect 26786 21496 26792 21508
rect 26844 21496 26850 21548
rect 28166 21536 28172 21548
rect 28079 21508 28172 21536
rect 28166 21496 28172 21508
rect 28224 21496 28230 21548
rect 29270 21536 29276 21548
rect 29231 21508 29276 21536
rect 29270 21496 29276 21508
rect 29328 21496 29334 21548
rect 24912 21440 25728 21468
rect 28445 21471 28503 21477
rect 24912 21428 24918 21440
rect 28445 21437 28457 21471
rect 28491 21468 28503 21471
rect 29362 21468 29368 21480
rect 28491 21440 29368 21468
rect 28491 21437 28503 21440
rect 28445 21431 28503 21437
rect 29362 21428 29368 21440
rect 29420 21468 29426 21480
rect 30190 21468 30196 21480
rect 29420 21440 30196 21468
rect 29420 21428 29426 21440
rect 30190 21428 30196 21440
rect 30248 21428 30254 21480
rect 24394 21400 24400 21412
rect 6886 21372 24400 21400
rect 24394 21360 24400 21372
rect 24452 21360 24458 21412
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 2133 21335 2191 21341
rect 2133 21332 2145 21335
rect 1452 21304 2145 21332
rect 1452 21292 1458 21304
rect 2133 21301 2145 21304
rect 2179 21301 2191 21335
rect 2133 21295 2191 21301
rect 16666 21292 16672 21344
rect 16724 21332 16730 21344
rect 16853 21335 16911 21341
rect 16853 21332 16865 21335
rect 16724 21304 16865 21332
rect 16724 21292 16730 21304
rect 16853 21301 16865 21304
rect 16899 21301 16911 21335
rect 18046 21332 18052 21344
rect 18007 21304 18052 21332
rect 16853 21295 16911 21301
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 18506 21332 18512 21344
rect 18467 21304 18512 21332
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 19245 21335 19303 21341
rect 19245 21301 19257 21335
rect 19291 21332 19303 21335
rect 19334 21332 19340 21344
rect 19291 21304 19340 21332
rect 19291 21301 19303 21304
rect 19245 21295 19303 21301
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 1104 21242 30820 21264
rect 1104 21190 5915 21242
rect 5967 21190 5979 21242
rect 6031 21190 6043 21242
rect 6095 21190 6107 21242
rect 6159 21190 6171 21242
rect 6223 21190 15846 21242
rect 15898 21190 15910 21242
rect 15962 21190 15974 21242
rect 16026 21190 16038 21242
rect 16090 21190 16102 21242
rect 16154 21190 25776 21242
rect 25828 21190 25840 21242
rect 25892 21190 25904 21242
rect 25956 21190 25968 21242
rect 26020 21190 26032 21242
rect 26084 21190 30820 21242
rect 1104 21168 30820 21190
rect 12710 21088 12716 21140
rect 12768 21128 12774 21140
rect 16945 21131 17003 21137
rect 16945 21128 16957 21131
rect 12768 21100 16957 21128
rect 12768 21088 12774 21100
rect 16945 21097 16957 21100
rect 16991 21097 17003 21131
rect 16945 21091 17003 21097
rect 23566 21088 23572 21140
rect 23624 21128 23630 21140
rect 24397 21131 24455 21137
rect 24397 21128 24409 21131
rect 23624 21100 24409 21128
rect 23624 21088 23630 21100
rect 24397 21097 24409 21100
rect 24443 21097 24455 21131
rect 27430 21128 27436 21140
rect 27391 21100 27436 21128
rect 24397 21091 24455 21097
rect 27430 21088 27436 21100
rect 27488 21088 27494 21140
rect 28077 21131 28135 21137
rect 28077 21097 28089 21131
rect 28123 21128 28135 21131
rect 29178 21128 29184 21140
rect 28123 21100 29184 21128
rect 28123 21097 28135 21100
rect 28077 21091 28135 21097
rect 29178 21088 29184 21100
rect 29236 21088 29242 21140
rect 30098 21128 30104 21140
rect 30059 21100 30104 21128
rect 30098 21088 30104 21100
rect 30156 21088 30162 21140
rect 17865 20995 17923 21001
rect 17865 20992 17877 20995
rect 16776 20964 17877 20992
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 16776 20933 16804 20964
rect 17865 20961 17877 20964
rect 17911 20961 17923 20995
rect 17865 20955 17923 20961
rect 18046 20952 18052 21004
rect 18104 20992 18110 21004
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 18104 20964 19257 20992
rect 18104 20952 18110 20964
rect 19245 20961 19257 20964
rect 19291 20961 19303 20995
rect 28997 20995 29055 21001
rect 28997 20992 29009 20995
rect 19245 20955 19303 20961
rect 25608 20964 29009 20992
rect 25608 20936 25636 20964
rect 28997 20961 29009 20964
rect 29043 20961 29055 20995
rect 28997 20955 29055 20961
rect 16761 20927 16819 20933
rect 16761 20893 16773 20927
rect 16807 20893 16819 20927
rect 16761 20887 16819 20893
rect 17589 20927 17647 20933
rect 17589 20893 17601 20927
rect 17635 20893 17647 20927
rect 17589 20887 17647 20893
rect 17681 20927 17739 20933
rect 17681 20893 17693 20927
rect 17727 20924 17739 20927
rect 17770 20924 17776 20936
rect 17727 20896 17776 20924
rect 17727 20893 17739 20896
rect 17681 20887 17739 20893
rect 17604 20856 17632 20887
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19501 20927 19559 20933
rect 19501 20924 19513 20927
rect 19392 20896 19513 20924
rect 19392 20884 19398 20896
rect 19501 20893 19513 20896
rect 19547 20893 19559 20927
rect 24578 20924 24584 20936
rect 24539 20896 24584 20924
rect 19501 20887 19559 20893
rect 24578 20884 24584 20896
rect 24636 20884 24642 20936
rect 24854 20924 24860 20936
rect 24815 20896 24860 20924
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 25041 20927 25099 20933
rect 25041 20893 25053 20927
rect 25087 20924 25099 20927
rect 25590 20924 25596 20936
rect 25087 20896 25596 20924
rect 25087 20893 25099 20896
rect 25041 20887 25099 20893
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 27614 20924 27620 20936
rect 27575 20896 27620 20924
rect 27614 20884 27620 20896
rect 27672 20884 27678 20936
rect 28258 20924 28264 20936
rect 28219 20896 28264 20924
rect 28258 20884 28264 20896
rect 28316 20884 28322 20936
rect 29914 20924 29920 20936
rect 29875 20896 29920 20924
rect 29914 20884 29920 20896
rect 29972 20884 29978 20936
rect 18046 20856 18052 20868
rect 17604 20828 18052 20856
rect 18046 20816 18052 20828
rect 18104 20816 18110 20868
rect 26418 20816 26424 20868
rect 26476 20856 26482 20868
rect 26878 20856 26884 20868
rect 26476 20828 26884 20856
rect 26476 20816 26482 20828
rect 26878 20816 26884 20828
rect 26936 20816 26942 20868
rect 28810 20856 28816 20868
rect 28771 20828 28816 20856
rect 28810 20816 28816 20828
rect 28868 20816 28874 20868
rect 29178 20816 29184 20868
rect 29236 20856 29242 20868
rect 29733 20859 29791 20865
rect 29733 20856 29745 20859
rect 29236 20828 29745 20856
rect 29236 20816 29242 20828
rect 29733 20825 29745 20828
rect 29779 20825 29791 20859
rect 29733 20819 29791 20825
rect 1578 20788 1584 20800
rect 1539 20760 1584 20788
rect 1578 20748 1584 20760
rect 1636 20748 1642 20800
rect 20622 20788 20628 20800
rect 20583 20760 20628 20788
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 1104 20698 30820 20720
rect 1104 20646 10880 20698
rect 10932 20646 10944 20698
rect 10996 20646 11008 20698
rect 11060 20646 11072 20698
rect 11124 20646 11136 20698
rect 11188 20646 20811 20698
rect 20863 20646 20875 20698
rect 20927 20646 20939 20698
rect 20991 20646 21003 20698
rect 21055 20646 21067 20698
rect 21119 20646 30820 20698
rect 1104 20624 30820 20646
rect 2314 20544 2320 20596
rect 2372 20584 2378 20596
rect 29439 20587 29497 20593
rect 29439 20584 29451 20587
rect 2372 20556 29451 20584
rect 2372 20544 2378 20556
rect 29439 20553 29451 20556
rect 29485 20553 29497 20587
rect 29439 20547 29497 20553
rect 29917 20587 29975 20593
rect 29917 20553 29929 20587
rect 29963 20584 29975 20587
rect 31570 20584 31576 20596
rect 29963 20556 31576 20584
rect 29963 20553 29975 20556
rect 29917 20547 29975 20553
rect 31570 20544 31576 20556
rect 31628 20544 31634 20596
rect 20073 20519 20131 20525
rect 20073 20485 20085 20519
rect 20119 20516 20131 20519
rect 20622 20516 20628 20528
rect 20119 20488 20628 20516
rect 20119 20485 20131 20488
rect 20073 20479 20131 20485
rect 20622 20476 20628 20488
rect 20680 20476 20686 20528
rect 28166 20476 28172 20528
rect 28224 20516 28230 20528
rect 28261 20519 28319 20525
rect 28261 20516 28273 20519
rect 28224 20488 28273 20516
rect 28224 20476 28230 20488
rect 28261 20485 28273 20488
rect 28307 20485 28319 20519
rect 28261 20479 28319 20485
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20448 1455 20451
rect 2130 20448 2136 20460
rect 1443 20420 2136 20448
rect 1443 20417 1455 20420
rect 1397 20411 1455 20417
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 16482 20448 16488 20460
rect 16163 20420 16488 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 16925 20451 16983 20457
rect 16925 20448 16937 20451
rect 16776 20420 16937 20448
rect 16776 20380 16804 20420
rect 16925 20417 16937 20420
rect 16971 20417 16983 20451
rect 16925 20411 16983 20417
rect 18046 20408 18052 20460
rect 18104 20448 18110 20460
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 18104 20420 18613 20448
rect 18104 20408 18110 20420
rect 18601 20417 18613 20420
rect 18647 20448 18659 20451
rect 19242 20448 19248 20460
rect 18647 20420 19248 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 19242 20408 19248 20420
rect 19300 20408 19306 20460
rect 29178 20408 29184 20460
rect 29236 20448 29242 20460
rect 29733 20451 29791 20457
rect 29733 20448 29745 20451
rect 29236 20420 29745 20448
rect 29236 20408 29242 20420
rect 29733 20417 29745 20420
rect 29779 20417 29791 20451
rect 29733 20411 29791 20417
rect 15948 20352 16804 20380
rect 15948 20321 15976 20352
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 20257 20383 20315 20389
rect 20257 20380 20269 20383
rect 17920 20352 20269 20380
rect 17920 20340 17926 20352
rect 20257 20349 20269 20352
rect 20303 20349 20315 20383
rect 30006 20380 30012 20392
rect 29967 20352 30012 20380
rect 20257 20343 20315 20349
rect 30006 20340 30012 20352
rect 30064 20340 30070 20392
rect 15933 20315 15991 20321
rect 15933 20281 15945 20315
rect 15979 20281 15991 20315
rect 18046 20312 18052 20324
rect 18007 20284 18052 20312
rect 15933 20275 15991 20281
rect 18046 20272 18052 20284
rect 18104 20272 18110 20324
rect 25774 20272 25780 20324
rect 25832 20312 25838 20324
rect 27430 20312 27436 20324
rect 25832 20284 27436 20312
rect 25832 20272 25838 20284
rect 27430 20272 27436 20284
rect 27488 20272 27494 20324
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 18693 20247 18751 20253
rect 18693 20244 18705 20247
rect 18288 20216 18705 20244
rect 18288 20204 18294 20216
rect 18693 20213 18705 20216
rect 18739 20213 18751 20247
rect 18693 20207 18751 20213
rect 28166 20204 28172 20256
rect 28224 20244 28230 20256
rect 28353 20247 28411 20253
rect 28353 20244 28365 20247
rect 28224 20216 28365 20244
rect 28224 20204 28230 20216
rect 28353 20213 28365 20216
rect 28399 20213 28411 20247
rect 28353 20207 28411 20213
rect 1104 20154 30820 20176
rect 1104 20102 5915 20154
rect 5967 20102 5979 20154
rect 6031 20102 6043 20154
rect 6095 20102 6107 20154
rect 6159 20102 6171 20154
rect 6223 20102 15846 20154
rect 15898 20102 15910 20154
rect 15962 20102 15974 20154
rect 16026 20102 16038 20154
rect 16090 20102 16102 20154
rect 16154 20102 25776 20154
rect 25828 20102 25840 20154
rect 25892 20102 25904 20154
rect 25956 20102 25968 20154
rect 26020 20102 26032 20154
rect 26084 20102 30820 20154
rect 1104 20080 30820 20102
rect 2130 20040 2136 20052
rect 2091 20012 2136 20040
rect 2130 20000 2136 20012
rect 2188 20000 2194 20052
rect 16482 20000 16488 20052
rect 16540 20040 16546 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16540 20012 16865 20040
rect 16540 20000 16546 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 19392 20012 23152 20040
rect 19392 20000 19398 20012
rect 9674 19932 9680 19984
rect 9732 19972 9738 19984
rect 17589 19975 17647 19981
rect 17589 19972 17601 19975
rect 9732 19944 17601 19972
rect 9732 19932 9738 19944
rect 17589 19941 17601 19944
rect 17635 19941 17647 19975
rect 23124 19972 23152 20012
rect 23198 20000 23204 20052
rect 23256 20040 23262 20052
rect 23293 20043 23351 20049
rect 23293 20040 23305 20043
rect 23256 20012 23305 20040
rect 23256 20000 23262 20012
rect 23293 20009 23305 20012
rect 23339 20040 23351 20043
rect 24026 20040 24032 20052
rect 23339 20012 24032 20040
rect 23339 20009 23351 20012
rect 23293 20003 23351 20009
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 28629 20043 28687 20049
rect 28629 20009 28641 20043
rect 28675 20040 28687 20043
rect 28718 20040 28724 20052
rect 28675 20012 28724 20040
rect 28675 20009 28687 20012
rect 28629 20003 28687 20009
rect 28718 20000 28724 20012
rect 28776 20000 28782 20052
rect 28994 20000 29000 20052
rect 29052 20040 29058 20052
rect 30009 20043 30067 20049
rect 30009 20040 30021 20043
rect 29052 20012 30021 20040
rect 29052 20000 29058 20012
rect 30009 20009 30021 20012
rect 30055 20040 30067 20043
rect 30282 20040 30288 20052
rect 30055 20012 30288 20040
rect 30055 20009 30067 20012
rect 30009 20003 30067 20009
rect 30282 20000 30288 20012
rect 30340 20000 30346 20052
rect 29454 19972 29460 19984
rect 23124 19944 29460 19972
rect 17589 19935 17647 19941
rect 29454 19932 29460 19944
rect 29512 19932 29518 19984
rect 29822 19932 29828 19984
rect 29880 19972 29886 19984
rect 30190 19972 30196 19984
rect 29880 19944 30196 19972
rect 29880 19932 29886 19944
rect 30190 19932 30196 19944
rect 30248 19932 30254 19984
rect 23474 19864 23480 19916
rect 23532 19904 23538 19916
rect 24118 19904 24124 19916
rect 23532 19876 24124 19904
rect 23532 19864 23538 19876
rect 24118 19864 24124 19876
rect 24176 19864 24182 19916
rect 25958 19904 25964 19916
rect 25056 19876 25964 19904
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19836 1455 19839
rect 2130 19836 2136 19848
rect 1443 19808 2136 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 2130 19796 2136 19808
rect 2188 19796 2194 19848
rect 2314 19836 2320 19848
rect 2275 19808 2320 19836
rect 2314 19796 2320 19808
rect 2372 19796 2378 19848
rect 16482 19836 16488 19848
rect 16443 19808 16488 19836
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 16666 19836 16672 19848
rect 16627 19808 16672 19836
rect 16666 19796 16672 19808
rect 16724 19796 16730 19848
rect 17770 19836 17776 19848
rect 17731 19808 17776 19836
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 18230 19836 18236 19848
rect 18191 19808 18236 19836
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 19242 19796 19248 19848
rect 19300 19836 19306 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 19300 19808 20177 19836
rect 19300 19796 19306 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 20622 19836 20628 19848
rect 20395 19808 20628 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 21913 19839 21971 19845
rect 21913 19805 21925 19839
rect 21959 19836 21971 19839
rect 22462 19836 22468 19848
rect 21959 19808 22468 19836
rect 21959 19805 21971 19808
rect 21913 19799 21971 19805
rect 22462 19796 22468 19808
rect 22520 19796 22526 19848
rect 24578 19836 24584 19848
rect 24539 19808 24584 19836
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 24854 19836 24860 19848
rect 24815 19808 24860 19836
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 25056 19845 25084 19876
rect 25958 19864 25964 19876
rect 26016 19864 26022 19916
rect 26050 19864 26056 19916
rect 26108 19904 26114 19916
rect 27062 19904 27068 19916
rect 26108 19876 27068 19904
rect 26108 19864 26114 19876
rect 27062 19864 27068 19876
rect 27120 19864 27126 19916
rect 28258 19864 28264 19916
rect 28316 19904 28322 19916
rect 31754 19904 31760 19916
rect 28316 19876 31760 19904
rect 28316 19864 28322 19876
rect 31754 19864 31760 19876
rect 31812 19864 31818 19916
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19805 25099 19839
rect 25041 19799 25099 19805
rect 25130 19796 25136 19848
rect 25188 19836 25194 19848
rect 27246 19836 27252 19848
rect 25188 19808 27252 19836
rect 25188 19796 25194 19808
rect 27246 19796 27252 19808
rect 27304 19796 27310 19848
rect 27982 19796 27988 19848
rect 28040 19836 28046 19848
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 28040 19808 28457 19836
rect 28040 19796 28046 19808
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 29822 19836 29828 19848
rect 29783 19808 29828 19836
rect 28445 19799 28503 19805
rect 29822 19796 29828 19808
rect 29880 19796 29886 19848
rect 20533 19771 20591 19777
rect 20533 19737 20545 19771
rect 20579 19768 20591 19771
rect 21450 19768 21456 19780
rect 20579 19740 21456 19768
rect 20579 19737 20591 19740
rect 20533 19731 20591 19737
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 22180 19771 22238 19777
rect 22180 19737 22192 19771
rect 22226 19768 22238 19771
rect 22922 19768 22928 19780
rect 22226 19740 22928 19768
rect 22226 19737 22238 19740
rect 22180 19731 22238 19737
rect 22922 19728 22928 19740
rect 22980 19728 22986 19780
rect 25498 19728 25504 19780
rect 25556 19768 25562 19780
rect 26786 19768 26792 19780
rect 25556 19740 26792 19768
rect 25556 19728 25562 19740
rect 26786 19728 26792 19740
rect 26844 19728 26850 19780
rect 27798 19728 27804 19780
rect 27856 19768 27862 19780
rect 28261 19771 28319 19777
rect 28261 19768 28273 19771
rect 27856 19740 28273 19768
rect 27856 19728 27862 19740
rect 28261 19737 28273 19740
rect 28307 19737 28319 19771
rect 30374 19768 30380 19780
rect 28261 19731 28319 19737
rect 28920 19740 30380 19768
rect 1578 19700 1584 19712
rect 1539 19672 1584 19700
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 24210 19700 24216 19712
rect 20772 19672 24216 19700
rect 20772 19660 20778 19672
rect 24210 19660 24216 19672
rect 24268 19660 24274 19712
rect 24394 19700 24400 19712
rect 24355 19672 24400 19700
rect 24394 19660 24400 19672
rect 24452 19660 24458 19712
rect 28920 19700 28948 19740
rect 30374 19728 30380 19740
rect 30432 19728 30438 19780
rect 29178 19700 29184 19712
rect 28920 19672 29184 19700
rect 29178 19660 29184 19672
rect 29236 19660 29242 19712
rect 1104 19610 30820 19632
rect 1104 19558 10880 19610
rect 10932 19558 10944 19610
rect 10996 19558 11008 19610
rect 11060 19558 11072 19610
rect 11124 19558 11136 19610
rect 11188 19558 20811 19610
rect 20863 19558 20875 19610
rect 20927 19558 20939 19610
rect 20991 19558 21003 19610
rect 21055 19558 21067 19610
rect 21119 19558 30820 19610
rect 1104 19536 30820 19558
rect 2130 19496 2136 19508
rect 2091 19468 2136 19496
rect 2130 19456 2136 19468
rect 2188 19456 2194 19508
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 17313 19499 17371 19505
rect 17313 19496 17325 19499
rect 16724 19468 17325 19496
rect 16724 19456 16730 19468
rect 17313 19465 17325 19468
rect 17359 19465 17371 19499
rect 22922 19496 22928 19508
rect 22883 19468 22928 19496
rect 17313 19459 17371 19465
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 24210 19456 24216 19508
rect 24268 19496 24274 19508
rect 27599 19499 27657 19505
rect 27599 19496 27611 19499
rect 24268 19468 27611 19496
rect 24268 19456 24274 19468
rect 27599 19465 27611 19468
rect 27645 19465 27657 19499
rect 27599 19459 27657 19465
rect 28077 19499 28135 19505
rect 28077 19465 28089 19499
rect 28123 19496 28135 19499
rect 28258 19496 28264 19508
rect 28123 19468 28264 19496
rect 28123 19465 28135 19468
rect 28077 19459 28135 19465
rect 28258 19456 28264 19468
rect 28316 19456 28322 19508
rect 28721 19499 28779 19505
rect 28721 19465 28733 19499
rect 28767 19496 28779 19499
rect 29178 19496 29184 19508
rect 28767 19468 29184 19496
rect 28767 19465 28779 19468
rect 28721 19459 28779 19465
rect 29178 19456 29184 19468
rect 29236 19456 29242 19508
rect 29917 19499 29975 19505
rect 29917 19465 29929 19499
rect 29963 19496 29975 19499
rect 31202 19496 31208 19508
rect 29963 19468 31208 19496
rect 29963 19465 29975 19468
rect 29917 19459 29975 19465
rect 31202 19456 31208 19468
rect 31260 19456 31266 19508
rect 17681 19431 17739 19437
rect 17681 19397 17693 19431
rect 17727 19428 17739 19431
rect 17862 19428 17868 19440
rect 17727 19400 17868 19428
rect 17727 19397 17739 19400
rect 17681 19391 17739 19397
rect 17862 19388 17868 19400
rect 17920 19428 17926 19440
rect 17920 19400 19104 19428
rect 17920 19388 17926 19400
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19360 2375 19363
rect 17773 19363 17831 19369
rect 2363 19332 11008 19360
rect 2363 19329 2375 19332
rect 2317 19323 2375 19329
rect 10980 19292 11008 19332
rect 17773 19329 17785 19363
rect 17819 19360 17831 19363
rect 18230 19360 18236 19372
rect 17819 19332 18236 19360
rect 17819 19329 17831 19332
rect 17773 19323 17831 19329
rect 18230 19320 18236 19332
rect 18288 19360 18294 19372
rect 18524 19369 18552 19400
rect 18509 19363 18567 19369
rect 18288 19332 18460 19360
rect 18288 19320 18294 19332
rect 17865 19295 17923 19301
rect 10980 19264 12434 19292
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 12406 19156 12434 19264
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 18046 19292 18052 19304
rect 17911 19264 18052 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18432 19292 18460 19332
rect 18509 19329 18521 19363
rect 18555 19329 18567 19363
rect 18509 19323 18567 19329
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18785 19363 18843 19369
rect 18785 19360 18797 19363
rect 18656 19332 18797 19360
rect 18656 19320 18662 19332
rect 18785 19329 18797 19332
rect 18831 19329 18843 19363
rect 18785 19323 18843 19329
rect 18966 19292 18972 19304
rect 18432 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19076 19292 19104 19400
rect 19242 19388 19248 19440
rect 19300 19428 19306 19440
rect 19300 19400 20116 19428
rect 19300 19388 19306 19400
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19360 19211 19363
rect 19610 19360 19616 19372
rect 19199 19332 19616 19360
rect 19199 19329 19211 19332
rect 19153 19323 19211 19329
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 20088 19369 20116 19400
rect 25406 19388 25412 19440
rect 25464 19428 25470 19440
rect 25464 19400 25820 19428
rect 25464 19388 25470 19400
rect 25792 19372 25820 19400
rect 27430 19388 27436 19440
rect 27488 19428 27494 19440
rect 27893 19431 27951 19437
rect 27893 19428 27905 19431
rect 27488 19400 27905 19428
rect 27488 19388 27494 19400
rect 27893 19397 27905 19400
rect 27939 19397 27951 19431
rect 27893 19391 27951 19397
rect 28166 19388 28172 19440
rect 28224 19428 28230 19440
rect 28994 19428 29000 19440
rect 28224 19400 29000 19428
rect 28224 19388 28230 19400
rect 28994 19388 29000 19400
rect 29052 19428 29058 19440
rect 30006 19428 30012 19440
rect 29052 19400 30012 19428
rect 29052 19388 29058 19400
rect 30006 19388 30012 19400
rect 30064 19388 30070 19440
rect 19889 19363 19947 19369
rect 19889 19360 19901 19363
rect 19720 19332 19901 19360
rect 19720 19292 19748 19332
rect 19889 19329 19901 19332
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 20073 19363 20131 19369
rect 20073 19329 20085 19363
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 21266 19360 21272 19372
rect 20303 19332 21272 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19360 23167 19363
rect 24394 19360 24400 19372
rect 23155 19332 24400 19360
rect 23155 19329 23167 19332
rect 23109 19323 23167 19329
rect 24394 19320 24400 19332
rect 24452 19320 24458 19372
rect 25590 19320 25596 19372
rect 25648 19360 25654 19372
rect 25685 19363 25743 19369
rect 25685 19360 25697 19363
rect 25648 19332 25697 19360
rect 25648 19320 25654 19332
rect 25685 19329 25697 19332
rect 25731 19329 25743 19363
rect 25685 19323 25743 19329
rect 25774 19320 25780 19372
rect 25832 19360 25838 19372
rect 25869 19363 25927 19369
rect 25869 19360 25881 19363
rect 25832 19332 25881 19360
rect 25832 19320 25838 19332
rect 25869 19329 25881 19332
rect 25915 19329 25927 19363
rect 25869 19323 25927 19329
rect 26145 19363 26203 19369
rect 26145 19329 26157 19363
rect 26191 19329 26203 19363
rect 26145 19323 26203 19329
rect 26329 19363 26387 19369
rect 26329 19329 26341 19363
rect 26375 19360 26387 19363
rect 26694 19360 26700 19372
rect 26375 19332 26700 19360
rect 26375 19329 26387 19332
rect 26329 19323 26387 19329
rect 19076 19264 19748 19292
rect 23198 19252 23204 19304
rect 23256 19292 23262 19304
rect 23385 19295 23443 19301
rect 23385 19292 23397 19295
rect 23256 19264 23397 19292
rect 23256 19252 23262 19264
rect 23385 19261 23397 19264
rect 23431 19261 23443 19295
rect 23385 19255 23443 19261
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 26160 19292 26188 19323
rect 26694 19320 26700 19332
rect 26752 19320 26758 19372
rect 28902 19360 28908 19372
rect 28863 19332 28908 19360
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29178 19320 29184 19372
rect 29236 19360 29242 19372
rect 29638 19360 29644 19372
rect 29236 19332 29644 19360
rect 29236 19320 29242 19332
rect 29638 19320 29644 19332
rect 29696 19360 29702 19372
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 29696 19332 29745 19360
rect 29696 19320 29702 19332
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 25188 19264 26188 19292
rect 25188 19252 25194 19264
rect 23293 19227 23351 19233
rect 23293 19193 23305 19227
rect 23339 19224 23351 19227
rect 23658 19224 23664 19236
rect 23339 19196 23664 19224
rect 23339 19193 23351 19196
rect 23293 19187 23351 19193
rect 23658 19184 23664 19196
rect 23716 19224 23722 19236
rect 24026 19224 24032 19236
rect 23716 19196 24032 19224
rect 23716 19184 23722 19196
rect 24026 19184 24032 19196
rect 24084 19184 24090 19236
rect 25866 19184 25872 19236
rect 25924 19224 25930 19236
rect 28902 19224 28908 19236
rect 25924 19196 28908 19224
rect 25924 19184 25930 19196
rect 28902 19184 28908 19196
rect 28960 19184 28966 19236
rect 29454 19224 29460 19236
rect 29415 19196 29460 19224
rect 29454 19184 29460 19196
rect 29512 19184 29518 19236
rect 23198 19156 23204 19168
rect 12406 19128 23204 19156
rect 23198 19116 23204 19128
rect 23256 19116 23262 19168
rect 1104 19066 30820 19088
rect 1104 19014 5915 19066
rect 5967 19014 5979 19066
rect 6031 19014 6043 19066
rect 6095 19014 6107 19066
rect 6159 19014 6171 19066
rect 6223 19014 15846 19066
rect 15898 19014 15910 19066
rect 15962 19014 15974 19066
rect 16026 19014 16038 19066
rect 16090 19014 16102 19066
rect 16154 19014 25776 19066
rect 25828 19014 25840 19066
rect 25892 19014 25904 19066
rect 25956 19014 25968 19066
rect 26020 19014 26032 19066
rect 26084 19014 30820 19066
rect 31570 19048 31576 19100
rect 31628 19088 31634 19100
rect 31754 19088 31760 19100
rect 31628 19060 31760 19088
rect 31628 19048 31634 19060
rect 31754 19048 31760 19060
rect 31812 19048 31818 19100
rect 1104 18992 30820 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 1452 18924 2329 18952
rect 1452 18912 1458 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 6886 18924 22094 18952
rect 6886 18884 6914 18924
rect 1872 18856 6914 18884
rect 22066 18884 22094 18924
rect 23198 18912 23204 18964
rect 23256 18952 23262 18964
rect 28353 18955 28411 18961
rect 28353 18952 28365 18955
rect 23256 18924 28365 18952
rect 23256 18912 23262 18924
rect 28353 18921 28365 18924
rect 28399 18921 28411 18955
rect 28353 18915 28411 18921
rect 29546 18912 29552 18964
rect 29604 18952 29610 18964
rect 29917 18955 29975 18961
rect 29917 18952 29929 18955
rect 29604 18924 29929 18952
rect 29604 18912 29610 18924
rect 29917 18921 29929 18924
rect 29963 18921 29975 18955
rect 29917 18915 29975 18921
rect 25406 18884 25412 18896
rect 22066 18856 25412 18884
rect 1872 18757 1900 18856
rect 25406 18844 25412 18856
rect 25464 18844 25470 18896
rect 26602 18844 26608 18896
rect 26660 18884 26666 18896
rect 26973 18887 27031 18893
rect 26973 18884 26985 18887
rect 26660 18856 26985 18884
rect 26660 18844 26666 18856
rect 26973 18853 26985 18856
rect 27019 18884 27031 18887
rect 27522 18884 27528 18896
rect 27019 18856 27528 18884
rect 27019 18853 27031 18856
rect 26973 18847 27031 18853
rect 27522 18844 27528 18856
rect 27580 18844 27586 18896
rect 28166 18844 28172 18896
rect 28224 18884 28230 18896
rect 28442 18884 28448 18896
rect 28224 18856 28448 18884
rect 28224 18844 28230 18856
rect 28442 18844 28448 18856
rect 28500 18844 28506 18896
rect 19334 18816 19340 18828
rect 6886 18788 19340 18816
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18717 1915 18751
rect 1857 18711 1915 18717
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18748 2559 18751
rect 6886 18748 6914 18788
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 22462 18776 22468 18828
rect 22520 18816 22526 18828
rect 25593 18819 25651 18825
rect 25593 18816 25605 18819
rect 22520 18788 25605 18816
rect 22520 18776 22526 18788
rect 25593 18785 25605 18788
rect 25639 18785 25651 18819
rect 25593 18779 25651 18785
rect 27982 18776 27988 18828
rect 28040 18816 28046 18828
rect 28905 18819 28963 18825
rect 28040 18788 28764 18816
rect 28040 18776 28046 18788
rect 24578 18748 24584 18760
rect 2547 18720 6914 18748
rect 24539 18720 24584 18748
rect 2547 18717 2559 18720
rect 2501 18711 2559 18717
rect 24578 18708 24584 18720
rect 24636 18708 24642 18760
rect 24854 18748 24860 18760
rect 24815 18720 24860 18748
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18748 25099 18751
rect 28626 18748 28632 18760
rect 25087 18720 26004 18748
rect 28587 18720 28632 18748
rect 25087 18717 25099 18720
rect 25041 18711 25099 18717
rect 25976 18692 26004 18720
rect 28626 18708 28632 18720
rect 28684 18708 28690 18760
rect 28736 18748 28764 18788
rect 28905 18785 28917 18819
rect 28951 18816 28963 18819
rect 28994 18816 29000 18828
rect 28951 18788 29000 18816
rect 28951 18785 28963 18788
rect 28905 18779 28963 18785
rect 28994 18776 29000 18788
rect 29052 18776 29058 18828
rect 29733 18751 29791 18757
rect 29733 18748 29745 18751
rect 28736 18720 29745 18748
rect 29733 18717 29745 18720
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 1486 18640 1492 18692
rect 1544 18680 1550 18692
rect 1544 18652 6914 18680
rect 1544 18640 1550 18652
rect 1394 18572 1400 18624
rect 1452 18612 1458 18624
rect 1673 18615 1731 18621
rect 1673 18612 1685 18615
rect 1452 18584 1685 18612
rect 1452 18572 1458 18584
rect 1673 18581 1685 18584
rect 1719 18581 1731 18615
rect 6886 18612 6914 18652
rect 25682 18640 25688 18692
rect 25740 18680 25746 18692
rect 25838 18683 25896 18689
rect 25838 18680 25850 18683
rect 25740 18652 25850 18680
rect 25740 18640 25746 18652
rect 25838 18649 25850 18652
rect 25884 18649 25896 18683
rect 25838 18643 25896 18649
rect 25958 18640 25964 18692
rect 26016 18640 26022 18692
rect 28442 18640 28448 18692
rect 28500 18680 28506 18692
rect 29549 18683 29607 18689
rect 29549 18680 29561 18683
rect 28500 18652 29561 18680
rect 28500 18640 28506 18652
rect 29549 18649 29561 18652
rect 29595 18649 29607 18683
rect 29549 18643 29607 18649
rect 21726 18612 21732 18624
rect 6886 18584 21732 18612
rect 1673 18575 1731 18581
rect 21726 18572 21732 18584
rect 21784 18572 21790 18624
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24397 18615 24455 18621
rect 24397 18612 24409 18615
rect 23900 18584 24409 18612
rect 23900 18572 23906 18584
rect 24397 18581 24409 18584
rect 24443 18581 24455 18615
rect 24397 18575 24455 18581
rect 28813 18615 28871 18621
rect 28813 18581 28825 18615
rect 28859 18612 28871 18615
rect 31754 18612 31760 18624
rect 28859 18584 31760 18612
rect 28859 18581 28871 18584
rect 28813 18575 28871 18581
rect 31754 18572 31760 18584
rect 31812 18572 31818 18624
rect 1104 18522 30820 18544
rect 1104 18470 10880 18522
rect 10932 18470 10944 18522
rect 10996 18470 11008 18522
rect 11060 18470 11072 18522
rect 11124 18470 11136 18522
rect 11188 18470 20811 18522
rect 20863 18470 20875 18522
rect 20927 18470 20939 18522
rect 20991 18470 21003 18522
rect 21055 18470 21067 18522
rect 21119 18470 30820 18522
rect 1104 18448 30820 18470
rect 22830 18368 22836 18420
rect 22888 18408 22894 18420
rect 23201 18411 23259 18417
rect 23201 18408 23213 18411
rect 22888 18380 23213 18408
rect 22888 18368 22894 18380
rect 23201 18377 23213 18380
rect 23247 18377 23259 18411
rect 23201 18371 23259 18377
rect 28350 18368 28356 18420
rect 28408 18408 28414 18420
rect 28629 18411 28687 18417
rect 28629 18408 28641 18411
rect 28408 18380 28641 18408
rect 28408 18368 28414 18380
rect 28629 18377 28641 18380
rect 28675 18377 28687 18411
rect 28629 18371 28687 18377
rect 29733 18411 29791 18417
rect 29733 18377 29745 18411
rect 29779 18408 29791 18411
rect 31662 18408 31668 18420
rect 29779 18380 31668 18408
rect 29779 18377 29791 18380
rect 29733 18371 29791 18377
rect 31662 18368 31668 18380
rect 31720 18368 31726 18420
rect 22462 18340 22468 18352
rect 21836 18312 22468 18340
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 20714 18272 20720 18284
rect 2363 18244 20720 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 21836 18281 21864 18312
rect 22462 18300 22468 18312
rect 22520 18300 22526 18352
rect 24118 18300 24124 18352
rect 24176 18300 24182 18352
rect 27982 18300 27988 18352
rect 28040 18340 28046 18352
rect 28445 18343 28503 18349
rect 28445 18340 28457 18343
rect 28040 18312 28457 18340
rect 28040 18300 28046 18312
rect 28445 18309 28457 18312
rect 28491 18309 28503 18343
rect 28445 18303 28503 18309
rect 29362 18300 29368 18352
rect 29420 18340 29426 18352
rect 29549 18343 29607 18349
rect 29549 18340 29561 18343
rect 29420 18312 29561 18340
rect 29420 18300 29426 18312
rect 29549 18309 29561 18312
rect 29595 18309 29607 18343
rect 29549 18303 29607 18309
rect 21821 18275 21879 18281
rect 21821 18241 21833 18275
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22088 18275 22146 18281
rect 22088 18241 22100 18275
rect 22134 18272 22146 18275
rect 22370 18272 22376 18284
rect 22134 18244 22376 18272
rect 22134 18241 22146 18244
rect 22088 18235 22146 18241
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 23842 18272 23848 18284
rect 23803 18244 23848 18272
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 24026 18272 24032 18284
rect 23987 18244 24032 18272
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 24136 18272 24164 18300
rect 24762 18272 24768 18284
rect 24136 18244 24768 18272
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 24854 18232 24860 18284
rect 24912 18272 24918 18284
rect 25501 18275 25559 18281
rect 25501 18272 25513 18275
rect 24912 18244 25513 18272
rect 24912 18232 24918 18244
rect 25501 18241 25513 18244
rect 25547 18241 25559 18275
rect 28258 18272 28264 18284
rect 28219 18244 28264 18272
rect 25501 18235 25559 18241
rect 28258 18232 28264 18244
rect 28316 18232 28322 18284
rect 28994 18232 29000 18284
rect 29052 18272 29058 18284
rect 29825 18275 29883 18281
rect 29825 18272 29837 18275
rect 29052 18244 29837 18272
rect 29052 18232 29058 18244
rect 29825 18241 29837 18244
rect 29871 18241 29883 18275
rect 29825 18235 29883 18241
rect 23106 18164 23112 18216
rect 23164 18204 23170 18216
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 23164 18176 24133 18204
rect 23164 18164 23170 18176
rect 23860 18148 23888 18176
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 24121 18167 24179 18173
rect 25130 18164 25136 18216
rect 25188 18204 25194 18216
rect 25225 18207 25283 18213
rect 25225 18204 25237 18207
rect 25188 18176 25237 18204
rect 25188 18164 25194 18176
rect 25225 18173 25237 18176
rect 25271 18173 25283 18207
rect 25958 18204 25964 18216
rect 25225 18167 25283 18173
rect 25332 18176 25964 18204
rect 1578 18136 1584 18148
rect 1539 18108 1584 18136
rect 1578 18096 1584 18108
rect 1636 18096 1642 18148
rect 23842 18096 23848 18148
rect 23900 18096 23906 18148
rect 25332 18136 25360 18176
rect 25958 18164 25964 18176
rect 26016 18164 26022 18216
rect 27338 18164 27344 18216
rect 27396 18204 27402 18216
rect 31018 18204 31024 18216
rect 27396 18176 31024 18204
rect 27396 18164 27402 18176
rect 31018 18164 31024 18176
rect 31076 18164 31082 18216
rect 25240 18108 25360 18136
rect 25240 18080 25268 18108
rect 25406 18096 25412 18148
rect 25464 18136 25470 18148
rect 29273 18139 29331 18145
rect 29273 18136 29285 18139
rect 25464 18108 29285 18136
rect 25464 18096 25470 18108
rect 29273 18105 29285 18108
rect 29319 18105 29331 18139
rect 29273 18099 29331 18105
rect 29914 18096 29920 18148
rect 29972 18136 29978 18148
rect 30282 18136 30288 18148
rect 29972 18108 30288 18136
rect 29972 18096 29978 18108
rect 30282 18096 30288 18108
rect 30340 18096 30346 18148
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 2133 18071 2191 18077
rect 2133 18068 2145 18071
rect 1452 18040 2145 18068
rect 1452 18028 1458 18040
rect 2133 18037 2145 18040
rect 2179 18037 2191 18071
rect 2133 18031 2191 18037
rect 18782 18028 18788 18080
rect 18840 18068 18846 18080
rect 19518 18068 19524 18080
rect 18840 18040 19524 18068
rect 18840 18028 18846 18040
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 23658 18068 23664 18080
rect 23619 18040 23664 18068
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 24210 18028 24216 18080
rect 24268 18068 24274 18080
rect 24578 18068 24584 18080
rect 24268 18040 24584 18068
rect 24268 18028 24274 18040
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 25222 18028 25228 18080
rect 25280 18028 25286 18080
rect 29362 18028 29368 18080
rect 29420 18068 29426 18080
rect 29822 18068 29828 18080
rect 29420 18040 29828 18068
rect 29420 18028 29426 18040
rect 29822 18028 29828 18040
rect 29880 18028 29886 18080
rect 1104 17978 30820 18000
rect 1104 17926 5915 17978
rect 5967 17926 5979 17978
rect 6031 17926 6043 17978
rect 6095 17926 6107 17978
rect 6159 17926 6171 17978
rect 6223 17926 15846 17978
rect 15898 17926 15910 17978
rect 15962 17926 15974 17978
rect 16026 17926 16038 17978
rect 16090 17926 16102 17978
rect 16154 17926 25776 17978
rect 25828 17926 25840 17978
rect 25892 17926 25904 17978
rect 25956 17926 25968 17978
rect 26020 17926 26032 17978
rect 26084 17926 30820 17978
rect 1104 17904 30820 17926
rect 22002 17824 22008 17876
rect 22060 17864 22066 17876
rect 22738 17864 22744 17876
rect 22060 17836 22744 17864
rect 22060 17824 22066 17836
rect 22738 17824 22744 17836
rect 22796 17824 22802 17876
rect 23842 17864 23848 17876
rect 23803 17836 23848 17864
rect 23842 17824 23848 17836
rect 23900 17824 23906 17876
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24949 17867 25007 17873
rect 24949 17864 24961 17867
rect 24084 17836 24961 17864
rect 24084 17824 24090 17836
rect 24949 17833 24961 17836
rect 24995 17833 25007 17867
rect 25682 17864 25688 17876
rect 25643 17836 25688 17864
rect 24949 17827 25007 17833
rect 25682 17824 25688 17836
rect 25740 17824 25746 17876
rect 28626 17824 28632 17876
rect 28684 17864 28690 17876
rect 28813 17867 28871 17873
rect 28813 17864 28825 17867
rect 28684 17836 28825 17864
rect 28684 17824 28690 17836
rect 28813 17833 28825 17836
rect 28859 17833 28871 17867
rect 28813 17827 28871 17833
rect 28169 17799 28227 17805
rect 28169 17765 28181 17799
rect 28215 17796 28227 17799
rect 29270 17796 29276 17808
rect 28215 17768 29276 17796
rect 28215 17765 28227 17768
rect 28169 17759 28227 17765
rect 29270 17756 29276 17768
rect 29328 17756 29334 17808
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 21085 17731 21143 17737
rect 21085 17728 21097 17731
rect 19484 17700 21097 17728
rect 19484 17688 19490 17700
rect 21085 17697 21097 17700
rect 21131 17697 21143 17731
rect 21085 17691 21143 17697
rect 26145 17731 26203 17737
rect 26145 17697 26157 17731
rect 26191 17728 26203 17731
rect 26602 17728 26608 17740
rect 26191 17700 26608 17728
rect 26191 17697 26203 17700
rect 26145 17691 26203 17697
rect 26602 17688 26608 17700
rect 26660 17688 26666 17740
rect 28626 17688 28632 17740
rect 28684 17728 28690 17740
rect 30926 17728 30932 17740
rect 28684 17700 30932 17728
rect 28684 17688 28690 17700
rect 30926 17688 30932 17700
rect 30984 17688 30990 17740
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17620 1458 17672
rect 19610 17660 19616 17672
rect 19571 17632 19616 17660
rect 19610 17620 19616 17632
rect 19668 17620 19674 17672
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17660 19947 17663
rect 20346 17660 20352 17672
rect 19935 17632 20352 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17660 20775 17663
rect 21450 17660 21456 17672
rect 20763 17632 21456 17660
rect 20763 17629 20775 17632
rect 20717 17623 20775 17629
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22462 17660 22468 17672
rect 22423 17632 22468 17660
rect 22462 17620 22468 17632
rect 22520 17620 22526 17672
rect 22732 17663 22790 17669
rect 22732 17629 22744 17663
rect 22778 17660 22790 17663
rect 23658 17660 23664 17672
rect 22778 17632 23664 17660
rect 22778 17629 22790 17632
rect 22732 17623 22790 17629
rect 23658 17620 23664 17632
rect 23716 17620 23722 17672
rect 25590 17620 25596 17672
rect 25648 17660 25654 17672
rect 25869 17663 25927 17669
rect 25869 17660 25881 17663
rect 25648 17632 25881 17660
rect 25648 17620 25654 17632
rect 25869 17629 25881 17632
rect 25915 17629 25927 17663
rect 26050 17660 26056 17672
rect 26011 17632 26056 17660
rect 25869 17623 25927 17629
rect 26050 17620 26056 17632
rect 26108 17660 26114 17672
rect 26234 17660 26240 17672
rect 26108 17632 26240 17660
rect 26108 17620 26114 17632
rect 26234 17620 26240 17632
rect 26292 17620 26298 17672
rect 28350 17660 28356 17672
rect 28311 17632 28356 17660
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 28997 17663 29055 17669
rect 28997 17660 29009 17663
rect 28868 17632 29009 17660
rect 28868 17620 28874 17632
rect 28997 17629 29009 17632
rect 29043 17629 29055 17663
rect 29914 17660 29920 17672
rect 29875 17632 29920 17660
rect 28997 17623 29055 17629
rect 29914 17620 29920 17632
rect 29972 17620 29978 17672
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 18966 17592 18972 17604
rect 18656 17564 18972 17592
rect 18656 17552 18662 17564
rect 18966 17552 18972 17564
rect 19024 17592 19030 17604
rect 19797 17595 19855 17601
rect 19797 17592 19809 17595
rect 19024 17564 19809 17592
rect 19024 17552 19030 17564
rect 19797 17561 19809 17564
rect 19843 17561 19855 17595
rect 19797 17555 19855 17561
rect 20901 17595 20959 17601
rect 20901 17561 20913 17595
rect 20947 17592 20959 17595
rect 22830 17592 22836 17604
rect 20947 17564 22836 17592
rect 20947 17561 20959 17564
rect 20901 17555 20959 17561
rect 22830 17552 22836 17564
rect 22888 17552 22894 17604
rect 24857 17595 24915 17601
rect 24857 17561 24869 17595
rect 24903 17592 24915 17595
rect 26068 17592 26096 17620
rect 24903 17564 26096 17592
rect 24903 17561 24915 17564
rect 24857 17555 24915 17561
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19702 17524 19708 17536
rect 19475 17496 19708 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 28902 17484 28908 17536
rect 28960 17524 28966 17536
rect 30009 17527 30067 17533
rect 30009 17524 30021 17527
rect 28960 17496 30021 17524
rect 28960 17484 28966 17496
rect 30009 17493 30021 17496
rect 30055 17493 30067 17527
rect 30009 17487 30067 17493
rect 1104 17434 30820 17456
rect 1104 17382 10880 17434
rect 10932 17382 10944 17434
rect 10996 17382 11008 17434
rect 11060 17382 11072 17434
rect 11124 17382 11136 17434
rect 11188 17382 20811 17434
rect 20863 17382 20875 17434
rect 20927 17382 20939 17434
rect 20991 17382 21003 17434
rect 21055 17382 21067 17434
rect 21119 17382 30820 17434
rect 1104 17360 30820 17382
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 21542 17320 21548 17332
rect 18104 17292 21548 17320
rect 18104 17280 18110 17292
rect 21542 17280 21548 17292
rect 21600 17280 21606 17332
rect 22370 17280 22376 17332
rect 22428 17320 22434 17332
rect 22465 17323 22523 17329
rect 22465 17320 22477 17323
rect 22428 17292 22477 17320
rect 22428 17280 22434 17292
rect 22465 17289 22477 17292
rect 22511 17289 22523 17323
rect 27522 17320 27528 17332
rect 27483 17292 27528 17320
rect 22465 17283 22523 17289
rect 27522 17280 27528 17292
rect 27580 17280 27586 17332
rect 27982 17280 27988 17332
rect 28040 17320 28046 17332
rect 28718 17320 28724 17332
rect 28040 17292 28724 17320
rect 28040 17280 28046 17292
rect 28718 17280 28724 17292
rect 28776 17280 28782 17332
rect 29178 17320 29184 17332
rect 29139 17292 29184 17320
rect 29178 17280 29184 17292
rect 29236 17280 29242 17332
rect 23382 17252 23388 17264
rect 18432 17224 19656 17252
rect 1397 17187 1455 17193
rect 1397 17153 1409 17187
rect 1443 17184 1455 17187
rect 2317 17187 2375 17193
rect 1443 17156 2176 17184
rect 1443 17153 1455 17156
rect 1397 17147 1455 17153
rect 2148 17057 2176 17156
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 2682 17184 2688 17196
rect 2363 17156 2688 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 17218 17144 17224 17196
rect 17276 17184 17282 17196
rect 18432 17193 18460 17224
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 17276 17156 17877 17184
rect 17276 17144 17282 17156
rect 17865 17153 17877 17156
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 18417 17187 18475 17193
rect 18417 17153 18429 17187
rect 18463 17153 18475 17187
rect 18598 17184 18604 17196
rect 18559 17156 18604 17184
rect 18417 17147 18475 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17184 19027 17187
rect 19518 17184 19524 17196
rect 19015 17156 19524 17184
rect 19015 17153 19027 17156
rect 18969 17147 19027 17153
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19628 17193 19656 17224
rect 19720 17224 23388 17252
rect 19720 17193 19748 17224
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 27430 17252 27436 17264
rect 24504 17224 27436 17252
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17153 19763 17187
rect 19886 17184 19892 17196
rect 19847 17156 19892 17184
rect 19705 17147 19763 17153
rect 18877 17119 18935 17125
rect 18877 17085 18889 17119
rect 18923 17116 18935 17119
rect 19334 17116 19340 17128
rect 18923 17088 19340 17116
rect 18923 17085 18935 17088
rect 18877 17079 18935 17085
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 19628 17116 19656 17147
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20714 17184 20720 17196
rect 20027 17156 20720 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20714 17144 20720 17156
rect 20772 17184 20778 17196
rect 21266 17184 21272 17196
rect 20772 17156 21272 17184
rect 20772 17144 20778 17156
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 22649 17187 22707 17193
rect 22649 17153 22661 17187
rect 22695 17184 22707 17187
rect 23845 17187 23903 17193
rect 23845 17184 23857 17187
rect 22695 17156 23857 17184
rect 22695 17153 22707 17156
rect 22649 17147 22707 17153
rect 23845 17153 23857 17156
rect 23891 17153 23903 17187
rect 23845 17147 23903 17153
rect 24029 17187 24087 17193
rect 24029 17153 24041 17187
rect 24075 17184 24087 17187
rect 24210 17184 24216 17196
rect 24075 17156 24216 17184
rect 24075 17153 24087 17156
rect 24029 17147 24087 17153
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 24504 17193 24532 17224
rect 27430 17212 27436 17224
rect 27488 17212 27494 17264
rect 28166 17212 28172 17264
rect 28224 17252 28230 17264
rect 28261 17255 28319 17261
rect 28261 17252 28273 17255
rect 28224 17224 28273 17252
rect 28224 17212 28230 17224
rect 28261 17221 28273 17224
rect 28307 17221 28319 17255
rect 28261 17215 28319 17221
rect 29917 17255 29975 17261
rect 29917 17221 29929 17255
rect 29963 17252 29975 17255
rect 30006 17252 30012 17264
rect 29963 17224 30012 17252
rect 29963 17221 29975 17224
rect 29917 17215 29975 17221
rect 30006 17212 30012 17224
rect 30064 17212 30070 17264
rect 24305 17187 24363 17193
rect 24305 17153 24317 17187
rect 24351 17153 24363 17187
rect 24305 17147 24363 17153
rect 24489 17187 24547 17193
rect 24489 17153 24501 17187
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 20346 17116 20352 17128
rect 19628 17088 20352 17116
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 22830 17076 22836 17128
rect 22888 17116 22894 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22888 17088 22937 17116
rect 22888 17076 22894 17088
rect 22925 17085 22937 17088
rect 22971 17085 22983 17119
rect 22925 17079 22983 17085
rect 24118 17076 24124 17128
rect 24176 17116 24182 17128
rect 24320 17116 24348 17147
rect 27062 17144 27068 17196
rect 27120 17184 27126 17196
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 27120 17156 27353 17184
rect 27120 17144 27126 17156
rect 27341 17153 27353 17156
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 28902 17144 28908 17196
rect 28960 17184 28966 17196
rect 29365 17187 29423 17193
rect 29365 17184 29377 17187
rect 28960 17156 29377 17184
rect 28960 17144 28966 17156
rect 29365 17153 29377 17156
rect 29411 17153 29423 17187
rect 29365 17147 29423 17153
rect 24176 17088 24348 17116
rect 27617 17119 27675 17125
rect 24176 17076 24182 17088
rect 27617 17085 27629 17119
rect 27663 17116 27675 17119
rect 27706 17116 27712 17128
rect 27663 17088 27712 17116
rect 27663 17085 27675 17088
rect 27617 17079 27675 17085
rect 27706 17076 27712 17088
rect 27764 17116 27770 17128
rect 28445 17119 28503 17125
rect 28445 17116 28457 17119
rect 27764 17088 28457 17116
rect 27764 17076 27770 17088
rect 28445 17085 28457 17088
rect 28491 17085 28503 17119
rect 28445 17079 28503 17085
rect 29178 17076 29184 17128
rect 29236 17116 29242 17128
rect 30098 17116 30104 17128
rect 29236 17088 30104 17116
rect 29236 17076 29242 17088
rect 30098 17076 30104 17088
rect 30156 17076 30162 17128
rect 2133 17051 2191 17057
rect 2133 17017 2145 17051
rect 2179 17017 2191 17051
rect 2133 17011 2191 17017
rect 18690 17008 18696 17060
rect 18748 17048 18754 17060
rect 27065 17051 27123 17057
rect 27065 17048 27077 17051
rect 18748 17020 27077 17048
rect 18748 17008 18754 17020
rect 27065 17017 27077 17020
rect 27111 17017 27123 17051
rect 27065 17011 27123 17017
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 17678 16980 17684 16992
rect 17639 16952 17684 16980
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18506 16980 18512 16992
rect 18012 16952 18512 16980
rect 18012 16940 18018 16952
rect 18506 16940 18512 16952
rect 18564 16940 18570 16992
rect 19429 16983 19487 16989
rect 19429 16949 19441 16983
rect 19475 16980 19487 16983
rect 19518 16980 19524 16992
rect 19475 16952 19524 16980
rect 19475 16949 19487 16952
rect 19429 16943 19487 16949
rect 19518 16940 19524 16952
rect 19576 16940 19582 16992
rect 22833 16983 22891 16989
rect 22833 16949 22845 16983
rect 22879 16980 22891 16983
rect 24026 16980 24032 16992
rect 22879 16952 24032 16980
rect 22879 16949 22891 16952
rect 22833 16943 22891 16949
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 25222 16940 25228 16992
rect 25280 16980 25286 16992
rect 30009 16983 30067 16989
rect 30009 16980 30021 16983
rect 25280 16952 30021 16980
rect 25280 16940 25286 16952
rect 30009 16949 30021 16952
rect 30055 16949 30067 16983
rect 30009 16943 30067 16949
rect 1104 16890 30820 16912
rect 1104 16838 5915 16890
rect 5967 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 15846 16890
rect 15898 16838 15910 16890
rect 15962 16838 15974 16890
rect 16026 16838 16038 16890
rect 16090 16838 16102 16890
rect 16154 16838 25776 16890
rect 25828 16838 25840 16890
rect 25892 16838 25904 16890
rect 25956 16838 25968 16890
rect 26020 16838 26032 16890
rect 26084 16838 30820 16890
rect 1104 16816 30820 16838
rect 17218 16776 17224 16788
rect 17179 16748 17224 16776
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 18095 16779 18153 16785
rect 18095 16745 18107 16779
rect 18141 16776 18153 16779
rect 18966 16776 18972 16788
rect 18141 16748 18972 16776
rect 18141 16745 18153 16748
rect 18095 16739 18153 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19886 16736 19892 16788
rect 19944 16776 19950 16788
rect 20349 16779 20407 16785
rect 20349 16776 20361 16779
rect 19944 16748 20361 16776
rect 19944 16736 19950 16748
rect 20349 16745 20361 16748
rect 20395 16745 20407 16779
rect 27614 16776 27620 16788
rect 27575 16748 27620 16776
rect 20349 16739 20407 16745
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 18690 16708 18696 16720
rect 6886 16680 18696 16708
rect 6886 16640 6914 16680
rect 18690 16668 18696 16680
rect 18748 16668 18754 16720
rect 18874 16668 18880 16720
rect 18932 16708 18938 16720
rect 18932 16680 19012 16708
rect 18932 16668 18938 16680
rect 2332 16612 6914 16640
rect 2332 16581 2360 16612
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 16540 16612 16804 16640
rect 16540 16600 16546 16612
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16572 1455 16575
rect 2317 16575 2375 16581
rect 1443 16544 2176 16572
rect 1443 16541 1455 16544
rect 1397 16535 1455 16541
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 2148 16445 2176 16544
rect 2317 16541 2329 16575
rect 2363 16574 2375 16575
rect 2363 16546 2397 16574
rect 16206 16572 16212 16584
rect 2363 16541 2375 16546
rect 16167 16544 16212 16572
rect 2317 16535 2375 16541
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16776 16572 16804 16612
rect 16850 16600 16856 16652
rect 16908 16640 16914 16652
rect 16908 16612 16953 16640
rect 16908 16600 16914 16612
rect 17037 16575 17095 16581
rect 17037 16572 17049 16575
rect 16776 16544 17049 16572
rect 17037 16541 17049 16544
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16572 17923 16575
rect 18598 16572 18604 16584
rect 17911 16544 18604 16572
rect 17911 16541 17923 16544
rect 17865 16535 17923 16541
rect 18598 16532 18604 16544
rect 18656 16572 18662 16584
rect 18984 16572 19012 16680
rect 19426 16668 19432 16720
rect 19484 16668 19490 16720
rect 19444 16581 19472 16668
rect 19886 16640 19892 16652
rect 19799 16612 19892 16640
rect 19886 16600 19892 16612
rect 19944 16600 19950 16652
rect 20438 16600 20444 16652
rect 20496 16640 20502 16652
rect 20717 16643 20775 16649
rect 20717 16640 20729 16643
rect 20496 16612 20729 16640
rect 20496 16600 20502 16612
rect 20717 16609 20729 16612
rect 20763 16609 20775 16643
rect 20717 16603 20775 16609
rect 26602 16600 26608 16652
rect 26660 16640 26666 16652
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 26660 16612 27077 16640
rect 26660 16600 26666 16612
rect 27065 16609 27077 16612
rect 27111 16640 27123 16643
rect 27522 16640 27528 16652
rect 27111 16612 27528 16640
rect 27111 16609 27123 16612
rect 27065 16603 27123 16609
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 28810 16600 28816 16652
rect 28868 16640 28874 16652
rect 31294 16640 31300 16652
rect 28868 16612 31300 16640
rect 28868 16600 28874 16612
rect 31294 16600 31300 16612
rect 31352 16600 31358 16652
rect 18656 16544 19012 16572
rect 19430 16575 19488 16581
rect 18656 16532 18662 16544
rect 19430 16541 19442 16575
rect 19476 16541 19488 16575
rect 19430 16535 19488 16541
rect 19702 16532 19708 16584
rect 19760 16581 19766 16584
rect 19760 16575 19789 16581
rect 19777 16541 19789 16575
rect 19916 16572 19944 16600
rect 19760 16535 19789 16541
rect 19904 16544 19944 16572
rect 19760 16532 19766 16535
rect 2682 16464 2688 16516
rect 2740 16504 2746 16516
rect 18690 16504 18696 16516
rect 2740 16476 18696 16504
rect 2740 16464 2746 16476
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 18874 16464 18880 16516
rect 18932 16504 18938 16516
rect 19521 16507 19579 16513
rect 19521 16504 19533 16507
rect 18932 16476 19533 16504
rect 18932 16464 18938 16476
rect 19521 16473 19533 16476
rect 19567 16473 19579 16507
rect 19521 16467 19579 16473
rect 19613 16507 19671 16513
rect 19613 16473 19625 16507
rect 19659 16473 19671 16507
rect 19904 16504 19932 16544
rect 20070 16532 20076 16584
rect 20128 16572 20134 16584
rect 20533 16575 20591 16581
rect 20533 16572 20545 16575
rect 20128 16544 20545 16572
rect 20128 16532 20134 16544
rect 20533 16541 20545 16544
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 20622 16532 20628 16584
rect 20680 16572 20686 16584
rect 20809 16575 20867 16581
rect 20680 16544 20725 16572
rect 20680 16532 20686 16544
rect 20809 16541 20821 16575
rect 20855 16541 20867 16575
rect 20809 16535 20867 16541
rect 20824 16504 20852 16535
rect 21174 16532 21180 16584
rect 21232 16572 21238 16584
rect 28059 16575 28117 16581
rect 28059 16572 28071 16575
rect 21232 16544 28071 16572
rect 21232 16532 21238 16544
rect 28059 16541 28071 16544
rect 28105 16541 28117 16575
rect 28059 16535 28117 16541
rect 28258 16532 28264 16584
rect 28316 16572 28322 16584
rect 28353 16575 28411 16581
rect 28353 16572 28365 16575
rect 28316 16544 28365 16572
rect 28316 16532 28322 16544
rect 28353 16541 28365 16544
rect 28399 16541 28411 16575
rect 30098 16572 30104 16584
rect 30059 16544 30104 16572
rect 28353 16535 28411 16541
rect 30098 16532 30104 16544
rect 30156 16532 30162 16584
rect 19904 16476 20852 16504
rect 19613 16467 19671 16473
rect 2133 16439 2191 16445
rect 2133 16405 2145 16439
rect 2179 16405 2191 16439
rect 2133 16399 2191 16405
rect 16393 16439 16451 16445
rect 16393 16405 16405 16439
rect 16439 16436 16451 16439
rect 16850 16436 16856 16448
rect 16439 16408 16856 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 16850 16396 16856 16408
rect 16908 16396 16914 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19625 16436 19653 16467
rect 25038 16464 25044 16516
rect 25096 16504 25102 16516
rect 25498 16504 25504 16516
rect 25096 16476 25504 16504
rect 25096 16464 25102 16476
rect 25498 16464 25504 16476
rect 25556 16464 25562 16516
rect 27249 16507 27307 16513
rect 27249 16473 27261 16507
rect 27295 16504 27307 16507
rect 27706 16504 27712 16516
rect 27295 16476 27712 16504
rect 27295 16473 27307 16476
rect 27249 16467 27307 16473
rect 27706 16464 27712 16476
rect 27764 16504 27770 16516
rect 28629 16507 28687 16513
rect 28629 16504 28641 16507
rect 27764 16476 28641 16504
rect 27764 16464 27770 16476
rect 28629 16473 28641 16476
rect 28675 16504 28687 16507
rect 28718 16504 28724 16516
rect 28675 16476 28724 16504
rect 28675 16473 28687 16476
rect 28629 16467 28687 16473
rect 28718 16464 28724 16476
rect 28776 16464 28782 16516
rect 19392 16408 19653 16436
rect 19392 16396 19398 16408
rect 19886 16396 19892 16448
rect 19944 16436 19950 16448
rect 26679 16439 26737 16445
rect 26679 16436 26691 16439
rect 19944 16408 26691 16436
rect 19944 16396 19950 16408
rect 26679 16405 26691 16408
rect 26725 16405 26737 16439
rect 26679 16399 26737 16405
rect 27157 16439 27215 16445
rect 27157 16405 27169 16439
rect 27203 16436 27215 16439
rect 27338 16436 27344 16448
rect 27203 16408 27344 16436
rect 27203 16405 27215 16408
rect 27157 16399 27215 16405
rect 27338 16396 27344 16408
rect 27396 16396 27402 16448
rect 27614 16396 27620 16448
rect 27672 16436 27678 16448
rect 28537 16439 28595 16445
rect 28537 16436 28549 16439
rect 27672 16408 28549 16436
rect 27672 16396 27678 16408
rect 28537 16405 28549 16408
rect 28583 16405 28595 16439
rect 28537 16399 28595 16405
rect 29822 16396 29828 16448
rect 29880 16436 29886 16448
rect 29917 16439 29975 16445
rect 29917 16436 29929 16439
rect 29880 16408 29929 16436
rect 29880 16396 29886 16408
rect 29917 16405 29929 16408
rect 29963 16405 29975 16439
rect 29917 16399 29975 16405
rect 1104 16346 30820 16368
rect 1104 16294 10880 16346
rect 10932 16294 10944 16346
rect 10996 16294 11008 16346
rect 11060 16294 11072 16346
rect 11124 16294 11136 16346
rect 11188 16294 20811 16346
rect 20863 16294 20875 16346
rect 20927 16294 20939 16346
rect 20991 16294 21003 16346
rect 21055 16294 21067 16346
rect 21119 16294 30820 16346
rect 1104 16272 30820 16294
rect 18230 16232 18236 16244
rect 1872 16204 18236 16232
rect 1872 16105 1900 16204
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 28151 16235 28209 16241
rect 28151 16232 28163 16235
rect 18472 16204 28163 16232
rect 18472 16192 18478 16204
rect 28151 16201 28163 16204
rect 28197 16201 28209 16235
rect 28151 16195 28209 16201
rect 28350 16192 28356 16244
rect 28408 16232 28414 16244
rect 31110 16232 31116 16244
rect 28408 16204 31116 16232
rect 28408 16192 28414 16204
rect 31110 16192 31116 16204
rect 31168 16192 31174 16244
rect 16942 16164 16948 16176
rect 6886 16136 16948 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 2501 16099 2559 16105
rect 2501 16065 2513 16099
rect 2547 16096 2559 16099
rect 6886 16096 6914 16136
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 17120 16167 17178 16173
rect 17120 16133 17132 16167
rect 17166 16164 17178 16167
rect 17678 16164 17684 16176
rect 17166 16136 17684 16164
rect 17166 16133 17178 16136
rect 17120 16127 17178 16133
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 17770 16124 17776 16176
rect 17828 16164 17834 16176
rect 17908 16164 17914 16176
rect 17828 16136 17914 16164
rect 17828 16124 17834 16136
rect 17908 16124 17914 16136
rect 17966 16124 17972 16176
rect 25317 16167 25375 16173
rect 25317 16133 25329 16167
rect 25363 16164 25375 16167
rect 26234 16164 26240 16176
rect 25363 16136 26240 16164
rect 25363 16133 25375 16136
rect 25317 16127 25375 16133
rect 26234 16124 26240 16136
rect 26292 16124 26298 16176
rect 27062 16124 27068 16176
rect 27120 16164 27126 16176
rect 27338 16164 27344 16176
rect 27120 16136 27344 16164
rect 27120 16124 27126 16136
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 27614 16124 27620 16176
rect 27672 16164 27678 16176
rect 27709 16167 27767 16173
rect 27709 16164 27721 16167
rect 27672 16136 27721 16164
rect 27672 16124 27678 16136
rect 27709 16133 27721 16136
rect 27755 16164 27767 16167
rect 28629 16167 28687 16173
rect 28629 16164 28641 16167
rect 27755 16136 28641 16164
rect 27755 16133 27767 16136
rect 27709 16127 27767 16133
rect 28629 16133 28641 16136
rect 28675 16133 28687 16167
rect 28629 16127 28687 16133
rect 28718 16124 28724 16176
rect 28776 16164 28782 16176
rect 28776 16136 28821 16164
rect 28776 16124 28782 16136
rect 16850 16096 16856 16108
rect 2547 16068 6914 16096
rect 16811 16068 16856 16096
rect 2547 16065 2559 16068
rect 2501 16059 2559 16065
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 19334 16096 19340 16108
rect 18739 16068 19340 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 19444 16068 20545 16096
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 19444 16028 19472 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 21818 16096 21824 16108
rect 21779 16068 21824 16096
rect 20533 16059 20591 16065
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 25038 16096 25044 16108
rect 24999 16068 25044 16096
rect 25038 16056 25044 16068
rect 25096 16056 25102 16108
rect 25222 16096 25228 16108
rect 25183 16068 25228 16096
rect 25222 16056 25228 16068
rect 25280 16056 25286 16108
rect 25409 16099 25467 16105
rect 25409 16065 25421 16099
rect 25455 16096 25467 16099
rect 25590 16096 25596 16108
rect 25455 16068 25596 16096
rect 25455 16065 25467 16068
rect 25409 16059 25467 16065
rect 25590 16056 25596 16068
rect 25648 16056 25654 16108
rect 28442 16096 28448 16108
rect 28403 16068 28448 16096
rect 28442 16056 28448 16068
rect 28500 16056 28506 16108
rect 29914 16096 29920 16108
rect 29875 16068 29920 16096
rect 29914 16056 29920 16068
rect 29972 16056 29978 16108
rect 18380 16000 19472 16028
rect 20257 16031 20315 16037
rect 18380 15988 18386 16000
rect 20257 15997 20269 16031
rect 20303 16028 20315 16031
rect 20346 16028 20352 16040
rect 20303 16000 20352 16028
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 27430 15988 27436 16040
rect 27488 16028 27494 16040
rect 30101 16031 30159 16037
rect 30101 16028 30113 16031
rect 27488 16000 30113 16028
rect 27488 15988 27494 16000
rect 30101 15997 30113 16000
rect 30147 15997 30159 16031
rect 30101 15991 30159 15997
rect 18233 15963 18291 15969
rect 18233 15929 18245 15963
rect 18279 15960 18291 15963
rect 18598 15960 18604 15972
rect 18279 15932 18604 15960
rect 18279 15929 18291 15932
rect 18233 15923 18291 15929
rect 18598 15920 18604 15932
rect 18656 15920 18662 15972
rect 21910 15920 21916 15972
rect 21968 15960 21974 15972
rect 22005 15963 22063 15969
rect 22005 15960 22017 15963
rect 21968 15932 22017 15960
rect 21968 15920 21974 15932
rect 22005 15929 22017 15932
rect 22051 15929 22063 15963
rect 22005 15923 22063 15929
rect 25593 15963 25651 15969
rect 25593 15929 25605 15963
rect 25639 15960 25651 15963
rect 26142 15960 26148 15972
rect 25639 15932 26148 15960
rect 25639 15929 25651 15932
rect 25593 15923 25651 15929
rect 26142 15920 26148 15932
rect 26200 15920 26206 15972
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1673 15895 1731 15901
rect 1673 15892 1685 15895
rect 1452 15864 1685 15892
rect 1452 15852 1458 15864
rect 1673 15861 1685 15864
rect 1719 15861 1731 15895
rect 1673 15855 1731 15861
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 2317 15895 2375 15901
rect 2317 15892 2329 15895
rect 1820 15864 2329 15892
rect 1820 15852 1826 15864
rect 2317 15861 2329 15864
rect 2363 15861 2375 15895
rect 2317 15855 2375 15861
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 18046 15892 18052 15904
rect 16724 15864 18052 15892
rect 16724 15852 16730 15864
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 19337 15895 19395 15901
rect 19337 15861 19349 15895
rect 19383 15892 19395 15895
rect 19702 15892 19708 15904
rect 19383 15864 19708 15892
rect 19383 15861 19395 15864
rect 19337 15855 19395 15861
rect 19702 15852 19708 15864
rect 19760 15852 19766 15904
rect 27982 15852 27988 15904
rect 28040 15892 28046 15904
rect 28442 15892 28448 15904
rect 28040 15864 28448 15892
rect 28040 15852 28046 15864
rect 28442 15852 28448 15864
rect 28500 15852 28506 15904
rect 1104 15802 30820 15824
rect 1104 15750 5915 15802
rect 5967 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 15846 15802
rect 15898 15750 15910 15802
rect 15962 15750 15974 15802
rect 16026 15750 16038 15802
rect 16090 15750 16102 15802
rect 16154 15750 25776 15802
rect 25828 15750 25840 15802
rect 25892 15750 25904 15802
rect 25956 15750 25968 15802
rect 26020 15750 26032 15802
rect 26084 15750 30820 15802
rect 1104 15728 30820 15750
rect 16666 15688 16672 15700
rect 6886 15660 16672 15688
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 1762 15484 1768 15496
rect 1443 15456 1768 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 1762 15444 1768 15456
rect 1820 15444 1826 15496
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 6886 15484 6914 15660
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 16942 15648 16948 15700
rect 17000 15688 17006 15700
rect 27157 15691 27215 15697
rect 27157 15688 27169 15691
rect 17000 15660 27169 15688
rect 17000 15648 17006 15660
rect 27157 15657 27169 15660
rect 27203 15657 27215 15691
rect 27157 15651 27215 15657
rect 28258 15648 28264 15700
rect 28316 15688 28322 15700
rect 28813 15691 28871 15697
rect 28813 15688 28825 15691
rect 28316 15660 28825 15688
rect 28316 15648 28322 15660
rect 28813 15657 28825 15660
rect 28859 15657 28871 15691
rect 28813 15651 28871 15657
rect 16853 15623 16911 15629
rect 16853 15589 16865 15623
rect 16899 15620 16911 15623
rect 18693 15623 18751 15629
rect 16899 15592 17356 15620
rect 16899 15589 16911 15592
rect 16853 15583 16911 15589
rect 17328 15561 17356 15592
rect 18693 15589 18705 15623
rect 18739 15620 18751 15623
rect 19334 15620 19340 15632
rect 18739 15592 19340 15620
rect 18739 15589 18751 15592
rect 18693 15583 18751 15589
rect 19334 15580 19340 15592
rect 19392 15580 19398 15632
rect 20346 15580 20352 15632
rect 20404 15620 20410 15632
rect 20625 15623 20683 15629
rect 20625 15620 20637 15623
rect 20404 15592 20637 15620
rect 20404 15580 20410 15592
rect 20625 15589 20637 15592
rect 20671 15589 20683 15623
rect 20625 15583 20683 15589
rect 25777 15623 25835 15629
rect 25777 15589 25789 15623
rect 25823 15620 25835 15623
rect 28994 15620 29000 15632
rect 25823 15592 29000 15620
rect 25823 15589 25835 15592
rect 25777 15583 25835 15589
rect 28994 15580 29000 15592
rect 29052 15580 29058 15632
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 20530 15552 20536 15564
rect 17313 15515 17371 15521
rect 20180 15524 20536 15552
rect 20180 15496 20208 15524
rect 20530 15512 20536 15524
rect 20588 15512 20594 15564
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15552 21327 15555
rect 21634 15552 21640 15564
rect 21315 15524 21640 15552
rect 21315 15521 21327 15524
rect 21269 15515 21327 15521
rect 21634 15512 21640 15524
rect 21692 15552 21698 15564
rect 21910 15552 21916 15564
rect 21692 15524 21916 15552
rect 21692 15512 21698 15524
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 26878 15552 26884 15564
rect 26660 15524 26884 15552
rect 26660 15512 26666 15524
rect 26878 15512 26884 15524
rect 26936 15512 26942 15564
rect 27706 15552 27712 15564
rect 27667 15524 27712 15552
rect 27706 15512 27712 15524
rect 27764 15512 27770 15564
rect 2363 15456 6914 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 16669 15487 16727 15493
rect 16669 15484 16681 15487
rect 16632 15456 16681 15484
rect 16632 15444 16638 15456
rect 16669 15453 16681 15456
rect 16715 15453 16727 15487
rect 16669 15447 16727 15453
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 19300 15456 19349 15484
rect 19300 15444 19306 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 19702 15484 19708 15496
rect 19663 15456 19708 15484
rect 19337 15447 19395 15453
rect 17580 15419 17638 15425
rect 17580 15385 17592 15419
rect 17626 15416 17638 15419
rect 18414 15416 18420 15428
rect 17626 15388 18420 15416
rect 17626 15385 17638 15388
rect 17580 15379 17638 15385
rect 18414 15376 18420 15388
rect 18472 15376 18478 15428
rect 19352 15416 19380 15447
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 20162 15484 20168 15496
rect 20123 15456 20168 15484
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 20438 15484 20444 15496
rect 20399 15456 20444 15484
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 21542 15484 21548 15496
rect 21503 15456 21548 15484
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 24486 15444 24492 15496
rect 24544 15484 24550 15496
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 24544 15456 25237 15484
rect 24544 15444 24550 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25590 15484 25596 15496
rect 25503 15456 25596 15484
rect 25225 15447 25283 15453
rect 25590 15444 25596 15456
rect 25648 15484 25654 15496
rect 26142 15484 26148 15496
rect 25648 15456 26148 15484
rect 25648 15444 25654 15456
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 26234 15444 26240 15496
rect 26292 15484 26298 15496
rect 27430 15484 27436 15496
rect 26292 15456 27436 15484
rect 26292 15444 26298 15456
rect 27430 15444 27436 15456
rect 27488 15444 27494 15496
rect 28994 15484 29000 15496
rect 28955 15456 29000 15484
rect 28994 15444 29000 15456
rect 29052 15444 29058 15496
rect 20622 15416 20628 15428
rect 19352 15388 20628 15416
rect 20622 15376 20628 15388
rect 20680 15376 20686 15428
rect 24210 15376 24216 15428
rect 24268 15416 24274 15428
rect 24670 15416 24676 15428
rect 24268 15388 24676 15416
rect 24268 15376 24274 15388
rect 24670 15376 24676 15388
rect 24728 15376 24734 15428
rect 25406 15416 25412 15428
rect 25367 15388 25412 15416
rect 25406 15376 25412 15388
rect 25464 15376 25470 15428
rect 25501 15419 25559 15425
rect 25501 15385 25513 15419
rect 25547 15416 25559 15419
rect 26878 15416 26884 15428
rect 25547 15388 26884 15416
rect 25547 15385 25559 15388
rect 25501 15379 25559 15385
rect 26878 15376 26884 15388
rect 26936 15376 26942 15428
rect 27614 15416 27620 15428
rect 27575 15388 27620 15416
rect 27614 15376 27620 15388
rect 27672 15376 27678 15428
rect 29914 15416 29920 15428
rect 29875 15388 29920 15416
rect 29914 15376 29920 15388
rect 29972 15376 29978 15428
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2130 15348 2136 15360
rect 2091 15320 2136 15348
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 27522 15308 27528 15360
rect 27580 15348 27586 15360
rect 30009 15351 30067 15357
rect 30009 15348 30021 15351
rect 27580 15320 30021 15348
rect 27580 15308 27586 15320
rect 30009 15317 30021 15320
rect 30055 15317 30067 15351
rect 30009 15311 30067 15317
rect 1104 15258 30820 15280
rect 1104 15206 10880 15258
rect 10932 15206 10944 15258
rect 10996 15206 11008 15258
rect 11060 15206 11072 15258
rect 11124 15206 11136 15258
rect 11188 15206 20811 15258
rect 20863 15206 20875 15258
rect 20927 15206 20939 15258
rect 20991 15206 21003 15258
rect 21055 15206 21067 15258
rect 21119 15206 30820 15258
rect 1104 15184 30820 15206
rect 22462 15144 22468 15156
rect 21836 15116 22468 15144
rect 19794 15036 19800 15088
rect 19852 15076 19858 15088
rect 20346 15076 20352 15088
rect 19852 15048 20352 15076
rect 19852 15036 19858 15048
rect 20346 15036 20352 15048
rect 20404 15076 20410 15088
rect 20404 15048 21128 15076
rect 20404 15036 20410 15048
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 19334 15008 19340 15020
rect 19295 14980 19340 15008
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 20772 14980 20821 15008
rect 20772 14968 20778 14980
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 21100 15017 21128 15048
rect 21085 15011 21143 15017
rect 20956 14980 21001 15008
rect 20956 14968 20962 14980
rect 21085 14977 21097 15011
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 21232 14980 21277 15008
rect 21232 14968 21238 14980
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19484 14912 19625 14940
rect 19484 14900 19490 14912
rect 19613 14909 19625 14912
rect 19659 14940 19671 14943
rect 20070 14940 20076 14952
rect 19659 14912 20076 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 21542 14900 21548 14952
rect 21600 14940 21606 14952
rect 21836 14949 21864 15116
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 23201 15147 23259 15153
rect 23201 15113 23213 15147
rect 23247 15144 23259 15147
rect 23474 15144 23480 15156
rect 23247 15116 23480 15144
rect 23247 15113 23259 15116
rect 23201 15107 23259 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 23753 15147 23811 15153
rect 23753 15113 23765 15147
rect 23799 15113 23811 15147
rect 23753 15107 23811 15113
rect 24673 15147 24731 15153
rect 24673 15113 24685 15147
rect 24719 15144 24731 15147
rect 25406 15144 25412 15156
rect 24719 15116 25412 15144
rect 24719 15113 24731 15116
rect 24673 15107 24731 15113
rect 23768 15076 23796 15107
rect 25406 15104 25412 15116
rect 25464 15104 25470 15156
rect 26237 15147 26295 15153
rect 26237 15113 26249 15147
rect 26283 15144 26295 15147
rect 26283 15116 26372 15144
rect 26283 15113 26295 15116
rect 26237 15107 26295 15113
rect 25222 15076 25228 15088
rect 23768 15048 25228 15076
rect 25222 15036 25228 15048
rect 25280 15036 25286 15088
rect 22088 15011 22146 15017
rect 22088 14977 22100 15011
rect 22134 15008 22146 15011
rect 22462 15008 22468 15020
rect 22134 14980 22468 15008
rect 22134 14977 22146 14980
rect 22088 14971 22146 14977
rect 22462 14968 22468 14980
rect 22520 14968 22526 15020
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 23808 14980 23949 15008
rect 23808 14968 23814 14980
rect 23937 14977 23949 14980
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 24026 14968 24032 15020
rect 24084 15008 24090 15020
rect 24857 15011 24915 15017
rect 24084 14980 24348 15008
rect 24084 14968 24090 14980
rect 21821 14943 21879 14949
rect 21821 14940 21833 14943
rect 21600 14912 21833 14940
rect 21600 14900 21606 14912
rect 21821 14909 21833 14912
rect 21867 14909 21879 14943
rect 21821 14903 21879 14909
rect 23198 14900 23204 14952
rect 23256 14940 23262 14952
rect 24213 14943 24271 14949
rect 24213 14940 24225 14943
rect 23256 14912 24225 14940
rect 23256 14900 23262 14912
rect 24213 14909 24225 14912
rect 24259 14909 24271 14943
rect 24320 14940 24348 14980
rect 24857 14977 24869 15011
rect 24903 15008 24915 15011
rect 25406 15008 25412 15020
rect 24903 14980 25412 15008
rect 24903 14977 24915 14980
rect 24857 14971 24915 14977
rect 25406 14968 25412 14980
rect 25464 14968 25470 15020
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24320 14912 25145 14940
rect 24213 14903 24271 14909
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 26344 14940 26372 15116
rect 27430 15104 27436 15156
rect 27488 15144 27494 15156
rect 28258 15144 28264 15156
rect 27488 15116 27752 15144
rect 28219 15116 28264 15144
rect 27488 15104 27494 15116
rect 27614 15076 27620 15088
rect 26436 15048 27620 15076
rect 26436 15017 26464 15048
rect 27614 15036 27620 15048
rect 27672 15036 27678 15088
rect 27724 15076 27752 15116
rect 28258 15104 28264 15116
rect 28316 15104 28322 15156
rect 27724 15048 29592 15076
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 27062 14968 27068 15020
rect 27120 15008 27126 15020
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 27120 14980 27169 15008
rect 27120 14968 27126 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 27982 15008 27988 15020
rect 27157 14971 27215 14977
rect 27448 14980 27988 15008
rect 27448 14940 27476 14980
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 28074 14968 28080 15020
rect 28132 15008 28138 15020
rect 29564 15017 29592 15048
rect 28169 15011 28227 15017
rect 28169 15008 28181 15011
rect 28132 14980 28181 15008
rect 28132 14968 28138 14980
rect 28169 14977 28181 14980
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 29549 15011 29607 15017
rect 29549 14977 29561 15011
rect 29595 14977 29607 15011
rect 29549 14971 29607 14977
rect 26344 14912 27476 14940
rect 25133 14903 25191 14909
rect 27522 14900 27528 14952
rect 27580 14940 27586 14952
rect 28353 14943 28411 14949
rect 28353 14940 28365 14943
rect 27580 14912 28365 14940
rect 27580 14900 27586 14912
rect 28353 14909 28365 14912
rect 28399 14909 28411 14943
rect 28353 14903 28411 14909
rect 28902 14900 28908 14952
rect 28960 14940 28966 14952
rect 29273 14943 29331 14949
rect 29273 14940 29285 14943
rect 28960 14912 29285 14940
rect 28960 14900 28966 14912
rect 29273 14909 29285 14912
rect 29319 14909 29331 14943
rect 29273 14903 29331 14909
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 27341 14875 27399 14881
rect 27341 14872 27353 14875
rect 17276 14844 20760 14872
rect 17276 14832 17282 14844
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 20036 14776 20637 14804
rect 20036 14764 20042 14776
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 20732 14804 20760 14844
rect 23124 14844 27353 14872
rect 23124 14804 23152 14844
rect 27341 14841 27353 14844
rect 27387 14841 27399 14875
rect 27341 14835 27399 14841
rect 20732 14776 23152 14804
rect 20625 14767 20683 14773
rect 23382 14764 23388 14816
rect 23440 14804 23446 14816
rect 24026 14804 24032 14816
rect 23440 14776 24032 14804
rect 23440 14764 23446 14776
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 24121 14807 24179 14813
rect 24121 14773 24133 14807
rect 24167 14804 24179 14807
rect 25038 14804 25044 14816
rect 24167 14776 25044 14804
rect 24167 14773 24179 14776
rect 24121 14767 24179 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 25406 14764 25412 14816
rect 25464 14804 25470 14816
rect 26326 14804 26332 14816
rect 25464 14776 26332 14804
rect 25464 14764 25470 14776
rect 26326 14764 26332 14776
rect 26384 14764 26390 14816
rect 27430 14764 27436 14816
rect 27488 14804 27494 14816
rect 27801 14807 27859 14813
rect 27801 14804 27813 14807
rect 27488 14776 27813 14804
rect 27488 14764 27494 14776
rect 27801 14773 27813 14776
rect 27847 14773 27859 14807
rect 27801 14767 27859 14773
rect 1104 14714 30820 14736
rect 1104 14662 5915 14714
rect 5967 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 15846 14714
rect 15898 14662 15910 14714
rect 15962 14662 15974 14714
rect 16026 14662 16038 14714
rect 16090 14662 16102 14714
rect 16154 14662 25776 14714
rect 25828 14662 25840 14714
rect 25892 14662 25904 14714
rect 25956 14662 25968 14714
rect 26020 14662 26032 14714
rect 26084 14662 30820 14714
rect 1104 14640 30820 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 17218 14600 17224 14612
rect 1452 14572 17224 14600
rect 1452 14560 1458 14572
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 18414 14560 18420 14612
rect 18472 14600 18478 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 18472 14572 19257 14600
rect 18472 14560 18478 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 19245 14563 19303 14569
rect 20070 14560 20076 14612
rect 20128 14600 20134 14612
rect 20349 14603 20407 14609
rect 20349 14600 20361 14603
rect 20128 14572 20361 14600
rect 20128 14560 20134 14572
rect 20349 14569 20361 14572
rect 20395 14569 20407 14603
rect 20349 14563 20407 14569
rect 20809 14603 20867 14609
rect 20809 14569 20821 14603
rect 20855 14600 20867 14603
rect 21818 14600 21824 14612
rect 20855 14572 21824 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 21818 14560 21824 14572
rect 21876 14560 21882 14612
rect 22462 14600 22468 14612
rect 22423 14572 22468 14600
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 25406 14600 25412 14612
rect 24912 14572 25412 14600
rect 24912 14560 24918 14572
rect 25406 14560 25412 14572
rect 25464 14560 25470 14612
rect 26329 14603 26387 14609
rect 26329 14569 26341 14603
rect 26375 14569 26387 14603
rect 30834 14600 30840 14612
rect 26329 14563 26387 14569
rect 27264 14572 30840 14600
rect 6270 14492 6276 14544
rect 6328 14532 6334 14544
rect 19518 14532 19524 14544
rect 6328 14504 19524 14532
rect 6328 14492 6334 14504
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 20254 14464 20260 14476
rect 19720 14436 20260 14464
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2130 14396 2136 14408
rect 1443 14368 2136 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 19426 14356 19432 14408
rect 19484 14405 19490 14408
rect 19484 14399 19533 14405
rect 19484 14365 19487 14399
rect 19521 14365 19533 14399
rect 19610 14396 19616 14408
rect 19571 14368 19616 14396
rect 19484 14359 19533 14365
rect 19484 14356 19490 14359
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 19720 14405 19748 14436
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14433 20499 14467
rect 20441 14427 20499 14433
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 19978 14396 19984 14408
rect 19935 14368 19984 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20162 14396 20168 14408
rect 20075 14368 20168 14396
rect 20162 14356 20168 14368
rect 20220 14396 20226 14408
rect 20456 14396 20484 14427
rect 20898 14424 20904 14476
rect 20956 14464 20962 14476
rect 22925 14467 22983 14473
rect 22925 14464 22937 14467
rect 20956 14436 22937 14464
rect 20956 14424 20962 14436
rect 22925 14433 22937 14436
rect 22971 14464 22983 14467
rect 23474 14464 23480 14476
rect 22971 14436 23480 14464
rect 22971 14433 22983 14436
rect 22925 14427 22983 14433
rect 23474 14424 23480 14436
rect 23532 14424 23538 14476
rect 20622 14396 20628 14408
rect 20220 14368 20484 14396
rect 20583 14368 20628 14396
rect 20220 14356 20226 14368
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14396 22891 14399
rect 23106 14396 23112 14408
rect 22879 14368 23112 14396
rect 22879 14365 22891 14368
rect 22833 14359 22891 14365
rect 1578 14260 1584 14272
rect 1539 14232 1584 14260
rect 1578 14220 1584 14232
rect 1636 14220 1642 14272
rect 19518 14220 19524 14272
rect 19576 14260 19582 14272
rect 20180 14260 20208 14356
rect 20349 14331 20407 14337
rect 20349 14297 20361 14331
rect 20395 14328 20407 14331
rect 20438 14328 20444 14340
rect 20395 14300 20444 14328
rect 20395 14297 20407 14300
rect 20349 14291 20407 14297
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 22664 14328 22692 14359
rect 23106 14356 23112 14368
rect 23164 14356 23170 14408
rect 25314 14356 25320 14408
rect 25372 14396 25378 14408
rect 25777 14399 25835 14405
rect 25777 14396 25789 14399
rect 25372 14368 25789 14396
rect 25372 14356 25378 14368
rect 25777 14365 25789 14368
rect 25823 14365 25835 14399
rect 26142 14396 26148 14408
rect 26103 14368 26148 14396
rect 25777 14359 25835 14365
rect 26142 14356 26148 14368
rect 26200 14356 26206 14408
rect 26344 14396 26372 14563
rect 27062 14492 27068 14544
rect 27120 14532 27126 14544
rect 27120 14504 27165 14532
rect 27120 14492 27126 14504
rect 27264 14396 27292 14572
rect 30834 14560 30840 14572
rect 30892 14560 30898 14612
rect 27338 14492 27344 14544
rect 27396 14532 27402 14544
rect 27396 14504 27752 14532
rect 27396 14492 27402 14504
rect 27522 14424 27528 14476
rect 27580 14464 27586 14476
rect 27617 14467 27675 14473
rect 27617 14464 27629 14467
rect 27580 14436 27629 14464
rect 27580 14424 27586 14436
rect 27617 14433 27629 14436
rect 27663 14433 27675 14467
rect 27724 14464 27752 14504
rect 27982 14492 27988 14544
rect 28040 14532 28046 14544
rect 28353 14535 28411 14541
rect 28353 14532 28365 14535
rect 28040 14504 28365 14532
rect 28040 14492 28046 14504
rect 28353 14501 28365 14504
rect 28399 14501 28411 14535
rect 30009 14535 30067 14541
rect 30009 14532 30021 14535
rect 28353 14495 28411 14501
rect 28460 14504 30021 14532
rect 28258 14464 28264 14476
rect 27724 14436 28264 14464
rect 27617 14427 27675 14433
rect 28258 14424 28264 14436
rect 28316 14464 28322 14476
rect 28460 14464 28488 14504
rect 30009 14501 30021 14504
rect 30055 14501 30067 14535
rect 30009 14495 30067 14501
rect 28316 14436 28488 14464
rect 28813 14467 28871 14473
rect 28316 14424 28322 14436
rect 28813 14433 28825 14467
rect 28859 14464 28871 14467
rect 30098 14464 30104 14476
rect 28859 14436 30104 14464
rect 28859 14433 28871 14436
rect 28813 14427 28871 14433
rect 30098 14424 30104 14436
rect 30156 14424 30162 14476
rect 26344 14368 27292 14396
rect 27433 14399 27491 14405
rect 27433 14365 27445 14399
rect 27479 14396 27491 14399
rect 27798 14396 27804 14408
rect 27479 14368 27804 14396
rect 27479 14365 27491 14368
rect 27433 14359 27491 14365
rect 27798 14356 27804 14368
rect 27856 14356 27862 14408
rect 29822 14396 29828 14408
rect 29783 14368 29828 14396
rect 29822 14356 29828 14368
rect 29880 14356 29886 14408
rect 24394 14328 24400 14340
rect 22664 14300 24400 14328
rect 24394 14288 24400 14300
rect 24452 14288 24458 14340
rect 24854 14288 24860 14340
rect 24912 14328 24918 14340
rect 25961 14331 26019 14337
rect 25961 14328 25973 14331
rect 24912 14300 25973 14328
rect 24912 14288 24918 14300
rect 25961 14297 25973 14300
rect 26007 14297 26019 14331
rect 25961 14291 26019 14297
rect 26053 14331 26111 14337
rect 26053 14297 26065 14331
rect 26099 14297 26111 14331
rect 26053 14291 26111 14297
rect 19576 14232 20208 14260
rect 19576 14220 19582 14232
rect 25774 14220 25780 14272
rect 25832 14260 25838 14272
rect 26068 14260 26096 14291
rect 28718 14288 28724 14340
rect 28776 14328 28782 14340
rect 28905 14331 28963 14337
rect 28905 14328 28917 14331
rect 28776 14300 28917 14328
rect 28776 14288 28782 14300
rect 28905 14297 28917 14300
rect 28951 14297 28963 14331
rect 28905 14291 28963 14297
rect 25832 14232 26096 14260
rect 25832 14220 25838 14232
rect 26786 14220 26792 14272
rect 26844 14260 26850 14272
rect 27525 14263 27583 14269
rect 27525 14260 27537 14263
rect 26844 14232 27537 14260
rect 26844 14220 26850 14232
rect 27525 14229 27537 14232
rect 27571 14229 27583 14263
rect 28810 14260 28816 14272
rect 28771 14232 28816 14260
rect 27525 14223 27583 14229
rect 28810 14220 28816 14232
rect 28868 14220 28874 14272
rect 1104 14170 30820 14192
rect 1104 14118 10880 14170
rect 10932 14118 10944 14170
rect 10996 14118 11008 14170
rect 11060 14118 11072 14170
rect 11124 14118 11136 14170
rect 11188 14118 20811 14170
rect 20863 14118 20875 14170
rect 20927 14118 20939 14170
rect 20991 14118 21003 14170
rect 21055 14118 21067 14170
rect 21119 14118 30820 14170
rect 1104 14096 30820 14118
rect 20530 14016 20536 14068
rect 20588 14056 20594 14068
rect 27525 14059 27583 14065
rect 27525 14056 27537 14059
rect 20588 14028 27537 14056
rect 20588 14016 20594 14028
rect 27525 14025 27537 14028
rect 27571 14025 27583 14059
rect 27525 14019 27583 14025
rect 28074 14016 28080 14068
rect 28132 14056 28138 14068
rect 28132 14028 29592 14056
rect 28132 14016 28138 14028
rect 21818 13988 21824 14000
rect 21779 13960 21824 13988
rect 21818 13948 21824 13960
rect 21876 13948 21882 14000
rect 26234 13988 26240 14000
rect 24412 13960 26240 13988
rect 1394 13920 1400 13932
rect 1355 13892 1400 13920
rect 1394 13880 1400 13892
rect 1452 13880 1458 13932
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13920 22063 13923
rect 23382 13920 23388 13932
rect 22051 13892 23388 13920
rect 22051 13889 22063 13892
rect 22005 13883 22063 13889
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 23952 13852 23980 13883
rect 24118 13880 24124 13932
rect 24176 13920 24182 13932
rect 24412 13929 24440 13960
rect 26234 13948 26240 13960
rect 26292 13948 26298 14000
rect 27430 13988 27436 14000
rect 27391 13960 27436 13988
rect 27430 13948 27436 13960
rect 27488 13948 27494 14000
rect 28445 13991 28503 13997
rect 28445 13957 28457 13991
rect 28491 13988 28503 13991
rect 28534 13988 28540 14000
rect 28491 13960 28540 13988
rect 28491 13957 28503 13960
rect 28445 13951 28503 13957
rect 28534 13948 28540 13960
rect 28592 13948 28598 14000
rect 28626 13948 28632 14000
rect 28684 13988 28690 14000
rect 28684 13960 28729 13988
rect 28684 13948 28690 13960
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 24176 13892 24225 13920
rect 24176 13880 24182 13892
rect 24213 13889 24225 13892
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 25222 13880 25228 13932
rect 25280 13920 25286 13932
rect 25498 13920 25504 13932
rect 25280 13892 25504 13920
rect 25280 13880 25286 13892
rect 25498 13880 25504 13892
rect 25556 13920 25562 13932
rect 29564 13929 29592 14028
rect 25593 13923 25651 13929
rect 25593 13920 25605 13923
rect 25556 13892 25605 13920
rect 25556 13880 25562 13892
rect 25593 13889 25605 13892
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 29549 13923 29607 13929
rect 29549 13889 29561 13923
rect 29595 13889 29607 13923
rect 29549 13883 29607 13889
rect 24578 13852 24584 13864
rect 23952 13824 24584 13852
rect 24578 13812 24584 13824
rect 24636 13812 24642 13864
rect 25869 13855 25927 13861
rect 25869 13821 25881 13855
rect 25915 13852 25927 13855
rect 26142 13852 26148 13864
rect 25915 13824 26148 13852
rect 25915 13821 25927 13824
rect 25869 13815 25927 13821
rect 26142 13812 26148 13824
rect 26200 13812 26206 13864
rect 28718 13852 28724 13864
rect 28679 13824 28724 13852
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 28902 13812 28908 13864
rect 28960 13852 28966 13864
rect 29273 13855 29331 13861
rect 29273 13852 29285 13855
rect 28960 13824 29285 13852
rect 28960 13812 28966 13824
rect 29273 13821 29285 13824
rect 29319 13821 29331 13855
rect 29273 13815 29331 13821
rect 22370 13744 22376 13796
rect 22428 13784 22434 13796
rect 22428 13756 23888 13784
rect 22428 13744 22434 13756
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 22186 13716 22192 13728
rect 22147 13688 22192 13716
rect 22186 13676 22192 13688
rect 22244 13676 22250 13728
rect 23750 13716 23756 13728
rect 23711 13688 23756 13716
rect 23750 13676 23756 13688
rect 23808 13676 23814 13728
rect 23860 13716 23888 13756
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 27706 13784 27712 13796
rect 26292 13756 27712 13784
rect 26292 13744 26298 13756
rect 27706 13744 27712 13756
rect 27764 13744 27770 13796
rect 28169 13719 28227 13725
rect 28169 13716 28181 13719
rect 23860 13688 28181 13716
rect 28169 13685 28181 13688
rect 28215 13685 28227 13719
rect 28169 13679 28227 13685
rect 1104 13626 30820 13648
rect 1104 13574 5915 13626
rect 5967 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 15846 13626
rect 15898 13574 15910 13626
rect 15962 13574 15974 13626
rect 16026 13574 16038 13626
rect 16090 13574 16102 13626
rect 16154 13574 25776 13626
rect 25828 13574 25840 13626
rect 25892 13574 25904 13626
rect 25956 13574 25968 13626
rect 26020 13574 26032 13626
rect 26084 13574 30820 13626
rect 1104 13552 30820 13574
rect 22186 13512 22192 13524
rect 21100 13484 22192 13512
rect 20346 13336 20352 13388
rect 20404 13376 20410 13388
rect 20404 13348 20760 13376
rect 20404 13336 20410 13348
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 20530 13308 20536 13320
rect 1443 13280 20536 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20732 13317 20760 13348
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 20810 13311 20868 13317
rect 20810 13277 20822 13311
rect 20856 13277 20868 13311
rect 20810 13271 20868 13277
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 21100 13308 21128 13484
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 23198 13512 23204 13524
rect 23159 13484 23204 13512
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 24394 13512 24400 13524
rect 24355 13484 24400 13512
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 26602 13472 26608 13524
rect 26660 13512 26666 13524
rect 27430 13512 27436 13524
rect 26660 13484 27436 13512
rect 26660 13472 26666 13484
rect 27430 13472 27436 13484
rect 27488 13472 27494 13524
rect 28718 13512 28724 13524
rect 28460 13484 28724 13512
rect 22922 13404 22928 13456
rect 22980 13444 22986 13456
rect 28353 13447 28411 13453
rect 28353 13444 28365 13447
rect 22980 13416 28365 13444
rect 22980 13404 22986 13416
rect 28353 13413 28365 13416
rect 28399 13413 28411 13447
rect 28353 13407 28411 13413
rect 24118 13336 24124 13388
rect 24176 13376 24182 13388
rect 25130 13376 25136 13388
rect 24176 13348 25136 13376
rect 24176 13336 24182 13348
rect 21266 13317 21272 13320
rect 21039 13280 21128 13308
rect 21223 13311 21272 13317
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 21223 13277 21235 13311
rect 21269 13277 21272 13311
rect 21223 13271 21272 13277
rect 20622 13200 20628 13252
rect 20680 13240 20686 13252
rect 20824 13240 20852 13271
rect 21266 13268 21272 13271
rect 21324 13268 21330 13320
rect 21542 13268 21548 13320
rect 21600 13308 21606 13320
rect 21821 13311 21879 13317
rect 21821 13308 21833 13311
rect 21600 13280 21833 13308
rect 21600 13268 21606 13280
rect 21821 13277 21833 13280
rect 21867 13277 21879 13311
rect 23198 13308 23204 13320
rect 21821 13271 21879 13277
rect 21928 13280 23204 13308
rect 20680 13212 20852 13240
rect 21085 13243 21143 13249
rect 20680 13200 20686 13212
rect 21085 13209 21097 13243
rect 21131 13240 21143 13243
rect 21928 13240 21956 13280
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 24578 13308 24584 13320
rect 24539 13280 24584 13308
rect 24578 13268 24584 13280
rect 24636 13268 24642 13320
rect 24872 13317 24900 13348
rect 25130 13336 25136 13348
rect 25188 13336 25194 13388
rect 26234 13376 26240 13388
rect 25332 13348 26240 13376
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13308 25099 13311
rect 25332 13308 25360 13348
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 26694 13336 26700 13388
rect 26752 13376 26758 13388
rect 27525 13379 27583 13385
rect 27525 13376 27537 13379
rect 26752 13348 27537 13376
rect 26752 13336 26758 13348
rect 27525 13345 27537 13348
rect 27571 13345 27583 13379
rect 27525 13339 27583 13345
rect 27709 13379 27767 13385
rect 27709 13345 27721 13379
rect 27755 13376 27767 13379
rect 28460 13376 28488 13484
rect 28718 13472 28724 13484
rect 28776 13472 28782 13524
rect 31386 13444 31392 13456
rect 27755 13348 28488 13376
rect 28552 13416 31392 13444
rect 27755 13345 27767 13348
rect 27709 13339 27767 13345
rect 25087 13280 25360 13308
rect 25087 13277 25099 13280
rect 25041 13271 25099 13277
rect 25406 13268 25412 13320
rect 25464 13308 25470 13320
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 25464 13280 26065 13308
rect 25464 13268 25470 13280
rect 26053 13277 26065 13280
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 26142 13268 26148 13320
rect 26200 13308 26206 13320
rect 26421 13311 26479 13317
rect 26421 13308 26433 13311
rect 26200 13280 26433 13308
rect 26200 13268 26206 13280
rect 26421 13277 26433 13280
rect 26467 13277 26479 13311
rect 26421 13271 26479 13277
rect 26786 13268 26792 13320
rect 26844 13308 26850 13320
rect 27433 13311 27491 13317
rect 27433 13308 27445 13311
rect 26844 13280 27445 13308
rect 26844 13268 26850 13280
rect 27433 13277 27445 13280
rect 27479 13277 27491 13311
rect 28552 13308 28580 13416
rect 31386 13404 31392 13416
rect 31444 13404 31450 13456
rect 28718 13336 28724 13388
rect 28776 13376 28782 13388
rect 28905 13379 28963 13385
rect 28905 13376 28917 13379
rect 28776 13348 28917 13376
rect 28776 13336 28782 13348
rect 28905 13345 28917 13348
rect 28951 13376 28963 13379
rect 30101 13379 30159 13385
rect 30101 13376 30113 13379
rect 28951 13348 30113 13376
rect 28951 13345 28963 13348
rect 28905 13339 28963 13345
rect 30101 13345 30113 13348
rect 30147 13345 30159 13379
rect 30101 13339 30159 13345
rect 27433 13271 27491 13277
rect 28092 13280 28580 13308
rect 28629 13311 28687 13317
rect 21131 13212 21956 13240
rect 22088 13243 22146 13249
rect 21131 13209 21143 13212
rect 21085 13203 21143 13209
rect 22088 13209 22100 13243
rect 22134 13240 22146 13243
rect 22646 13240 22652 13252
rect 22134 13212 22652 13240
rect 22134 13209 22146 13212
rect 22088 13203 22146 13209
rect 22646 13200 22652 13212
rect 22704 13200 22710 13252
rect 26234 13240 26240 13252
rect 26195 13212 26240 13240
rect 26234 13200 26240 13212
rect 26292 13200 26298 13252
rect 26329 13243 26387 13249
rect 26329 13209 26341 13243
rect 26375 13240 26387 13243
rect 26694 13240 26700 13252
rect 26375 13212 26700 13240
rect 26375 13209 26387 13212
rect 26329 13203 26387 13209
rect 26694 13200 26700 13212
rect 26752 13200 26758 13252
rect 28092 13240 28120 13280
rect 28629 13277 28641 13311
rect 28675 13308 28687 13311
rect 30006 13308 30012 13320
rect 28675 13280 30012 13308
rect 28675 13277 28687 13280
rect 28629 13271 28687 13277
rect 30006 13268 30012 13280
rect 30064 13268 30070 13320
rect 26896 13212 28120 13240
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19518 13172 19524 13184
rect 19392 13144 19524 13172
rect 19392 13132 19398 13144
rect 19518 13132 19524 13144
rect 19576 13132 19582 13184
rect 21358 13172 21364 13184
rect 21319 13144 21364 13172
rect 21358 13132 21364 13144
rect 21416 13132 21422 13184
rect 24210 13132 24216 13184
rect 24268 13172 24274 13184
rect 25498 13172 25504 13184
rect 24268 13144 25504 13172
rect 24268 13132 24274 13144
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 26605 13175 26663 13181
rect 26605 13141 26617 13175
rect 26651 13172 26663 13175
rect 26896 13172 26924 13212
rect 28166 13200 28172 13252
rect 28224 13240 28230 13252
rect 29917 13243 29975 13249
rect 29917 13240 29929 13243
rect 28224 13212 29929 13240
rect 28224 13200 28230 13212
rect 29917 13209 29929 13212
rect 29963 13209 29975 13243
rect 29917 13203 29975 13209
rect 27062 13172 27068 13184
rect 26651 13144 26924 13172
rect 27023 13144 27068 13172
rect 26651 13141 26663 13144
rect 26605 13135 26663 13141
rect 27062 13132 27068 13144
rect 27120 13132 27126 13184
rect 27430 13132 27436 13184
rect 27488 13172 27494 13184
rect 28813 13175 28871 13181
rect 28813 13172 28825 13175
rect 27488 13144 28825 13172
rect 27488 13132 27494 13144
rect 28813 13141 28825 13144
rect 28859 13141 28871 13175
rect 28813 13135 28871 13141
rect 1104 13082 30820 13104
rect 1104 13030 10880 13082
rect 10932 13030 10944 13082
rect 10996 13030 11008 13082
rect 11060 13030 11072 13082
rect 11124 13030 11136 13082
rect 11188 13030 20811 13082
rect 20863 13030 20875 13082
rect 20927 13030 20939 13082
rect 20991 13030 21003 13082
rect 21055 13030 21067 13082
rect 21119 13030 30820 13082
rect 1104 13008 30820 13030
rect 20622 12968 20628 12980
rect 20583 12940 20628 12968
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 22278 12968 22284 12980
rect 22152 12940 22284 12968
rect 22152 12928 22158 12940
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 22646 12928 22652 12980
rect 22704 12968 22710 12980
rect 22741 12971 22799 12977
rect 22741 12968 22753 12971
rect 22704 12940 22753 12968
rect 22704 12928 22710 12940
rect 22741 12937 22753 12940
rect 22787 12937 22799 12971
rect 22741 12931 22799 12937
rect 24673 12971 24731 12977
rect 24673 12937 24685 12971
rect 24719 12968 24731 12971
rect 24854 12968 24860 12980
rect 24719 12940 24860 12968
rect 24719 12937 24731 12940
rect 24673 12931 24731 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 25406 12928 25412 12980
rect 25464 12968 25470 12980
rect 26326 12968 26332 12980
rect 25464 12940 26332 12968
rect 25464 12928 25470 12940
rect 26326 12928 26332 12940
rect 26384 12928 26390 12980
rect 27246 12928 27252 12980
rect 27304 12968 27310 12980
rect 28258 12968 28264 12980
rect 27304 12940 28264 12968
rect 27304 12928 27310 12940
rect 28258 12928 28264 12940
rect 28316 12928 28322 12980
rect 28350 12928 28356 12980
rect 28408 12968 28414 12980
rect 28629 12971 28687 12977
rect 28629 12968 28641 12971
rect 28408 12940 28641 12968
rect 28408 12928 28414 12940
rect 28629 12937 28641 12940
rect 28675 12937 28687 12971
rect 28629 12931 28687 12937
rect 2038 12860 2044 12912
rect 2096 12900 2102 12912
rect 27617 12903 27675 12909
rect 27617 12900 27629 12903
rect 2096 12872 27629 12900
rect 2096 12860 2102 12872
rect 27617 12869 27629 12872
rect 27663 12869 27675 12903
rect 28442 12900 28448 12912
rect 28403 12872 28448 12900
rect 27617 12863 27675 12869
rect 28442 12860 28448 12872
rect 28500 12860 28506 12912
rect 28718 12900 28724 12912
rect 28679 12872 28724 12900
rect 28718 12860 28724 12872
rect 28776 12860 28782 12912
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 20548 12764 20576 12795
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 20717 12835 20775 12841
rect 20717 12832 20729 12835
rect 20680 12804 20729 12832
rect 20680 12792 20686 12804
rect 20717 12801 20729 12804
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 22925 12835 22983 12841
rect 22925 12801 22937 12835
rect 22971 12832 22983 12835
rect 23750 12832 23756 12844
rect 22971 12804 23756 12832
rect 22971 12801 22983 12804
rect 22925 12795 22983 12801
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 24854 12832 24860 12844
rect 24767 12804 24860 12832
rect 24854 12792 24860 12804
rect 24912 12832 24918 12844
rect 25406 12832 25412 12844
rect 24912 12804 25412 12832
rect 24912 12792 24918 12804
rect 25406 12792 25412 12804
rect 25464 12792 25470 12844
rect 25498 12792 25504 12844
rect 25556 12832 25562 12844
rect 25593 12835 25651 12841
rect 25593 12832 25605 12835
rect 25556 12804 25605 12832
rect 25556 12792 25562 12804
rect 25593 12801 25605 12804
rect 25639 12832 25651 12835
rect 26326 12832 26332 12844
rect 25639 12804 26332 12832
rect 25639 12801 25651 12804
rect 25593 12795 25651 12801
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 27430 12832 27436 12844
rect 27391 12804 27436 12832
rect 27430 12792 27436 12804
rect 27488 12792 27494 12844
rect 20806 12764 20812 12776
rect 20548 12736 20812 12764
rect 20806 12724 20812 12736
rect 20864 12764 20870 12776
rect 21266 12764 21272 12776
rect 20864 12736 21272 12764
rect 20864 12724 20870 12736
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 23106 12764 23112 12776
rect 23067 12736 23112 12764
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 23198 12724 23204 12776
rect 23256 12764 23262 12776
rect 23256 12736 23301 12764
rect 23256 12724 23262 12736
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 23440 12736 25145 12764
rect 23440 12724 23446 12736
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 29273 12767 29331 12773
rect 29273 12733 29285 12767
rect 29319 12764 29331 12767
rect 29362 12764 29368 12776
rect 29319 12736 29368 12764
rect 29319 12733 29331 12736
rect 29273 12727 29331 12733
rect 29362 12724 29368 12736
rect 29420 12724 29426 12776
rect 29546 12764 29552 12776
rect 29507 12736 29552 12764
rect 29546 12724 29552 12736
rect 29604 12724 29610 12776
rect 2314 12656 2320 12708
rect 2372 12696 2378 12708
rect 28169 12699 28227 12705
rect 28169 12696 28181 12699
rect 2372 12668 28181 12696
rect 2372 12656 2378 12668
rect 28169 12665 28181 12668
rect 28215 12665 28227 12699
rect 28169 12659 28227 12665
rect 25038 12628 25044 12640
rect 24999 12600 25044 12628
rect 25038 12588 25044 12600
rect 25096 12628 25102 12640
rect 25823 12631 25881 12637
rect 25823 12628 25835 12631
rect 25096 12600 25835 12628
rect 25096 12588 25102 12600
rect 25823 12597 25835 12600
rect 25869 12597 25881 12631
rect 25823 12591 25881 12597
rect 1104 12538 30820 12560
rect 1104 12486 5915 12538
rect 5967 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 15846 12538
rect 15898 12486 15910 12538
rect 15962 12486 15974 12538
rect 16026 12486 16038 12538
rect 16090 12486 16102 12538
rect 16154 12486 25776 12538
rect 25828 12486 25840 12538
rect 25892 12486 25904 12538
rect 25956 12486 25968 12538
rect 26020 12486 26032 12538
rect 26084 12486 30820 12538
rect 1104 12464 30820 12486
rect 2038 12424 2044 12436
rect 1999 12396 2044 12424
rect 2038 12384 2044 12396
rect 2096 12384 2102 12436
rect 25777 12427 25835 12433
rect 25777 12393 25789 12427
rect 25823 12424 25835 12427
rect 26418 12424 26424 12436
rect 25823 12396 26424 12424
rect 25823 12393 25835 12396
rect 25777 12387 25835 12393
rect 26418 12384 26424 12396
rect 26476 12384 26482 12436
rect 26973 12427 27031 12433
rect 26973 12393 26985 12427
rect 27019 12424 27031 12427
rect 27430 12424 27436 12436
rect 27019 12396 27436 12424
rect 27019 12393 27031 12396
rect 26973 12387 27031 12393
rect 27430 12384 27436 12396
rect 27488 12384 27494 12436
rect 26786 12316 26792 12368
rect 26844 12356 26850 12368
rect 30101 12359 30159 12365
rect 30101 12356 30113 12359
rect 26844 12328 30113 12356
rect 26844 12316 26850 12328
rect 30101 12325 30113 12328
rect 30147 12325 30159 12359
rect 30101 12319 30159 12325
rect 20346 12248 20352 12300
rect 20404 12288 20410 12300
rect 27522 12288 27528 12300
rect 20404 12260 21036 12288
rect 27483 12260 27528 12288
rect 20404 12248 20410 12260
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 2038 12220 2044 12232
rect 1443 12192 2044 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2682 12180 2688 12232
rect 2740 12220 2746 12232
rect 6270 12220 6276 12232
rect 2740 12192 6276 12220
rect 2740 12180 2746 12192
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18506 12220 18512 12232
rect 18003 12192 18512 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 20714 12220 20720 12232
rect 20675 12192 20720 12220
rect 20714 12180 20720 12192
rect 20772 12180 20778 12232
rect 21008 12229 21036 12260
rect 27522 12248 27528 12260
rect 27580 12248 27586 12300
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12189 20867 12223
rect 20809 12183 20867 12189
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12189 21051 12223
rect 20993 12183 21051 12189
rect 21085 12223 21143 12229
rect 21085 12189 21097 12223
rect 21131 12220 21143 12223
rect 21910 12220 21916 12232
rect 21131 12192 21916 12220
rect 21131 12189 21143 12192
rect 21085 12183 21143 12189
rect 20824 12152 20852 12183
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 23566 12180 23572 12232
rect 23624 12220 23630 12232
rect 25225 12223 25283 12229
rect 25225 12220 25237 12223
rect 23624 12192 25237 12220
rect 23624 12180 23630 12192
rect 25225 12189 25237 12192
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 25593 12223 25651 12229
rect 25593 12189 25605 12223
rect 25639 12220 25651 12223
rect 26142 12220 26148 12232
rect 25639 12192 26148 12220
rect 25639 12189 25651 12192
rect 25593 12183 25651 12189
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 28166 12220 28172 12232
rect 28127 12192 28172 12220
rect 28166 12180 28172 12192
rect 28224 12180 28230 12232
rect 22830 12152 22836 12164
rect 20824 12124 22836 12152
rect 22830 12112 22836 12124
rect 22888 12112 22894 12164
rect 24670 12112 24676 12164
rect 24728 12152 24734 12164
rect 25409 12155 25467 12161
rect 25409 12152 25421 12155
rect 24728 12124 25421 12152
rect 24728 12112 24734 12124
rect 25409 12121 25421 12124
rect 25455 12121 25467 12155
rect 25409 12115 25467 12121
rect 25501 12155 25559 12161
rect 25501 12121 25513 12155
rect 25547 12152 25559 12155
rect 25958 12152 25964 12164
rect 25547 12124 25964 12152
rect 25547 12121 25559 12124
rect 25501 12115 25559 12121
rect 25958 12112 25964 12124
rect 26016 12112 26022 12164
rect 26697 12155 26755 12161
rect 26697 12121 26709 12155
rect 26743 12152 26755 12155
rect 27433 12155 27491 12161
rect 27433 12152 27445 12155
rect 26743 12124 27445 12152
rect 26743 12121 26755 12124
rect 26697 12115 26755 12121
rect 27433 12121 27445 12124
rect 27479 12152 27491 12155
rect 29638 12152 29644 12164
rect 27479 12124 29644 12152
rect 27479 12121 27491 12124
rect 27433 12115 27491 12121
rect 29638 12112 29644 12124
rect 29696 12112 29702 12164
rect 29914 12152 29920 12164
rect 29875 12124 29920 12152
rect 29914 12112 29920 12124
rect 29972 12112 29978 12164
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 17494 12084 17500 12096
rect 17455 12056 17500 12084
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18141 12087 18199 12093
rect 18141 12084 18153 12087
rect 17920 12056 18153 12084
rect 17920 12044 17926 12056
rect 18141 12053 18153 12056
rect 18187 12053 18199 12087
rect 18141 12047 18199 12053
rect 20346 12044 20352 12096
rect 20404 12084 20410 12096
rect 20533 12087 20591 12093
rect 20533 12084 20545 12087
rect 20404 12056 20545 12084
rect 20404 12044 20410 12056
rect 20533 12053 20545 12056
rect 20579 12053 20591 12087
rect 20533 12047 20591 12053
rect 25038 12044 25044 12096
rect 25096 12084 25102 12096
rect 25866 12084 25872 12096
rect 25096 12056 25872 12084
rect 25096 12044 25102 12056
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 26878 12044 26884 12096
rect 26936 12084 26942 12096
rect 27341 12087 27399 12093
rect 27341 12084 27353 12087
rect 26936 12056 27353 12084
rect 26936 12044 26942 12056
rect 27341 12053 27353 12056
rect 27387 12084 27399 12087
rect 28399 12087 28457 12093
rect 28399 12084 28411 12087
rect 27387 12056 28411 12084
rect 27387 12053 27399 12056
rect 27341 12047 27399 12053
rect 28399 12053 28411 12056
rect 28445 12053 28457 12087
rect 28399 12047 28457 12053
rect 1104 11994 30820 12016
rect 1104 11942 10880 11994
rect 10932 11942 10944 11994
rect 10996 11942 11008 11994
rect 11060 11942 11072 11994
rect 11124 11942 11136 11994
rect 11188 11942 20811 11994
rect 20863 11942 20875 11994
rect 20927 11942 20939 11994
rect 20991 11942 21003 11994
rect 21055 11942 21067 11994
rect 21119 11942 30820 11994
rect 1104 11920 30820 11942
rect 19245 11883 19303 11889
rect 19245 11849 19257 11883
rect 19291 11880 19303 11883
rect 19334 11880 19340 11892
rect 19291 11852 19340 11880
rect 19291 11849 19303 11852
rect 19245 11843 19303 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20622 11880 20628 11892
rect 20036 11852 20628 11880
rect 20036 11840 20042 11852
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 25685 11883 25743 11889
rect 25685 11849 25697 11883
rect 25731 11880 25743 11883
rect 26234 11880 26240 11892
rect 25731 11852 26240 11880
rect 25731 11849 25743 11852
rect 25685 11843 25743 11849
rect 26234 11840 26240 11852
rect 26292 11840 26298 11892
rect 27614 11840 27620 11892
rect 27672 11840 27678 11892
rect 27798 11840 27804 11892
rect 27856 11880 27862 11892
rect 28629 11883 28687 11889
rect 28629 11880 28641 11883
rect 27856 11852 28641 11880
rect 27856 11840 27862 11852
rect 28629 11849 28641 11852
rect 28675 11849 28687 11883
rect 28629 11843 28687 11849
rect 4798 11772 4804 11824
rect 4856 11812 4862 11824
rect 27632 11812 27660 11840
rect 4856 11784 21496 11812
rect 4856 11772 4862 11784
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 17862 11744 17868 11756
rect 17823 11716 17868 11744
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 18132 11747 18190 11753
rect 18132 11713 18144 11747
rect 18178 11744 18190 11747
rect 19242 11744 19248 11756
rect 18178 11716 19248 11744
rect 18178 11713 18190 11716
rect 18132 11707 18190 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 19978 11744 19984 11756
rect 19939 11716 19984 11744
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11744 20223 11747
rect 20254 11744 20260 11756
rect 20211 11716 20260 11744
rect 20211 11713 20223 11716
rect 20165 11707 20223 11713
rect 19610 11636 19616 11688
rect 19668 11676 19674 11688
rect 19794 11676 19800 11688
rect 19668 11648 19800 11676
rect 19668 11636 19674 11648
rect 19794 11636 19800 11648
rect 19852 11676 19858 11688
rect 20088 11676 20116 11707
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11744 20407 11747
rect 21358 11744 21364 11756
rect 20395 11716 21364 11744
rect 20395 11713 20407 11716
rect 20349 11707 20407 11713
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 19852 11648 20116 11676
rect 19852 11636 19858 11648
rect 21468 11608 21496 11784
rect 22066 11784 27660 11812
rect 27709 11815 27767 11821
rect 22066 11608 22094 11784
rect 27709 11781 27721 11815
rect 27755 11812 27767 11815
rect 28353 11815 28411 11821
rect 28353 11812 28365 11815
rect 27755 11784 28365 11812
rect 27755 11781 27767 11784
rect 27709 11775 27767 11781
rect 28353 11781 28365 11784
rect 28399 11812 28411 11815
rect 29730 11812 29736 11824
rect 28399 11784 29736 11812
rect 28399 11781 28411 11784
rect 28353 11775 28411 11781
rect 29730 11772 29736 11784
rect 29788 11772 29794 11824
rect 24854 11744 24860 11756
rect 24815 11716 24860 11744
rect 24854 11704 24860 11716
rect 24912 11744 24918 11756
rect 25869 11747 25927 11753
rect 25869 11744 25881 11747
rect 24912 11716 25881 11744
rect 24912 11704 24918 11716
rect 25869 11713 25881 11716
rect 25915 11713 25927 11747
rect 25869 11707 25927 11713
rect 25958 11704 25964 11756
rect 26016 11744 26022 11756
rect 27617 11747 27675 11753
rect 27617 11744 27629 11747
rect 26016 11716 27629 11744
rect 26016 11704 26022 11716
rect 27617 11713 27629 11716
rect 27663 11744 27675 11747
rect 28810 11744 28816 11756
rect 27663 11716 27936 11744
rect 28771 11716 28816 11744
rect 27663 11713 27675 11716
rect 27617 11707 27675 11713
rect 25038 11676 25044 11688
rect 24999 11648 25044 11676
rect 25038 11636 25044 11648
rect 25096 11636 25102 11688
rect 25133 11679 25191 11685
rect 25133 11645 25145 11679
rect 25179 11676 25191 11679
rect 25179 11648 25360 11676
rect 25179 11645 25191 11648
rect 25133 11639 25191 11645
rect 21468 11580 22094 11608
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 19702 11540 19708 11552
rect 19663 11512 19708 11540
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 23198 11500 23204 11552
rect 23256 11540 23262 11552
rect 25332 11540 25360 11648
rect 25406 11636 25412 11688
rect 25464 11676 25470 11688
rect 25976 11676 26004 11704
rect 25464 11648 26004 11676
rect 26145 11679 26203 11685
rect 25464 11636 25470 11648
rect 26145 11645 26157 11679
rect 26191 11645 26203 11679
rect 26145 11639 26203 11645
rect 27801 11679 27859 11685
rect 27801 11645 27813 11679
rect 27847 11645 27859 11679
rect 27908 11676 27936 11716
rect 28810 11704 28816 11716
rect 28868 11704 28874 11756
rect 29454 11744 29460 11756
rect 28920 11716 29460 11744
rect 28920 11676 28948 11716
rect 29454 11704 29460 11716
rect 29512 11704 29518 11756
rect 29270 11676 29276 11688
rect 27908 11648 28948 11676
rect 29231 11648 29276 11676
rect 27801 11639 27859 11645
rect 25866 11568 25872 11620
rect 25924 11608 25930 11620
rect 26053 11611 26111 11617
rect 26053 11608 26065 11611
rect 25924 11580 26065 11608
rect 25924 11568 25930 11580
rect 26053 11577 26065 11580
rect 26099 11577 26111 11611
rect 26053 11571 26111 11577
rect 23256 11512 25360 11540
rect 23256 11500 23262 11512
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 26160 11540 26188 11639
rect 26694 11568 26700 11620
rect 26752 11608 26758 11620
rect 26752 11580 27476 11608
rect 26752 11568 26758 11580
rect 25556 11512 26188 11540
rect 25556 11500 25562 11512
rect 26602 11500 26608 11552
rect 26660 11540 26666 11552
rect 27249 11543 27307 11549
rect 27249 11540 27261 11543
rect 26660 11512 27261 11540
rect 26660 11500 26666 11512
rect 27249 11509 27261 11512
rect 27295 11509 27307 11543
rect 27448 11540 27476 11580
rect 27522 11568 27528 11620
rect 27580 11608 27586 11620
rect 27816 11608 27844 11639
rect 29270 11636 29276 11648
rect 29328 11636 29334 11688
rect 29549 11679 29607 11685
rect 29549 11645 29561 11679
rect 29595 11645 29607 11679
rect 29549 11639 29607 11645
rect 29564 11608 29592 11639
rect 27580 11580 27844 11608
rect 27908 11580 29592 11608
rect 27580 11568 27586 11580
rect 27908 11540 27936 11580
rect 27448 11512 27936 11540
rect 27249 11503 27307 11509
rect 1104 11450 30820 11472
rect 1104 11398 5915 11450
rect 5967 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 15846 11450
rect 15898 11398 15910 11450
rect 15962 11398 15974 11450
rect 16026 11398 16038 11450
rect 16090 11398 16102 11450
rect 16154 11398 25776 11450
rect 25828 11398 25840 11450
rect 25892 11398 25904 11450
rect 25956 11398 25968 11450
rect 26020 11398 26032 11450
rect 26084 11398 30820 11450
rect 1104 11376 30820 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 19242 11336 19248 11348
rect 1452 11308 6914 11336
rect 19203 11308 19248 11336
rect 1452 11296 1458 11308
rect 6886 11268 6914 11308
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21269 11339 21327 11345
rect 21269 11336 21281 11339
rect 21232 11308 21281 11336
rect 21232 11296 21238 11308
rect 21269 11305 21281 11308
rect 21315 11305 21327 11339
rect 21269 11299 21327 11305
rect 21358 11296 21364 11348
rect 21416 11336 21422 11348
rect 26697 11339 26755 11345
rect 26697 11336 26709 11339
rect 21416 11308 26709 11336
rect 21416 11296 21422 11308
rect 26697 11305 26709 11308
rect 26743 11305 26755 11339
rect 26697 11299 26755 11305
rect 27522 11296 27528 11348
rect 27580 11336 27586 11348
rect 28169 11339 28227 11345
rect 28169 11336 28181 11339
rect 27580 11308 28181 11336
rect 27580 11296 27586 11308
rect 28169 11305 28181 11308
rect 28215 11305 28227 11339
rect 28169 11299 28227 11305
rect 28442 11296 28448 11348
rect 28500 11336 28506 11348
rect 28905 11339 28963 11345
rect 28905 11336 28917 11339
rect 28500 11308 28917 11336
rect 28500 11296 28506 11308
rect 28905 11305 28917 11308
rect 28951 11305 28963 11339
rect 28905 11299 28963 11305
rect 30009 11339 30067 11345
rect 30009 11305 30021 11339
rect 30055 11336 30067 11339
rect 30098 11336 30104 11348
rect 30055 11308 30104 11336
rect 30055 11305 30067 11308
rect 30009 11299 30067 11305
rect 30098 11296 30104 11308
rect 30156 11296 30162 11348
rect 19610 11268 19616 11280
rect 6886 11240 19616 11268
rect 19610 11228 19616 11240
rect 19668 11228 19674 11280
rect 20162 11200 20168 11212
rect 19720 11172 20168 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 2314 11132 2320 11144
rect 2275 11104 2320 11132
rect 1397 11095 1455 11101
rect 1412 11064 1440 11095
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 19426 11092 19432 11144
rect 19484 11141 19490 11144
rect 19720 11141 19748 11172
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 20312 11172 20821 11200
rect 20312 11160 20318 11172
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 20809 11163 20867 11169
rect 20901 11203 20959 11209
rect 20901 11169 20913 11203
rect 20947 11200 20959 11203
rect 21634 11200 21640 11212
rect 20947 11172 21640 11200
rect 20947 11169 20959 11172
rect 20901 11163 20959 11169
rect 21634 11160 21640 11172
rect 21692 11160 21698 11212
rect 25130 11200 25136 11212
rect 24872 11172 25136 11200
rect 19484 11135 19533 11141
rect 19484 11101 19487 11135
rect 19521 11101 19533 11135
rect 19484 11095 19533 11101
rect 19594 11135 19652 11141
rect 19594 11101 19606 11135
rect 19640 11134 19652 11135
rect 19705 11135 19763 11141
rect 19640 11132 19656 11134
rect 19640 11101 19657 11132
rect 19594 11095 19657 11101
rect 19705 11101 19717 11135
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 19901 11135 19959 11141
rect 19901 11101 19913 11135
rect 19947 11132 19959 11135
rect 20346 11132 20352 11144
rect 19947 11104 20352 11132
rect 19947 11101 19959 11104
rect 19901 11095 19959 11101
rect 19484 11092 19490 11095
rect 19629 11064 19657 11095
rect 20346 11092 20352 11104
rect 20404 11092 20410 11144
rect 20533 11135 20591 11141
rect 20533 11101 20545 11135
rect 20579 11101 20591 11135
rect 20533 11095 20591 11101
rect 19794 11064 19800 11076
rect 1412 11036 2728 11064
rect 19629 11036 19800 11064
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 2700 10996 2728 11036
rect 19794 11024 19800 11036
rect 19852 11024 19858 11076
rect 20548 11064 20576 11095
rect 20622 11092 20628 11144
rect 20680 11132 20686 11144
rect 20717 11135 20775 11141
rect 20717 11132 20729 11135
rect 20680 11104 20729 11132
rect 20680 11092 20686 11104
rect 20717 11101 20729 11104
rect 20763 11101 20775 11135
rect 20717 11095 20775 11101
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 23198 11132 23204 11144
rect 21131 11104 23204 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 24026 11092 24032 11144
rect 24084 11132 24090 11144
rect 24394 11132 24400 11144
rect 24084 11104 24400 11132
rect 24084 11092 24090 11104
rect 24394 11092 24400 11104
rect 24452 11132 24458 11144
rect 24872 11141 24900 11172
rect 25130 11160 25136 11172
rect 25188 11200 25194 11212
rect 25777 11203 25835 11209
rect 25777 11200 25789 11203
rect 25188 11172 25789 11200
rect 25188 11160 25194 11172
rect 25777 11169 25789 11172
rect 25823 11169 25835 11203
rect 25777 11163 25835 11169
rect 27154 11160 27160 11212
rect 27212 11200 27218 11212
rect 27430 11200 27436 11212
rect 27212 11172 27436 11200
rect 27212 11160 27218 11172
rect 27430 11160 27436 11172
rect 27488 11160 27494 11212
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 24452 11104 24593 11132
rect 24452 11092 24458 11104
rect 24581 11101 24593 11104
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 24857 11095 24915 11101
rect 25041 11135 25099 11141
rect 25041 11101 25053 11135
rect 25087 11101 25099 11135
rect 25041 11095 25099 11101
rect 21174 11064 21180 11076
rect 20548 11036 21180 11064
rect 21174 11024 21180 11036
rect 21232 11064 21238 11076
rect 21450 11064 21456 11076
rect 21232 11036 21456 11064
rect 21232 11024 21238 11036
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 22830 11024 22836 11076
rect 22888 11064 22894 11076
rect 23014 11064 23020 11076
rect 22888 11036 23020 11064
rect 22888 11024 22894 11036
rect 23014 11024 23020 11036
rect 23072 11024 23078 11076
rect 25056 11064 25084 11095
rect 25314 11092 25320 11144
rect 25372 11132 25378 11144
rect 25593 11135 25651 11141
rect 25593 11132 25605 11135
rect 25372 11104 25605 11132
rect 25372 11092 25378 11104
rect 25593 11101 25605 11104
rect 25639 11101 25651 11135
rect 26602 11132 26608 11144
rect 26563 11104 26608 11132
rect 25593 11095 25651 11101
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 28077 11135 28135 11141
rect 28077 11101 28089 11135
rect 28123 11132 28135 11135
rect 28258 11132 28264 11144
rect 28123 11104 28264 11132
rect 28123 11101 28135 11104
rect 28077 11095 28135 11101
rect 28258 11092 28264 11104
rect 28316 11092 28322 11144
rect 28718 11132 28724 11144
rect 28679 11104 28724 11132
rect 28718 11092 28724 11104
rect 28776 11092 28782 11144
rect 28902 11092 28908 11144
rect 28960 11132 28966 11144
rect 29825 11135 29883 11141
rect 29825 11132 29837 11135
rect 28960 11104 29837 11132
rect 28960 11092 28966 11104
rect 29825 11101 29837 11104
rect 29871 11101 29883 11135
rect 29825 11095 29883 11101
rect 25406 11064 25412 11076
rect 25056 11036 25412 11064
rect 25406 11024 25412 11036
rect 25464 11024 25470 11076
rect 25682 11024 25688 11076
rect 25740 11064 25746 11076
rect 26234 11064 26240 11076
rect 25740 11036 26240 11064
rect 25740 11024 25746 11036
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 24210 10996 24216 11008
rect 2700 10968 24216 10996
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 24394 10996 24400 11008
rect 24355 10968 24400 10996
rect 24394 10956 24400 10968
rect 24452 10956 24458 11008
rect 1104 10906 30820 10928
rect 1104 10854 10880 10906
rect 10932 10854 10944 10906
rect 10996 10854 11008 10906
rect 11060 10854 11072 10906
rect 11124 10854 11136 10906
rect 11188 10854 20811 10906
rect 20863 10854 20875 10906
rect 20927 10854 20939 10906
rect 20991 10854 21003 10906
rect 21055 10854 21067 10906
rect 21119 10854 30820 10906
rect 1104 10832 30820 10854
rect 19245 10795 19303 10801
rect 19245 10761 19257 10795
rect 19291 10792 19303 10795
rect 20346 10792 20352 10804
rect 19291 10764 20352 10792
rect 19291 10761 19303 10764
rect 19245 10755 19303 10761
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 23198 10792 23204 10804
rect 23159 10764 23204 10792
rect 23198 10752 23204 10764
rect 23256 10752 23262 10804
rect 25130 10792 25136 10804
rect 24136 10764 25136 10792
rect 17954 10724 17960 10736
rect 6886 10696 17960 10724
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 6886 10656 6914 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18132 10727 18190 10733
rect 18132 10693 18144 10727
rect 18178 10724 18190 10727
rect 19702 10724 19708 10736
rect 18178 10696 19708 10724
rect 18178 10693 18190 10696
rect 18132 10687 18190 10693
rect 19702 10684 19708 10696
rect 19760 10684 19766 10736
rect 20438 10724 20444 10736
rect 20088 10696 20444 10724
rect 1443 10628 6914 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17552 10628 17877 10656
rect 17552 10616 17558 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 20088 10665 20116 10696
rect 20438 10684 20444 10696
rect 20496 10724 20502 10736
rect 20496 10696 21312 10724
rect 20496 10684 20502 10696
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 19484 10628 20085 10656
rect 19484 10616 19490 10628
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 21284 10665 21312 10696
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 20588 10628 21097 10656
rect 20588 10616 20594 10628
rect 21085 10625 21097 10628
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 22088 10659 22146 10665
rect 22088 10625 22100 10659
rect 22134 10656 22146 10659
rect 22646 10656 22652 10668
rect 22134 10628 22652 10656
rect 22134 10625 22146 10628
rect 22088 10619 22146 10625
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 24026 10656 24032 10668
rect 23987 10628 24032 10656
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 24136 10656 24164 10764
rect 25130 10752 25136 10764
rect 25188 10752 25194 10804
rect 27065 10795 27123 10801
rect 27065 10792 27077 10795
rect 26252 10764 27077 10792
rect 24210 10684 24216 10736
rect 24268 10724 24274 10736
rect 26252 10733 26280 10764
rect 27065 10761 27077 10764
rect 27111 10761 27123 10795
rect 27065 10755 27123 10761
rect 27525 10795 27583 10801
rect 27525 10761 27537 10795
rect 27571 10792 27583 10795
rect 28074 10792 28080 10804
rect 27571 10764 28080 10792
rect 27571 10761 27583 10764
rect 27525 10755 27583 10761
rect 28074 10752 28080 10764
rect 28132 10752 28138 10804
rect 29362 10792 29368 10804
rect 29323 10764 29368 10792
rect 29362 10752 29368 10764
rect 29420 10792 29426 10804
rect 30650 10792 30656 10804
rect 29420 10764 30656 10792
rect 29420 10752 29426 10764
rect 30650 10752 30656 10764
rect 30708 10752 30714 10804
rect 26237 10727 26295 10733
rect 24268 10696 24624 10724
rect 24268 10684 24274 10696
rect 24305 10659 24363 10665
rect 24305 10656 24317 10659
rect 24136 10628 24317 10656
rect 24305 10625 24317 10628
rect 24351 10625 24363 10659
rect 24305 10619 24363 10625
rect 24489 10659 24547 10665
rect 24489 10625 24501 10659
rect 24535 10625 24547 10659
rect 24596 10656 24624 10696
rect 26237 10693 26249 10727
rect 26283 10693 26295 10727
rect 26237 10687 26295 10693
rect 27614 10684 27620 10736
rect 27672 10724 27678 10736
rect 28353 10727 28411 10733
rect 28353 10724 28365 10727
rect 27672 10696 28365 10724
rect 27672 10684 27678 10696
rect 28353 10693 28365 10696
rect 28399 10693 28411 10727
rect 28353 10687 28411 10693
rect 26421 10659 26479 10665
rect 26421 10656 26433 10659
rect 24596 10628 26433 10656
rect 24489 10619 24547 10625
rect 26421 10625 26433 10628
rect 26467 10625 26479 10659
rect 26421 10619 26479 10625
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19797 10591 19855 10597
rect 19797 10588 19809 10591
rect 19392 10560 19809 10588
rect 19392 10548 19398 10560
rect 19797 10557 19809 10560
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 21821 10591 21879 10597
rect 21821 10588 21833 10591
rect 21600 10560 21833 10588
rect 21600 10548 21606 10560
rect 21821 10557 21833 10560
rect 21867 10557 21879 10591
rect 21821 10551 21879 10557
rect 24504 10520 24532 10619
rect 26786 10616 26792 10668
rect 26844 10656 26850 10668
rect 27433 10659 27491 10665
rect 27433 10656 27445 10659
rect 26844 10628 27445 10656
rect 26844 10616 26850 10628
rect 27433 10625 27445 10628
rect 27479 10625 27491 10659
rect 27433 10619 27491 10625
rect 27522 10548 27528 10600
rect 27580 10588 27586 10600
rect 27617 10591 27675 10597
rect 27617 10588 27629 10591
rect 27580 10560 27629 10588
rect 27580 10548 27586 10560
rect 27617 10557 27629 10560
rect 27663 10557 27675 10591
rect 27617 10551 27675 10557
rect 26878 10520 26884 10532
rect 24504 10492 26884 10520
rect 26878 10480 26884 10492
rect 26936 10480 26942 10532
rect 27246 10480 27252 10532
rect 27304 10520 27310 10532
rect 29104 10520 29132 10642
rect 29178 10548 29184 10600
rect 29236 10588 29242 10600
rect 29236 10560 29394 10588
rect 29236 10548 29242 10560
rect 27304 10492 29132 10520
rect 27304 10480 27310 10492
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 21085 10455 21143 10461
rect 21085 10421 21097 10455
rect 21131 10452 21143 10455
rect 21450 10452 21456 10464
rect 21131 10424 21456 10452
rect 21131 10421 21143 10424
rect 21085 10415 21143 10421
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 23842 10452 23848 10464
rect 23803 10424 23848 10452
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 1104 10362 30820 10384
rect 1104 10310 5915 10362
rect 5967 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 15846 10362
rect 15898 10310 15910 10362
rect 15962 10310 15974 10362
rect 16026 10310 16038 10362
rect 16090 10310 16102 10362
rect 16154 10310 25776 10362
rect 25828 10310 25840 10362
rect 25892 10310 25904 10362
rect 25956 10310 25968 10362
rect 26020 10310 26032 10362
rect 26084 10310 30820 10362
rect 1104 10288 30820 10310
rect 21910 10248 21916 10260
rect 21871 10220 21916 10248
rect 21910 10208 21916 10220
rect 21968 10208 21974 10260
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 22741 10251 22799 10257
rect 22741 10248 22753 10251
rect 22704 10220 22753 10248
rect 22704 10208 22710 10220
rect 22741 10217 22753 10220
rect 22787 10217 22799 10251
rect 23106 10248 23112 10260
rect 23067 10220 23112 10248
rect 22741 10211 22799 10217
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 26326 10248 26332 10260
rect 26287 10220 26332 10248
rect 26326 10208 26332 10220
rect 26384 10208 26390 10260
rect 17954 10140 17960 10192
rect 18012 10180 18018 10192
rect 28077 10183 28135 10189
rect 28077 10180 28089 10183
rect 18012 10152 28089 10180
rect 18012 10140 18018 10152
rect 28077 10149 28089 10152
rect 28123 10149 28135 10183
rect 28077 10143 28135 10149
rect 20165 10115 20223 10121
rect 20165 10081 20177 10115
rect 20211 10112 20223 10115
rect 20530 10112 20536 10124
rect 20211 10084 20536 10112
rect 20211 10081 20223 10084
rect 20165 10075 20223 10081
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 21450 10112 21456 10124
rect 21411 10084 21456 10112
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 21545 10115 21603 10121
rect 21545 10081 21557 10115
rect 21591 10112 21603 10115
rect 21634 10112 21640 10124
rect 21591 10084 21640 10112
rect 21591 10081 21603 10084
rect 21545 10075 21603 10081
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 24394 10112 24400 10124
rect 22940 10084 24400 10112
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2130 10044 2136 10056
rect 1443 10016 2136 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2682 10044 2688 10056
rect 2363 10016 2688 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20346 10044 20352 10056
rect 19935 10016 20352 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 21174 10044 21180 10056
rect 21135 10016 21180 10044
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21358 10044 21364 10056
rect 21319 10016 21364 10044
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 22940 10053 22968 10084
rect 24394 10072 24400 10084
rect 24452 10072 24458 10124
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10013 21787 10047
rect 21729 10007 21787 10013
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10013 22983 10047
rect 23198 10044 23204 10056
rect 23159 10016 23204 10044
rect 22925 10007 22983 10013
rect 21744 9976 21772 10007
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 27062 10004 27068 10056
rect 27120 10044 27126 10056
rect 27893 10047 27951 10053
rect 27893 10044 27905 10047
rect 27120 10016 27905 10044
rect 27120 10004 27126 10016
rect 27893 10013 27905 10016
rect 27939 10013 27951 10047
rect 27893 10007 27951 10013
rect 28258 10004 28264 10056
rect 28316 10044 28322 10056
rect 28721 10047 28779 10053
rect 28721 10044 28733 10047
rect 28316 10016 28733 10044
rect 28316 10004 28322 10016
rect 28721 10013 28733 10016
rect 28767 10013 28779 10047
rect 28721 10007 28779 10013
rect 25498 9976 25504 9988
rect 21744 9948 25504 9976
rect 25498 9936 25504 9948
rect 25556 9936 25562 9988
rect 26234 9976 26240 9988
rect 26147 9948 26240 9976
rect 26234 9936 26240 9948
rect 26292 9976 26298 9988
rect 29730 9976 29736 9988
rect 26292 9948 28948 9976
rect 29691 9948 29736 9976
rect 26292 9936 26298 9948
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 2130 9908 2136 9920
rect 2091 9880 2136 9908
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 28810 9908 28816 9920
rect 28771 9880 28816 9908
rect 28810 9868 28816 9880
rect 28868 9868 28874 9920
rect 28920 9908 28948 9948
rect 29730 9936 29736 9948
rect 29788 9936 29794 9988
rect 29825 9911 29883 9917
rect 29825 9908 29837 9911
rect 28920 9880 29837 9908
rect 29825 9877 29837 9880
rect 29871 9877 29883 9911
rect 29825 9871 29883 9877
rect 1104 9818 30820 9840
rect 1104 9766 10880 9818
rect 10932 9766 10944 9818
rect 10996 9766 11008 9818
rect 11060 9766 11072 9818
rect 11124 9766 11136 9818
rect 11188 9766 20811 9818
rect 20863 9766 20875 9818
rect 20927 9766 20939 9818
rect 20991 9766 21003 9818
rect 21055 9766 21067 9818
rect 21119 9766 30820 9818
rect 1104 9744 30820 9766
rect 20346 9664 20352 9716
rect 20404 9704 20410 9716
rect 21269 9707 21327 9713
rect 20404 9676 20760 9704
rect 20404 9664 20410 9676
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 19981 9639 20039 9645
rect 7616 9608 19932 9636
rect 7616 9596 7622 9608
rect 2314 9392 2320 9444
rect 2372 9432 2378 9444
rect 19904 9432 19932 9608
rect 19981 9605 19993 9639
rect 20027 9636 20039 9639
rect 20622 9636 20628 9648
rect 20027 9608 20628 9636
rect 20027 9605 20039 9608
rect 19981 9599 20039 9605
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 20732 9636 20760 9676
rect 21269 9673 21281 9707
rect 21315 9704 21327 9707
rect 21358 9704 21364 9716
rect 21315 9676 21364 9704
rect 21315 9673 21327 9676
rect 21269 9667 21327 9673
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 24026 9664 24032 9716
rect 24084 9704 24090 9716
rect 24121 9707 24179 9713
rect 24121 9704 24133 9707
rect 24084 9676 24133 9704
rect 24084 9664 24090 9676
rect 24121 9673 24133 9676
rect 24167 9673 24179 9707
rect 24121 9667 24179 9673
rect 29365 9707 29423 9713
rect 29365 9673 29377 9707
rect 29411 9704 29423 9707
rect 29411 9676 29868 9704
rect 29411 9673 29423 9676
rect 29365 9667 29423 9673
rect 29840 9636 29868 9676
rect 30374 9636 30380 9648
rect 20732 9608 21128 9636
rect 29840 9608 30380 9636
rect 20162 9568 20168 9580
rect 20123 9540 20168 9568
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 20438 9568 20444 9580
rect 20399 9540 20444 9568
rect 20438 9528 20444 9540
rect 20496 9568 20502 9580
rect 21100 9577 21128 9608
rect 30374 9596 30380 9608
rect 30432 9636 30438 9648
rect 31846 9636 31852 9648
rect 30432 9608 31852 9636
rect 30432 9596 30438 9608
rect 31846 9596 31852 9608
rect 31904 9596 31910 9648
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20496 9540 20913 9568
rect 20496 9528 20502 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9537 21143 9571
rect 21085 9531 21143 9537
rect 22833 9571 22891 9577
rect 22833 9537 22845 9571
rect 22879 9568 22891 9571
rect 23842 9568 23848 9580
rect 22879 9540 23848 9568
rect 22879 9537 22891 9540
rect 22833 9531 22891 9537
rect 23842 9528 23848 9540
rect 23900 9528 23906 9580
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9568 24363 9571
rect 25590 9568 25596 9580
rect 24351 9540 25596 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 27062 9568 27068 9580
rect 27023 9540 27068 9568
rect 27062 9528 27068 9540
rect 27120 9528 27126 9580
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9568 27215 9571
rect 27430 9568 27436 9580
rect 27203 9540 27436 9568
rect 27203 9537 27215 9540
rect 27157 9531 27215 9537
rect 20349 9503 20407 9509
rect 20349 9469 20361 9503
rect 20395 9500 20407 9503
rect 20530 9500 20536 9512
rect 20395 9472 20536 9500
rect 20395 9469 20407 9472
rect 20349 9463 20407 9469
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 23109 9503 23167 9509
rect 23109 9469 23121 9503
rect 23155 9500 23167 9503
rect 23290 9500 23296 9512
rect 23155 9472 23296 9500
rect 23155 9469 23167 9472
rect 23109 9463 23167 9469
rect 23290 9460 23296 9472
rect 23348 9460 23354 9512
rect 26694 9460 26700 9512
rect 26752 9500 26758 9512
rect 27172 9500 27200 9531
rect 27430 9528 27436 9540
rect 27488 9528 27494 9580
rect 28626 9528 28632 9580
rect 28684 9568 28690 9580
rect 28684 9540 29118 9568
rect 28684 9528 28690 9540
rect 26752 9472 27200 9500
rect 28353 9503 28411 9509
rect 26752 9460 26758 9472
rect 28353 9469 28365 9503
rect 28399 9469 28411 9503
rect 28353 9463 28411 9469
rect 28368 9432 28396 9463
rect 29178 9460 29184 9512
rect 29236 9500 29242 9512
rect 29236 9472 29394 9500
rect 29236 9460 29242 9472
rect 2372 9404 6914 9432
rect 19904 9404 28396 9432
rect 2372 9392 2378 9404
rect 6886 9364 6914 9404
rect 22370 9364 22376 9376
rect 6886 9336 22376 9364
rect 22370 9324 22376 9336
rect 22428 9324 22434 9376
rect 22646 9364 22652 9376
rect 22607 9336 22652 9364
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23017 9367 23075 9373
rect 23017 9333 23029 9367
rect 23063 9364 23075 9367
rect 23106 9364 23112 9376
rect 23063 9336 23112 9364
rect 23063 9333 23075 9336
rect 23017 9327 23075 9333
rect 23106 9324 23112 9336
rect 23164 9324 23170 9376
rect 25314 9324 25320 9376
rect 25372 9364 25378 9376
rect 27065 9367 27123 9373
rect 27065 9364 27077 9367
rect 25372 9336 27077 9364
rect 25372 9324 25378 9336
rect 27065 9333 27077 9336
rect 27111 9333 27123 9367
rect 27065 9327 27123 9333
rect 1104 9274 30820 9296
rect 1104 9222 5915 9274
rect 5967 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 15846 9274
rect 15898 9222 15910 9274
rect 15962 9222 15974 9274
rect 16026 9222 16038 9274
rect 16090 9222 16102 9274
rect 16154 9222 25776 9274
rect 25828 9222 25840 9274
rect 25892 9222 25904 9274
rect 25956 9222 25968 9274
rect 26020 9222 26032 9274
rect 26084 9222 30820 9274
rect 1104 9200 30820 9222
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 20254 9160 20260 9172
rect 2740 9132 6914 9160
rect 20215 9132 20260 9160
rect 2740 9120 2746 9132
rect 6886 9024 6914 9132
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 22830 9160 22836 9172
rect 20548 9132 22836 9160
rect 20165 9095 20223 9101
rect 20165 9061 20177 9095
rect 20211 9092 20223 9095
rect 20438 9092 20444 9104
rect 20211 9064 20444 9092
rect 20211 9061 20223 9064
rect 20165 9055 20223 9061
rect 20438 9052 20444 9064
rect 20496 9052 20502 9104
rect 20548 9024 20576 9132
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 22925 9163 22983 9169
rect 22925 9129 22937 9163
rect 22971 9160 22983 9163
rect 23290 9160 23296 9172
rect 22971 9132 23296 9160
rect 22971 9129 22983 9132
rect 22925 9123 22983 9129
rect 23290 9120 23296 9132
rect 23348 9120 23354 9172
rect 30006 9160 30012 9172
rect 29967 9132 30012 9160
rect 30006 9120 30012 9132
rect 30064 9120 30070 9172
rect 27065 9095 27123 9101
rect 27065 9061 27077 9095
rect 27111 9092 27123 9095
rect 28718 9092 28724 9104
rect 27111 9064 28724 9092
rect 27111 9061 27123 9064
rect 27065 9055 27123 9061
rect 28718 9052 28724 9064
rect 28776 9052 28782 9104
rect 6886 8996 20576 9024
rect 24578 8984 24584 9036
rect 24636 9024 24642 9036
rect 25409 9027 25467 9033
rect 25409 9024 25421 9027
rect 24636 8996 25421 9024
rect 24636 8984 24642 8996
rect 25409 8993 25421 8996
rect 25455 8993 25467 9027
rect 25409 8987 25467 8993
rect 27709 9027 27767 9033
rect 27709 8993 27721 9027
rect 27755 9024 27767 9027
rect 28810 9024 28816 9036
rect 27755 8996 28816 9024
rect 27755 8993 27767 8996
rect 27709 8987 27767 8993
rect 28810 8984 28816 8996
rect 28868 8984 28874 9036
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 2130 8956 2136 8968
rect 1443 8928 2136 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 20073 8959 20131 8965
rect 20073 8925 20085 8959
rect 20119 8956 20131 8959
rect 20530 8956 20536 8968
rect 20119 8928 20536 8956
rect 20119 8925 20131 8928
rect 20073 8919 20131 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 21542 8956 21548 8968
rect 21503 8928 21548 8956
rect 21542 8916 21548 8928
rect 21600 8916 21606 8968
rect 21812 8959 21870 8965
rect 21812 8925 21824 8959
rect 21858 8956 21870 8959
rect 22646 8956 22652 8968
rect 21858 8928 22652 8956
rect 21858 8925 21870 8928
rect 21812 8919 21870 8925
rect 22646 8916 22652 8928
rect 22704 8916 22710 8968
rect 25133 8959 25191 8965
rect 25133 8925 25145 8959
rect 25179 8956 25191 8959
rect 25314 8956 25320 8968
rect 25179 8928 25320 8956
rect 25179 8925 25191 8928
rect 25133 8919 25191 8925
rect 25314 8916 25320 8928
rect 25372 8916 25378 8968
rect 27430 8916 27436 8968
rect 27488 8956 27494 8968
rect 28626 8956 28632 8968
rect 27488 8928 28632 8956
rect 27488 8916 27494 8928
rect 28626 8916 28632 8928
rect 28684 8916 28690 8968
rect 29822 8956 29828 8968
rect 29783 8928 29828 8956
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 20162 8848 20168 8900
rect 20220 8888 20226 8900
rect 20349 8891 20407 8897
rect 20349 8888 20361 8891
rect 20220 8860 20361 8888
rect 20220 8848 20226 8860
rect 20349 8857 20361 8860
rect 20395 8857 20407 8891
rect 20349 8851 20407 8857
rect 24489 8891 24547 8897
rect 24489 8857 24501 8891
rect 24535 8888 24547 8891
rect 26142 8888 26148 8900
rect 24535 8860 26148 8888
rect 24535 8857 24547 8860
rect 24489 8851 24547 8857
rect 26142 8848 26148 8860
rect 26200 8848 26206 8900
rect 27525 8891 27583 8897
rect 27525 8857 27537 8891
rect 27571 8888 27583 8891
rect 28721 8891 28779 8897
rect 27571 8860 28672 8888
rect 27571 8857 27583 8860
rect 27525 8851 27583 8857
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2130 8820 2136 8832
rect 2091 8792 2136 8820
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 23106 8780 23112 8832
rect 23164 8820 23170 8832
rect 24581 8823 24639 8829
rect 24581 8820 24593 8823
rect 23164 8792 24593 8820
rect 23164 8780 23170 8792
rect 24581 8789 24593 8792
rect 24627 8789 24639 8823
rect 24581 8783 24639 8789
rect 27246 8780 27252 8832
rect 27304 8820 27310 8832
rect 27433 8823 27491 8829
rect 27433 8820 27445 8823
rect 27304 8792 27445 8820
rect 27304 8780 27310 8792
rect 27433 8789 27445 8792
rect 27479 8789 27491 8823
rect 28258 8820 28264 8832
rect 28219 8792 28264 8820
rect 27433 8783 27491 8789
rect 28258 8780 28264 8792
rect 28316 8780 28322 8832
rect 28644 8820 28672 8860
rect 28721 8857 28733 8891
rect 28767 8888 28779 8891
rect 30374 8888 30380 8900
rect 28767 8860 30380 8888
rect 28767 8857 28779 8860
rect 28721 8851 28779 8857
rect 30374 8848 30380 8860
rect 30432 8848 30438 8900
rect 29362 8820 29368 8832
rect 28644 8792 29368 8820
rect 29362 8780 29368 8792
rect 29420 8780 29426 8832
rect 1104 8730 30820 8752
rect 1104 8678 10880 8730
rect 10932 8678 10944 8730
rect 10996 8678 11008 8730
rect 11060 8678 11072 8730
rect 11124 8678 11136 8730
rect 11188 8678 20811 8730
rect 20863 8678 20875 8730
rect 20927 8678 20939 8730
rect 20991 8678 21003 8730
rect 21055 8678 21067 8730
rect 21119 8678 30820 8730
rect 1104 8656 30820 8678
rect 24688 8588 26096 8616
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8480 1455 8483
rect 2130 8480 2136 8492
rect 1443 8452 2136 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 24026 8440 24032 8492
rect 24084 8480 24090 8492
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 24084 8452 24225 8480
rect 24084 8440 24090 8452
rect 24213 8449 24225 8452
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24489 8483 24547 8489
rect 24489 8449 24501 8483
rect 24535 8480 24547 8483
rect 24578 8480 24584 8492
rect 24535 8452 24584 8480
rect 24535 8449 24547 8452
rect 24489 8443 24547 8449
rect 24578 8440 24584 8452
rect 24636 8440 24642 8492
rect 24688 8489 24716 8588
rect 25409 8551 25467 8557
rect 25409 8517 25421 8551
rect 25455 8548 25467 8551
rect 25590 8548 25596 8560
rect 25455 8520 25596 8548
rect 25455 8517 25467 8520
rect 25409 8511 25467 8517
rect 25590 8508 25596 8520
rect 25648 8508 25654 8560
rect 26068 8548 26096 8588
rect 26142 8576 26148 8628
rect 26200 8616 26206 8628
rect 26329 8619 26387 8625
rect 26329 8616 26341 8619
rect 26200 8588 26341 8616
rect 26200 8576 26206 8588
rect 26329 8585 26341 8588
rect 26375 8585 26387 8619
rect 26329 8579 26387 8585
rect 27062 8576 27068 8628
rect 27120 8616 27126 8628
rect 27525 8619 27583 8625
rect 27525 8616 27537 8619
rect 27120 8588 27537 8616
rect 27120 8576 27126 8588
rect 27525 8585 27537 8588
rect 27571 8585 27583 8619
rect 27525 8579 27583 8585
rect 29089 8619 29147 8625
rect 29089 8585 29101 8619
rect 29135 8616 29147 8619
rect 29362 8616 29368 8628
rect 29135 8588 29368 8616
rect 29135 8585 29147 8588
rect 29089 8579 29147 8585
rect 29362 8576 29368 8588
rect 29420 8616 29426 8628
rect 30742 8616 30748 8628
rect 29420 8588 30748 8616
rect 29420 8576 29426 8588
rect 30742 8576 30748 8588
rect 30800 8576 30806 8628
rect 26510 8548 26516 8560
rect 26068 8520 26516 8548
rect 26510 8508 26516 8520
rect 26568 8508 26574 8560
rect 26602 8508 26608 8560
rect 26660 8548 26666 8560
rect 27341 8551 27399 8557
rect 27341 8548 27353 8551
rect 26660 8520 27353 8548
rect 26660 8508 26666 8520
rect 27341 8517 27353 8520
rect 27387 8517 27399 8551
rect 27341 8511 27399 8517
rect 24673 8483 24731 8489
rect 24673 8449 24685 8483
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 25038 8480 25044 8492
rect 24820 8452 25044 8480
rect 24820 8440 24826 8452
rect 25038 8440 25044 8452
rect 25096 8480 25102 8492
rect 25225 8483 25283 8489
rect 25225 8480 25237 8483
rect 25096 8452 25237 8480
rect 25096 8440 25102 8452
rect 25225 8449 25237 8452
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 26145 8483 26203 8489
rect 26145 8449 26157 8483
rect 26191 8480 26203 8483
rect 27062 8480 27068 8492
rect 26191 8452 27068 8480
rect 26191 8449 26203 8452
rect 26145 8443 26203 8449
rect 27062 8440 27068 8452
rect 27120 8440 27126 8492
rect 27356 8480 27384 8511
rect 27522 8480 27528 8492
rect 27356 8452 27528 8480
rect 27522 8440 27528 8452
rect 27580 8440 27586 8492
rect 29270 8440 29276 8492
rect 29328 8440 29334 8492
rect 25590 8372 25596 8424
rect 25648 8412 25654 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 25648 8384 25973 8412
rect 25648 8372 25654 8384
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 25961 8375 26019 8381
rect 26068 8384 28089 8412
rect 1578 8344 1584 8356
rect 1539 8316 1584 8344
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 14274 8304 14280 8356
rect 14332 8344 14338 8356
rect 26068 8344 26096 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 29178 8372 29184 8424
rect 29236 8372 29242 8424
rect 14332 8316 26096 8344
rect 14332 8304 14338 8316
rect 26418 8304 26424 8356
rect 26476 8344 26482 8356
rect 26973 8347 27031 8353
rect 26973 8344 26985 8347
rect 26476 8316 26985 8344
rect 26476 8304 26482 8316
rect 26973 8313 26985 8316
rect 27019 8313 27031 8347
rect 26973 8307 27031 8313
rect 24026 8276 24032 8288
rect 23987 8248 24032 8276
rect 24026 8236 24032 8248
rect 24084 8236 24090 8288
rect 27338 8276 27344 8288
rect 27251 8248 27344 8276
rect 27338 8236 27344 8248
rect 27396 8276 27402 8288
rect 27890 8276 27896 8288
rect 27396 8248 27896 8276
rect 27396 8236 27402 8248
rect 27890 8236 27896 8248
rect 27948 8236 27954 8288
rect 1104 8186 30820 8208
rect 1104 8134 5915 8186
rect 5967 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 15846 8186
rect 15898 8134 15910 8186
rect 15962 8134 15974 8186
rect 16026 8134 16038 8186
rect 16090 8134 16102 8186
rect 16154 8134 25776 8186
rect 25828 8134 25840 8186
rect 25892 8134 25904 8186
rect 25956 8134 25968 8186
rect 26020 8134 26032 8186
rect 26084 8134 30820 8186
rect 1104 8112 30820 8134
rect 23017 8075 23075 8081
rect 23017 8041 23029 8075
rect 23063 8072 23075 8075
rect 23106 8072 23112 8084
rect 23063 8044 23112 8072
rect 23063 8041 23075 8044
rect 23017 8035 23075 8041
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 2133 8007 2191 8013
rect 2133 7973 2145 8007
rect 2179 7973 2191 8007
rect 2133 7967 2191 7973
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 2148 7868 2176 7967
rect 27062 7964 27068 8016
rect 27120 7964 27126 8016
rect 24026 7936 24032 7948
rect 22848 7908 24032 7936
rect 1443 7840 2176 7868
rect 2317 7871 2375 7877
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2682 7868 2688 7880
rect 2363 7840 2688 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 22848 7877 22876 7908
rect 24026 7896 24032 7908
rect 24084 7896 24090 7948
rect 25498 7936 25504 7948
rect 25459 7908 25504 7936
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 26789 7939 26847 7945
rect 26789 7905 26801 7939
rect 26835 7936 26847 7939
rect 27080 7936 27108 7964
rect 26835 7908 27108 7936
rect 26835 7905 26847 7908
rect 26789 7899 26847 7905
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23382 7868 23388 7880
rect 23155 7840 23388 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 25682 7828 25688 7880
rect 25740 7868 25746 7880
rect 25777 7871 25835 7877
rect 25777 7868 25789 7871
rect 25740 7840 25789 7868
rect 25740 7828 25746 7840
rect 25777 7837 25789 7840
rect 25823 7837 25835 7871
rect 25777 7831 25835 7837
rect 26050 7828 26056 7880
rect 26108 7868 26114 7880
rect 27065 7871 27123 7877
rect 27065 7868 27077 7871
rect 26108 7840 27077 7868
rect 26108 7828 26114 7840
rect 27065 7837 27077 7840
rect 27111 7837 27123 7871
rect 28258 7868 28264 7880
rect 28219 7840 28264 7868
rect 27065 7831 27123 7837
rect 28258 7828 28264 7840
rect 28316 7828 28322 7880
rect 28718 7828 28724 7880
rect 28776 7868 28782 7880
rect 29917 7871 29975 7877
rect 29917 7868 29929 7871
rect 28776 7840 29929 7868
rect 28776 7828 28782 7840
rect 29917 7837 29929 7840
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 25958 7760 25964 7812
rect 26016 7800 26022 7812
rect 30101 7803 30159 7809
rect 30101 7800 30113 7803
rect 26016 7772 30113 7800
rect 26016 7760 26022 7772
rect 30101 7769 30113 7772
rect 30147 7769 30159 7803
rect 30101 7763 30159 7769
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 22646 7732 22652 7744
rect 22607 7704 22652 7732
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 25222 7692 25228 7744
rect 25280 7732 25286 7744
rect 26142 7732 26148 7744
rect 25280 7704 26148 7732
rect 25280 7692 25286 7704
rect 26142 7692 26148 7704
rect 26200 7692 26206 7744
rect 28350 7732 28356 7744
rect 28311 7704 28356 7732
rect 28350 7692 28356 7704
rect 28408 7692 28414 7744
rect 1104 7642 30820 7664
rect 1104 7590 10880 7642
rect 10932 7590 10944 7642
rect 10996 7590 11008 7642
rect 11060 7590 11072 7642
rect 11124 7590 11136 7642
rect 11188 7590 20811 7642
rect 20863 7590 20875 7642
rect 20927 7590 20939 7642
rect 20991 7590 21003 7642
rect 21055 7590 21067 7642
rect 21119 7590 30820 7642
rect 1104 7568 30820 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 28350 7528 28356 7540
rect 2096 7500 28356 7528
rect 2096 7488 2102 7500
rect 28350 7488 28356 7500
rect 28408 7488 28414 7540
rect 29086 7528 29092 7540
rect 28999 7500 29092 7528
rect 29086 7488 29092 7500
rect 29144 7528 29150 7540
rect 30466 7528 30472 7540
rect 29144 7500 30472 7528
rect 29144 7488 29150 7500
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 28077 7463 28135 7469
rect 28077 7460 28089 7463
rect 6420 7432 28089 7460
rect 6420 7420 6426 7432
rect 28077 7429 28089 7432
rect 28123 7429 28135 7463
rect 28077 7423 28135 7429
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 24305 7395 24363 7401
rect 1443 7364 6914 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 6886 7256 6914 7364
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24486 7392 24492 7404
rect 24447 7364 24492 7392
rect 24305 7355 24363 7361
rect 24320 7324 24348 7355
rect 24486 7352 24492 7364
rect 24544 7352 24550 7404
rect 24578 7352 24584 7404
rect 24636 7392 24642 7404
rect 24636 7364 24681 7392
rect 24636 7352 24642 7364
rect 25682 7352 25688 7404
rect 25740 7392 25746 7404
rect 26329 7395 26387 7401
rect 26329 7392 26341 7395
rect 25740 7364 26341 7392
rect 25740 7352 25746 7364
rect 26329 7361 26341 7364
rect 26375 7361 26387 7395
rect 26970 7392 26976 7404
rect 26931 7364 26976 7392
rect 26329 7355 26387 7361
rect 26970 7352 26976 7364
rect 27028 7352 27034 7404
rect 28994 7352 29000 7404
rect 29052 7352 29058 7404
rect 25406 7324 25412 7336
rect 24320 7296 25412 7324
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 25498 7284 25504 7336
rect 25556 7324 25562 7336
rect 26050 7324 26056 7336
rect 25556 7296 26056 7324
rect 25556 7284 25562 7296
rect 26050 7284 26056 7296
rect 26108 7284 26114 7336
rect 26145 7327 26203 7333
rect 26145 7293 26157 7327
rect 26191 7293 26203 7327
rect 26145 7287 26203 7293
rect 26237 7327 26295 7333
rect 26237 7293 26249 7327
rect 26283 7324 26295 7327
rect 26786 7324 26792 7336
rect 26283 7296 26792 7324
rect 26283 7293 26295 7296
rect 26237 7287 26295 7293
rect 25958 7256 25964 7268
rect 6886 7228 25964 7256
rect 25958 7216 25964 7228
rect 26016 7216 26022 7268
rect 26160 7200 26188 7287
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 29178 7284 29184 7336
rect 29236 7284 29242 7336
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 24118 7188 24124 7200
rect 24079 7160 24124 7188
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 25222 7148 25228 7200
rect 25280 7188 25286 7200
rect 25869 7191 25927 7197
rect 25869 7188 25881 7191
rect 25280 7160 25881 7188
rect 25280 7148 25286 7160
rect 25869 7157 25881 7160
rect 25915 7157 25927 7191
rect 25869 7151 25927 7157
rect 26142 7148 26148 7200
rect 26200 7188 26206 7200
rect 27157 7191 27215 7197
rect 27157 7188 27169 7191
rect 26200 7160 27169 7188
rect 26200 7148 26206 7160
rect 27157 7157 27169 7160
rect 27203 7157 27215 7191
rect 27157 7151 27215 7157
rect 1104 7098 30820 7120
rect 1104 7046 5915 7098
rect 5967 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 15846 7098
rect 15898 7046 15910 7098
rect 15962 7046 15974 7098
rect 16026 7046 16038 7098
rect 16090 7046 16102 7098
rect 16154 7046 25776 7098
rect 25828 7046 25840 7098
rect 25892 7046 25904 7098
rect 25956 7046 25968 7098
rect 26020 7046 26032 7098
rect 26084 7046 30820 7098
rect 1104 7024 30820 7046
rect 22925 6987 22983 6993
rect 22925 6953 22937 6987
rect 22971 6984 22983 6987
rect 23382 6984 23388 6996
rect 22971 6956 23388 6984
rect 22971 6953 22983 6956
rect 22925 6947 22983 6953
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 28534 6944 28540 6996
rect 28592 6984 28598 6996
rect 30009 6987 30067 6993
rect 30009 6984 30021 6987
rect 28592 6956 30021 6984
rect 28592 6944 28598 6956
rect 30009 6953 30021 6956
rect 30055 6953 30067 6987
rect 30009 6947 30067 6953
rect 25590 6876 25596 6928
rect 25648 6916 25654 6928
rect 26142 6916 26148 6928
rect 25648 6888 26148 6916
rect 25648 6876 25654 6888
rect 26142 6876 26148 6888
rect 26200 6916 26206 6928
rect 26970 6916 26976 6928
rect 26200 6888 26976 6916
rect 26200 6876 26206 6888
rect 26970 6876 26976 6888
rect 27028 6876 27034 6928
rect 25406 6848 25412 6860
rect 25367 6820 25412 6848
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 25608 6848 25636 6876
rect 25685 6851 25743 6857
rect 25685 6848 25697 6851
rect 25608 6820 25697 6848
rect 25685 6817 25697 6820
rect 25731 6817 25743 6851
rect 25685 6811 25743 6817
rect 25777 6851 25835 6857
rect 25777 6817 25789 6851
rect 25823 6848 25835 6851
rect 27706 6848 27712 6860
rect 25823 6820 26924 6848
rect 25823 6817 25835 6820
rect 25777 6811 25835 6817
rect 21542 6780 21548 6792
rect 21455 6752 21548 6780
rect 21542 6740 21548 6752
rect 21600 6780 21606 6792
rect 21600 6752 22048 6780
rect 21600 6740 21606 6752
rect 22020 6724 22048 6752
rect 25498 6740 25504 6792
rect 25556 6780 25562 6792
rect 25593 6783 25651 6789
rect 25593 6780 25605 6783
rect 25556 6752 25605 6780
rect 25556 6740 25562 6752
rect 25593 6749 25605 6752
rect 25639 6749 25651 6783
rect 25593 6743 25651 6749
rect 25869 6783 25927 6789
rect 25869 6749 25881 6783
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 21812 6715 21870 6721
rect 21812 6681 21824 6715
rect 21858 6712 21870 6715
rect 21858 6684 21956 6712
rect 21858 6681 21870 6684
rect 21812 6675 21870 6681
rect 21928 6644 21956 6684
rect 22002 6672 22008 6724
rect 22060 6672 22066 6724
rect 25884 6712 25912 6743
rect 25700 6684 25912 6712
rect 26896 6712 26924 6820
rect 26988 6820 27712 6848
rect 26988 6789 27016 6820
rect 27706 6808 27712 6820
rect 27764 6808 27770 6860
rect 28718 6848 28724 6860
rect 28679 6820 28724 6848
rect 28718 6808 28724 6820
rect 28776 6808 28782 6860
rect 30190 6848 30196 6860
rect 28828 6820 30196 6848
rect 26973 6783 27031 6789
rect 26973 6749 26985 6783
rect 27019 6749 27031 6783
rect 27614 6780 27620 6792
rect 27575 6752 27620 6780
rect 26973 6743 27031 6749
rect 27614 6740 27620 6752
rect 27672 6740 27678 6792
rect 28828 6780 28856 6820
rect 30190 6808 30196 6820
rect 30248 6808 30254 6860
rect 28368 6752 28856 6780
rect 28368 6712 28396 6752
rect 28902 6740 28908 6792
rect 28960 6780 28966 6792
rect 29825 6783 29883 6789
rect 29825 6780 29837 6783
rect 28960 6752 29837 6780
rect 28960 6740 28966 6752
rect 29825 6749 29837 6752
rect 29871 6749 29883 6783
rect 29825 6743 29883 6749
rect 26896 6684 28396 6712
rect 28445 6715 28503 6721
rect 25700 6656 25728 6684
rect 28445 6681 28457 6715
rect 28491 6712 28503 6715
rect 28994 6712 29000 6724
rect 28491 6684 29000 6712
rect 28491 6681 28503 6684
rect 28445 6675 28503 6681
rect 28994 6672 29000 6684
rect 29052 6672 29058 6724
rect 22646 6644 22652 6656
rect 21928 6616 22652 6644
rect 22646 6604 22652 6616
rect 22704 6604 22710 6656
rect 25682 6604 25688 6656
rect 25740 6604 25746 6656
rect 26789 6647 26847 6653
rect 26789 6613 26801 6647
rect 26835 6644 26847 6647
rect 27246 6644 27252 6656
rect 26835 6616 27252 6644
rect 26835 6613 26847 6616
rect 26789 6607 26847 6613
rect 27246 6604 27252 6616
rect 27304 6604 27310 6656
rect 27430 6644 27436 6656
rect 27391 6616 27436 6644
rect 27430 6604 27436 6616
rect 27488 6604 27494 6656
rect 28074 6644 28080 6656
rect 28035 6616 28080 6644
rect 28074 6604 28080 6616
rect 28132 6604 28138 6656
rect 28537 6647 28595 6653
rect 28537 6613 28549 6647
rect 28583 6644 28595 6647
rect 29086 6644 29092 6656
rect 28583 6616 29092 6644
rect 28583 6613 28595 6616
rect 28537 6607 28595 6613
rect 29086 6604 29092 6616
rect 29144 6604 29150 6656
rect 1104 6554 30820 6576
rect 1104 6502 10880 6554
rect 10932 6502 10944 6554
rect 10996 6502 11008 6554
rect 11060 6502 11072 6554
rect 11124 6502 11136 6554
rect 11188 6502 20811 6554
rect 20863 6502 20875 6554
rect 20927 6502 20939 6554
rect 20991 6502 21003 6554
rect 21055 6502 21067 6554
rect 21119 6502 30820 6554
rect 1104 6480 30820 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 24486 6400 24492 6452
rect 24544 6440 24550 6452
rect 24673 6443 24731 6449
rect 24673 6440 24685 6443
rect 24544 6412 24685 6440
rect 24544 6400 24550 6412
rect 24673 6409 24685 6412
rect 24719 6409 24731 6443
rect 24673 6403 24731 6409
rect 28537 6443 28595 6449
rect 28537 6409 28549 6443
rect 28583 6440 28595 6443
rect 29270 6440 29276 6452
rect 28583 6412 29276 6440
rect 28583 6409 28595 6412
rect 28537 6403 28595 6409
rect 29270 6400 29276 6412
rect 29328 6400 29334 6452
rect 29822 6440 29828 6452
rect 29783 6412 29828 6440
rect 29822 6400 29828 6412
rect 29880 6400 29886 6452
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 2056 6304 2084 6400
rect 23560 6375 23618 6381
rect 23560 6341 23572 6375
rect 23606 6372 23618 6375
rect 24118 6372 24124 6384
rect 23606 6344 24124 6372
rect 23606 6341 23618 6344
rect 23560 6335 23618 6341
rect 24118 6332 24124 6344
rect 24176 6332 24182 6384
rect 27433 6375 27491 6381
rect 27433 6341 27445 6375
rect 27479 6372 27491 6375
rect 28074 6372 28080 6384
rect 27479 6344 28080 6372
rect 27479 6341 27491 6344
rect 27433 6335 27491 6341
rect 28074 6332 28080 6344
rect 28132 6332 28138 6384
rect 28629 6375 28687 6381
rect 28629 6341 28641 6375
rect 28675 6372 28687 6375
rect 29362 6372 29368 6384
rect 28675 6344 29368 6372
rect 28675 6341 28687 6344
rect 28629 6335 28687 6341
rect 29362 6332 29368 6344
rect 29420 6332 29426 6384
rect 1443 6276 2084 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 29086 6264 29092 6316
rect 29144 6304 29150 6316
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 29144 6276 29745 6304
rect 29144 6264 29150 6276
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 22002 6196 22008 6248
rect 22060 6236 22066 6248
rect 23293 6239 23351 6245
rect 23293 6236 23305 6239
rect 22060 6208 23305 6236
rect 22060 6196 22066 6208
rect 23293 6205 23305 6208
rect 23339 6205 23351 6239
rect 23293 6199 23351 6205
rect 28718 6196 28724 6248
rect 28776 6236 28782 6248
rect 28813 6239 28871 6245
rect 28813 6236 28825 6239
rect 28776 6208 28825 6236
rect 28776 6196 28782 6208
rect 28813 6205 28825 6208
rect 28859 6236 28871 6239
rect 29917 6239 29975 6245
rect 29917 6236 29929 6239
rect 28859 6208 29929 6236
rect 28859 6205 28871 6208
rect 28813 6199 28871 6205
rect 29917 6205 29929 6208
rect 29963 6205 29975 6239
rect 29917 6199 29975 6205
rect 1578 6168 1584 6180
rect 1539 6140 1584 6168
rect 1578 6128 1584 6140
rect 1636 6128 1642 6180
rect 24762 6060 24768 6112
rect 24820 6100 24826 6112
rect 27525 6103 27583 6109
rect 27525 6100 27537 6103
rect 24820 6072 27537 6100
rect 24820 6060 24826 6072
rect 27525 6069 27537 6072
rect 27571 6069 27583 6103
rect 27525 6063 27583 6069
rect 27982 6060 27988 6112
rect 28040 6100 28046 6112
rect 28169 6103 28227 6109
rect 28169 6100 28181 6103
rect 28040 6072 28181 6100
rect 28040 6060 28046 6072
rect 28169 6069 28181 6072
rect 28215 6069 28227 6103
rect 29362 6100 29368 6112
rect 29323 6072 29368 6100
rect 28169 6063 28227 6069
rect 29362 6060 29368 6072
rect 29420 6060 29426 6112
rect 1104 6010 30820 6032
rect 1104 5958 5915 6010
rect 5967 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 15846 6010
rect 15898 5958 15910 6010
rect 15962 5958 15974 6010
rect 16026 5958 16038 6010
rect 16090 5958 16102 6010
rect 16154 5958 25776 6010
rect 25828 5958 25840 6010
rect 25892 5958 25904 6010
rect 25956 5958 25968 6010
rect 26020 5958 26032 6010
rect 26084 5958 30820 6010
rect 1104 5936 30820 5958
rect 28077 5899 28135 5905
rect 28077 5896 28089 5899
rect 6886 5868 28089 5896
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 6886 5760 6914 5868
rect 28077 5865 28089 5868
rect 28123 5865 28135 5899
rect 28077 5859 28135 5865
rect 28813 5899 28871 5905
rect 28813 5865 28825 5899
rect 28859 5896 28871 5899
rect 28994 5896 29000 5908
rect 28859 5868 29000 5896
rect 28859 5865 28871 5868
rect 28813 5859 28871 5865
rect 28994 5856 29000 5868
rect 29052 5856 29058 5908
rect 29270 5856 29276 5908
rect 29328 5896 29334 5908
rect 29917 5899 29975 5905
rect 29917 5896 29929 5899
rect 29328 5868 29929 5896
rect 29328 5856 29334 5868
rect 29917 5865 29929 5868
rect 29963 5865 29975 5899
rect 29917 5859 29975 5865
rect 25590 5760 25596 5772
rect 2740 5732 6914 5760
rect 25503 5732 25596 5760
rect 2740 5720 2746 5732
rect 25590 5720 25596 5732
rect 25648 5760 25654 5772
rect 26142 5760 26148 5772
rect 25648 5732 26148 5760
rect 25648 5720 25654 5732
rect 26142 5720 26148 5732
rect 26200 5760 26206 5772
rect 26881 5763 26939 5769
rect 26881 5760 26893 5763
rect 26200 5732 26893 5760
rect 26200 5720 26206 5732
rect 26881 5729 26893 5732
rect 26927 5729 26939 5763
rect 26881 5723 26939 5729
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 25498 5692 25504 5704
rect 1443 5664 6914 5692
rect 25459 5664 25504 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 6886 5624 6914 5664
rect 25498 5652 25504 5664
rect 25556 5652 25562 5704
rect 25685 5695 25743 5701
rect 25685 5661 25697 5695
rect 25731 5661 25743 5695
rect 25685 5655 25743 5661
rect 24762 5624 24768 5636
rect 6886 5596 24768 5624
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 25314 5556 25320 5568
rect 25275 5528 25320 5556
rect 25314 5516 25320 5528
rect 25372 5516 25378 5568
rect 25700 5556 25728 5655
rect 25774 5652 25780 5704
rect 25832 5692 25838 5704
rect 26602 5692 26608 5704
rect 25832 5664 25877 5692
rect 26563 5664 26608 5692
rect 25832 5652 25838 5664
rect 26602 5652 26608 5664
rect 26660 5652 26666 5704
rect 27982 5692 27988 5704
rect 27943 5664 27988 5692
rect 27982 5652 27988 5664
rect 28040 5652 28046 5704
rect 28810 5652 28816 5704
rect 28868 5692 28874 5704
rect 28997 5695 29055 5701
rect 28997 5692 29009 5695
rect 28868 5664 29009 5692
rect 28868 5652 28874 5664
rect 28997 5661 29009 5664
rect 29043 5661 29055 5695
rect 30098 5692 30104 5704
rect 30059 5664 30104 5692
rect 28997 5655 29055 5661
rect 30098 5652 30104 5664
rect 30156 5652 30162 5704
rect 27154 5556 27160 5568
rect 25700 5528 27160 5556
rect 27154 5516 27160 5528
rect 27212 5516 27218 5568
rect 1104 5466 30820 5488
rect 1104 5414 10880 5466
rect 10932 5414 10944 5466
rect 10996 5414 11008 5466
rect 11060 5414 11072 5466
rect 11124 5414 11136 5466
rect 11188 5414 20811 5466
rect 20863 5414 20875 5466
rect 20927 5414 20939 5466
rect 20991 5414 21003 5466
rect 21055 5414 21067 5466
rect 21119 5414 30820 5466
rect 1104 5392 30820 5414
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 23293 5355 23351 5361
rect 23293 5352 23305 5355
rect 22336 5324 23305 5352
rect 22336 5312 22342 5324
rect 23293 5321 23305 5324
rect 23339 5321 23351 5355
rect 23293 5315 23351 5321
rect 23934 5312 23940 5364
rect 23992 5352 23998 5364
rect 27985 5355 28043 5361
rect 23992 5324 27936 5352
rect 23992 5312 23998 5324
rect 22186 5244 22192 5296
rect 22244 5284 22250 5296
rect 24397 5287 24455 5293
rect 24397 5284 24409 5287
rect 22244 5256 24409 5284
rect 22244 5244 22250 5256
rect 24397 5253 24409 5256
rect 24443 5284 24455 5287
rect 24670 5284 24676 5296
rect 24443 5256 24676 5284
rect 24443 5253 24455 5256
rect 24397 5247 24455 5253
rect 24670 5244 24676 5256
rect 24728 5244 24734 5296
rect 25498 5244 25504 5296
rect 25556 5284 25562 5296
rect 27157 5287 27215 5293
rect 27157 5284 27169 5287
rect 25556 5256 27169 5284
rect 25556 5244 25562 5256
rect 27157 5253 27169 5256
rect 27203 5253 27215 5287
rect 27908 5284 27936 5324
rect 27985 5321 27997 5355
rect 28031 5352 28043 5355
rect 29086 5352 29092 5364
rect 28031 5324 29092 5352
rect 28031 5321 28043 5324
rect 27985 5315 28043 5321
rect 29086 5312 29092 5324
rect 29144 5312 29150 5364
rect 29822 5352 29828 5364
rect 29783 5324 29828 5352
rect 29822 5312 29828 5324
rect 29880 5312 29886 5364
rect 28721 5287 28779 5293
rect 27908 5256 28672 5284
rect 27157 5247 27215 5253
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 2682 5216 2688 5228
rect 1443 5188 2688 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 23198 5216 23204 5228
rect 23159 5188 23204 5216
rect 23198 5176 23204 5188
rect 23256 5176 23262 5228
rect 24213 5219 24271 5225
rect 24213 5185 24225 5219
rect 24259 5185 24271 5219
rect 24213 5179 24271 5185
rect 24489 5219 24547 5225
rect 24489 5185 24501 5219
rect 24535 5216 24547 5219
rect 24578 5216 24584 5228
rect 24535 5188 24584 5216
rect 24535 5185 24547 5188
rect 24489 5179 24547 5185
rect 24228 5148 24256 5179
rect 24578 5176 24584 5188
rect 24636 5176 24642 5228
rect 25590 5216 25596 5228
rect 25551 5188 25596 5216
rect 25590 5176 25596 5188
rect 25648 5176 25654 5228
rect 26973 5219 27031 5225
rect 26973 5185 26985 5219
rect 27019 5216 27031 5219
rect 27062 5216 27068 5228
rect 27019 5188 27068 5216
rect 27019 5185 27031 5188
rect 26973 5179 27031 5185
rect 27062 5176 27068 5188
rect 27120 5216 27126 5228
rect 27617 5219 27675 5225
rect 27617 5216 27629 5219
rect 27120 5188 27629 5216
rect 27120 5176 27126 5188
rect 27617 5185 27629 5188
rect 27663 5185 27675 5219
rect 28166 5216 28172 5228
rect 28127 5188 28172 5216
rect 27617 5179 27675 5185
rect 28166 5176 28172 5188
rect 28224 5176 28230 5228
rect 28644 5216 28672 5256
rect 28721 5253 28733 5287
rect 28767 5284 28779 5287
rect 29362 5284 29368 5296
rect 28767 5256 29368 5284
rect 28767 5253 28779 5256
rect 28721 5247 28779 5253
rect 29362 5244 29368 5256
rect 29420 5244 29426 5296
rect 28994 5216 29000 5228
rect 28644 5188 29000 5216
rect 28994 5176 29000 5188
rect 29052 5176 29058 5228
rect 29086 5176 29092 5228
rect 29144 5216 29150 5228
rect 29733 5219 29791 5225
rect 29733 5216 29745 5219
rect 29144 5188 29745 5216
rect 29144 5176 29150 5188
rect 29733 5185 29745 5188
rect 29779 5185 29791 5219
rect 29733 5179 29791 5185
rect 25317 5151 25375 5157
rect 25317 5148 25329 5151
rect 24228 5120 25329 5148
rect 25317 5117 25329 5120
rect 25363 5117 25375 5151
rect 25498 5148 25504 5160
rect 25459 5120 25504 5148
rect 25317 5111 25375 5117
rect 25498 5108 25504 5120
rect 25556 5108 25562 5160
rect 25685 5151 25743 5157
rect 25685 5117 25697 5151
rect 25731 5117 25743 5151
rect 25685 5111 25743 5117
rect 24946 5040 24952 5092
rect 25004 5080 25010 5092
rect 25700 5080 25728 5111
rect 25774 5108 25780 5160
rect 25832 5148 25838 5160
rect 26142 5148 26148 5160
rect 25832 5120 26148 5148
rect 25832 5108 25838 5120
rect 26142 5108 26148 5120
rect 26200 5108 26206 5160
rect 29012 5148 29040 5176
rect 29914 5148 29920 5160
rect 29012 5120 29920 5148
rect 29914 5108 29920 5120
rect 29972 5108 29978 5160
rect 25004 5052 25728 5080
rect 25004 5040 25010 5052
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 24026 5012 24032 5024
rect 23987 4984 24032 5012
rect 24026 4972 24032 4984
rect 24084 4972 24090 5024
rect 27341 5015 27399 5021
rect 27341 4981 27353 5015
rect 27387 5012 27399 5015
rect 27430 5012 27436 5024
rect 27387 4984 27436 5012
rect 27387 4981 27399 4984
rect 27341 4975 27399 4981
rect 27430 4972 27436 4984
rect 27488 4972 27494 5024
rect 27706 4972 27712 5024
rect 27764 5012 27770 5024
rect 28813 5015 28871 5021
rect 28813 5012 28825 5015
rect 27764 4984 28825 5012
rect 27764 4972 27770 4984
rect 28813 4981 28825 4984
rect 28859 4981 28871 5015
rect 29362 5012 29368 5024
rect 29323 4984 29368 5012
rect 28813 4975 28871 4981
rect 29362 4972 29368 4984
rect 29420 4972 29426 5024
rect 1104 4922 30820 4944
rect 1104 4870 5915 4922
rect 5967 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 15846 4922
rect 15898 4870 15910 4922
rect 15962 4870 15974 4922
rect 16026 4870 16038 4922
rect 16090 4870 16102 4922
rect 16154 4870 25776 4922
rect 25828 4870 25840 4922
rect 25892 4870 25904 4922
rect 25956 4870 25968 4922
rect 26020 4870 26032 4922
rect 26084 4870 30820 4922
rect 1104 4848 30820 4870
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 26973 4811 27031 4817
rect 26973 4808 26985 4811
rect 23256 4780 26985 4808
rect 23256 4768 23262 4780
rect 26973 4777 26985 4780
rect 27019 4777 27031 4811
rect 26973 4771 27031 4777
rect 24578 4700 24584 4752
rect 24636 4740 24642 4752
rect 26878 4740 26884 4752
rect 24636 4712 25544 4740
rect 26839 4712 26884 4740
rect 24636 4700 24642 4712
rect 25314 4672 25320 4684
rect 23584 4644 25320 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1443 4576 6914 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 6886 4536 6914 4576
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23474 4604 23480 4616
rect 23072 4576 23480 4604
rect 23072 4564 23078 4576
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 23584 4613 23612 4644
rect 25314 4632 25320 4644
rect 25372 4632 25378 4684
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 23845 4607 23903 4613
rect 23845 4573 23857 4607
rect 23891 4604 23903 4607
rect 24578 4604 24584 4616
rect 23891 4576 24584 4604
rect 23891 4573 23903 4576
rect 23845 4567 23903 4573
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 25222 4604 25228 4616
rect 25183 4576 25228 4604
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 25406 4604 25412 4616
rect 25367 4576 25412 4604
rect 25406 4564 25412 4576
rect 25464 4564 25470 4616
rect 25516 4613 25544 4712
rect 26878 4700 26884 4712
rect 26936 4700 26942 4752
rect 28261 4743 28319 4749
rect 28261 4709 28273 4743
rect 28307 4709 28319 4743
rect 28261 4703 28319 4709
rect 26142 4632 26148 4684
rect 26200 4672 26206 4684
rect 26513 4675 26571 4681
rect 26513 4672 26525 4675
rect 26200 4644 26525 4672
rect 26200 4632 26206 4644
rect 26513 4641 26525 4644
rect 26559 4641 26571 4675
rect 27706 4672 27712 4684
rect 26513 4635 26571 4641
rect 26620 4644 27712 4672
rect 25501 4607 25559 4613
rect 25501 4573 25513 4607
rect 25547 4573 25559 4607
rect 25501 4567 25559 4573
rect 26620 4536 26648 4644
rect 27706 4632 27712 4644
rect 27764 4632 27770 4684
rect 27798 4604 27804 4616
rect 27759 4576 27804 4604
rect 27798 4564 27804 4576
rect 27856 4564 27862 4616
rect 28276 4604 28304 4703
rect 28718 4672 28724 4684
rect 28679 4644 28724 4672
rect 28718 4632 28724 4644
rect 28776 4632 28782 4684
rect 28905 4675 28963 4681
rect 28905 4641 28917 4675
rect 28951 4672 28963 4675
rect 28994 4672 29000 4684
rect 28951 4644 29000 4672
rect 28951 4641 28963 4644
rect 28905 4635 28963 4641
rect 28994 4632 29000 4644
rect 29052 4632 29058 4684
rect 29917 4607 29975 4613
rect 29917 4604 29929 4607
rect 28276 4576 29929 4604
rect 29917 4573 29929 4576
rect 29963 4573 29975 4607
rect 29917 4567 29975 4573
rect 28629 4539 28687 4545
rect 28629 4536 28641 4539
rect 6886 4508 26648 4536
rect 27632 4508 28641 4536
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 23382 4468 23388 4480
rect 23343 4440 23388 4468
rect 23382 4428 23388 4440
rect 23440 4428 23446 4480
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 23753 4471 23811 4477
rect 23753 4468 23765 4471
rect 23532 4440 23765 4468
rect 23532 4428 23538 4440
rect 23753 4437 23765 4440
rect 23799 4437 23811 4471
rect 23753 4431 23811 4437
rect 25041 4471 25099 4477
rect 25041 4437 25053 4471
rect 25087 4468 25099 4471
rect 25130 4468 25136 4480
rect 25087 4440 25136 4468
rect 25087 4437 25099 4440
rect 25041 4431 25099 4437
rect 25130 4428 25136 4440
rect 25188 4428 25194 4480
rect 27632 4477 27660 4508
rect 28629 4505 28641 4508
rect 28675 4505 28687 4539
rect 28629 4499 28687 4505
rect 27617 4471 27675 4477
rect 27617 4437 27629 4471
rect 27663 4437 27675 4471
rect 27617 4431 27675 4437
rect 27706 4428 27712 4480
rect 27764 4468 27770 4480
rect 30009 4471 30067 4477
rect 30009 4468 30021 4471
rect 27764 4440 30021 4468
rect 27764 4428 27770 4440
rect 30009 4437 30021 4440
rect 30055 4437 30067 4471
rect 30009 4431 30067 4437
rect 1104 4378 30820 4400
rect 1104 4326 10880 4378
rect 10932 4326 10944 4378
rect 10996 4326 11008 4378
rect 11060 4326 11072 4378
rect 11124 4326 11136 4378
rect 11188 4326 20811 4378
rect 20863 4326 20875 4378
rect 20927 4326 20939 4378
rect 20991 4326 21003 4378
rect 21055 4326 21067 4378
rect 21119 4326 30820 4378
rect 1104 4304 30820 4326
rect 2041 4267 2099 4273
rect 2041 4233 2053 4267
rect 2087 4264 2099 4267
rect 27706 4264 27712 4276
rect 2087 4236 27712 4264
rect 2087 4233 2099 4236
rect 2041 4227 2099 4233
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 2056 4128 2084 4227
rect 27706 4224 27712 4236
rect 27764 4224 27770 4276
rect 29365 4267 29423 4273
rect 29365 4233 29377 4267
rect 29411 4233 29423 4267
rect 29365 4227 29423 4233
rect 22272 4199 22330 4205
rect 22272 4165 22284 4199
rect 22318 4196 22330 4199
rect 23382 4196 23388 4208
rect 22318 4168 23388 4196
rect 22318 4165 22330 4168
rect 22272 4159 22330 4165
rect 23382 4156 23388 4168
rect 23440 4156 23446 4208
rect 24026 4156 24032 4208
rect 24084 4196 24090 4208
rect 24182 4199 24240 4205
rect 24182 4196 24194 4199
rect 24084 4168 24194 4196
rect 24084 4156 24090 4168
rect 24182 4165 24194 4168
rect 24228 4165 24240 4199
rect 24182 4159 24240 4165
rect 28537 4199 28595 4205
rect 28537 4165 28549 4199
rect 28583 4196 28595 4199
rect 29380 4196 29408 4227
rect 28583 4168 29408 4196
rect 28583 4165 28595 4168
rect 28537 4159 28595 4165
rect 16666 4128 16672 4140
rect 1443 4100 2084 4128
rect 16627 4100 16672 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 27430 4128 27436 4140
rect 27391 4100 27436 4128
rect 27430 4088 27436 4100
rect 27488 4088 27494 4140
rect 28166 4128 28172 4140
rect 28127 4100 28172 4128
rect 28166 4088 28172 4100
rect 28224 4088 28230 4140
rect 29730 4128 29736 4140
rect 29691 4100 29736 4128
rect 29730 4088 29736 4100
rect 29788 4088 29794 4140
rect 22002 4060 22008 4072
rect 21915 4032 22008 4060
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 23934 4060 23940 4072
rect 23308 4032 23940 4060
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 22020 3924 22048 4020
rect 23308 3924 23336 4032
rect 23934 4020 23940 4032
rect 23992 4020 23998 4072
rect 28997 4063 29055 4069
rect 28997 4029 29009 4063
rect 29043 4060 29055 4063
rect 29822 4060 29828 4072
rect 29043 4032 29828 4060
rect 29043 4029 29055 4032
rect 28997 4023 29055 4029
rect 29822 4020 29828 4032
rect 29880 4020 29886 4072
rect 29914 4020 29920 4072
rect 29972 4060 29978 4072
rect 29972 4032 30017 4060
rect 29972 4020 29978 4032
rect 23382 3952 23388 4004
rect 23440 3992 23446 4004
rect 27985 3995 28043 4001
rect 23440 3964 23485 3992
rect 23440 3952 23446 3964
rect 27985 3961 27997 3995
rect 28031 3992 28043 3995
rect 29086 3992 29092 4004
rect 28031 3964 29092 3992
rect 28031 3961 28043 3964
rect 27985 3955 28043 3961
rect 29086 3952 29092 3964
rect 29144 3952 29150 4004
rect 22020 3896 23336 3924
rect 24670 3884 24676 3936
rect 24728 3924 24734 3936
rect 25317 3927 25375 3933
rect 25317 3924 25329 3927
rect 24728 3896 25329 3924
rect 24728 3884 24734 3896
rect 25317 3893 25329 3896
rect 25363 3893 25375 3927
rect 27246 3924 27252 3936
rect 27207 3896 27252 3924
rect 25317 3887 25375 3893
rect 27246 3884 27252 3896
rect 27304 3884 27310 3936
rect 28626 3924 28632 3936
rect 28587 3896 28632 3924
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 1104 3834 30820 3856
rect 1104 3782 5915 3834
rect 5967 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 15846 3834
rect 15898 3782 15910 3834
rect 15962 3782 15974 3834
rect 16026 3782 16038 3834
rect 16090 3782 16102 3834
rect 16154 3782 25776 3834
rect 25828 3782 25840 3834
rect 25892 3782 25904 3834
rect 25956 3782 25968 3834
rect 26020 3782 26032 3834
rect 26084 3782 30820 3834
rect 1104 3760 30820 3782
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 28626 3720 28632 3732
rect 2188 3692 28632 3720
rect 2188 3680 2194 3692
rect 28626 3680 28632 3692
rect 28684 3680 28690 3732
rect 28077 3655 28135 3661
rect 28077 3621 28089 3655
rect 28123 3652 28135 3655
rect 29730 3652 29736 3664
rect 28123 3624 29736 3652
rect 28123 3621 28135 3624
rect 28077 3615 28135 3621
rect 29730 3612 29736 3624
rect 29788 3612 29794 3664
rect 23934 3544 23940 3596
rect 23992 3584 23998 3596
rect 24857 3587 24915 3593
rect 24857 3584 24869 3587
rect 23992 3556 24869 3584
rect 23992 3544 23998 3556
rect 24857 3553 24869 3556
rect 24903 3553 24915 3587
rect 24857 3547 24915 3553
rect 27246 3544 27252 3596
rect 27304 3584 27310 3596
rect 27304 3556 28764 3584
rect 27304 3544 27310 3556
rect 25130 3525 25136 3528
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3516 1455 3519
rect 25124 3516 25136 3525
rect 1443 3488 6914 3516
rect 25091 3488 25136 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 6886 3448 6914 3488
rect 25124 3479 25136 3488
rect 25130 3476 25136 3479
rect 25188 3476 25194 3528
rect 28258 3516 28264 3528
rect 28219 3488 28264 3516
rect 28258 3476 28264 3488
rect 28316 3476 28322 3528
rect 28736 3525 28764 3556
rect 28721 3519 28779 3525
rect 28721 3485 28733 3519
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 29362 3476 29368 3528
rect 29420 3516 29426 3528
rect 29917 3519 29975 3525
rect 29917 3516 29929 3519
rect 29420 3488 29929 3516
rect 29420 3476 29426 3488
rect 29917 3485 29929 3488
rect 29963 3485 29975 3519
rect 29917 3479 29975 3485
rect 6886 3420 29040 3448
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 25406 3340 25412 3392
rect 25464 3380 25470 3392
rect 26237 3383 26295 3389
rect 26237 3380 26249 3383
rect 25464 3352 26249 3380
rect 25464 3340 25470 3352
rect 26237 3349 26249 3352
rect 26283 3349 26295 3383
rect 28902 3380 28908 3392
rect 28863 3352 28908 3380
rect 26237 3343 26295 3349
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 29012 3380 29040 3420
rect 30009 3383 30067 3389
rect 30009 3380 30021 3383
rect 29012 3352 30021 3380
rect 30009 3349 30021 3352
rect 30055 3349 30067 3383
rect 30009 3343 30067 3349
rect 1104 3290 30820 3312
rect 1104 3238 10880 3290
rect 10932 3238 10944 3290
rect 10996 3238 11008 3290
rect 11060 3238 11072 3290
rect 11124 3238 11136 3290
rect 11188 3238 20811 3290
rect 20863 3238 20875 3290
rect 20927 3238 20939 3290
rect 20991 3238 21003 3290
rect 21055 3238 21067 3290
rect 21119 3238 30820 3290
rect 1104 3216 30820 3238
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 29089 3179 29147 3185
rect 29089 3176 29101 3179
rect 27580 3148 29101 3176
rect 27580 3136 27586 3148
rect 29089 3145 29101 3148
rect 29135 3145 29147 3179
rect 29089 3139 29147 3145
rect 29825 3179 29883 3185
rect 29825 3145 29837 3179
rect 29871 3145 29883 3179
rect 29825 3139 29883 3145
rect 26602 3068 26608 3120
rect 26660 3108 26666 3120
rect 29840 3108 29868 3139
rect 26660 3080 29868 3108
rect 26660 3068 26666 3080
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 1486 3040 1492 3052
rect 1443 3012 1492 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 1486 3000 1492 3012
rect 1544 3000 1550 3052
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28868 3012 28917 3040
rect 28868 3000 28874 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 29730 3040 29736 3052
rect 29691 3012 29736 3040
rect 28905 3003 28963 3009
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1452 2808 1593 2836
rect 1452 2796 1458 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 1104 2746 30820 2768
rect 1104 2694 5915 2746
rect 5967 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 15846 2746
rect 15898 2694 15910 2746
rect 15962 2694 15974 2746
rect 16026 2694 16038 2746
rect 16090 2694 16102 2746
rect 16154 2694 25776 2746
rect 25828 2694 25840 2746
rect 25892 2694 25904 2746
rect 25956 2694 25968 2746
rect 26020 2694 26032 2746
rect 26084 2694 30820 2746
rect 1104 2672 30820 2694
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 28077 2635 28135 2641
rect 28077 2632 28089 2635
rect 26936 2604 28089 2632
rect 26936 2592 26942 2604
rect 28077 2601 28089 2604
rect 28123 2601 28135 2635
rect 28077 2595 28135 2601
rect 27890 2524 27896 2576
rect 27948 2564 27954 2576
rect 28905 2567 28963 2573
rect 28905 2564 28917 2567
rect 27948 2536 28917 2564
rect 27948 2524 27954 2536
rect 28905 2533 28917 2536
rect 28951 2533 28963 2567
rect 28905 2527 28963 2533
rect 18690 2496 18696 2508
rect 1412 2468 18696 2496
rect 1412 2437 1440 2468
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 2130 2428 2136 2440
rect 2091 2400 2136 2428
rect 1397 2391 1455 2397
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 16850 2428 16856 2440
rect 3099 2400 16856 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 28258 2428 28264 2440
rect 28219 2400 28264 2428
rect 28258 2388 28264 2400
rect 28316 2388 28322 2440
rect 28718 2428 28724 2440
rect 28679 2400 28724 2428
rect 28718 2388 28724 2400
rect 28776 2388 28782 2440
rect 29638 2428 29644 2440
rect 29599 2400 29644 2428
rect 29638 2388 29644 2400
rect 29696 2388 29702 2440
rect 25038 2320 25044 2372
rect 25096 2360 25102 2372
rect 29917 2363 29975 2369
rect 29917 2360 29929 2363
rect 25096 2332 29929 2360
rect 25096 2320 25102 2332
rect 29917 2329 29929 2332
rect 29963 2329 29975 2363
rect 29917 2323 29975 2329
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 2314 2292 2320 2304
rect 2275 2264 2320 2292
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 1104 2202 30820 2224
rect 1104 2150 10880 2202
rect 10932 2150 10944 2202
rect 10996 2150 11008 2202
rect 11060 2150 11072 2202
rect 11124 2150 11136 2202
rect 11188 2150 20811 2202
rect 20863 2150 20875 2202
rect 20927 2150 20939 2202
rect 20991 2150 21003 2202
rect 21055 2150 21067 2202
rect 21119 2150 30820 2202
rect 1104 2128 30820 2150
rect 22738 1300 22744 1352
rect 22796 1340 22802 1352
rect 28718 1340 28724 1352
rect 22796 1312 28724 1340
rect 22796 1300 22802 1312
rect 28718 1300 28724 1312
rect 28776 1300 28782 1352
<< via1 >>
rect 5915 77766 5967 77818
rect 5979 77766 6031 77818
rect 6043 77766 6095 77818
rect 6107 77766 6159 77818
rect 6171 77766 6223 77818
rect 15846 77766 15898 77818
rect 15910 77766 15962 77818
rect 15974 77766 16026 77818
rect 16038 77766 16090 77818
rect 16102 77766 16154 77818
rect 25776 77766 25828 77818
rect 25840 77766 25892 77818
rect 25904 77766 25956 77818
rect 25968 77766 26020 77818
rect 26032 77766 26084 77818
rect 27896 77664 27948 77716
rect 28172 77707 28224 77716
rect 28172 77673 28181 77707
rect 28181 77673 28215 77707
rect 28215 77673 28224 77707
rect 28172 77664 28224 77673
rect 1400 77571 1452 77580
rect 1400 77537 1409 77571
rect 1409 77537 1443 77571
rect 1443 77537 1452 77571
rect 1400 77528 1452 77537
rect 3792 77571 3844 77580
rect 3792 77537 3801 77571
rect 3801 77537 3835 77571
rect 3835 77537 3844 77571
rect 3792 77528 3844 77537
rect 11704 77460 11756 77512
rect 27252 77503 27304 77512
rect 27252 77469 27261 77503
rect 27261 77469 27295 77503
rect 27295 77469 27304 77503
rect 27252 77460 27304 77469
rect 27712 77460 27764 77512
rect 27160 77392 27212 77444
rect 29368 77460 29420 77512
rect 11796 77324 11848 77376
rect 28908 77367 28960 77376
rect 28908 77333 28917 77367
rect 28917 77333 28951 77367
rect 28951 77333 28960 77367
rect 28908 77324 28960 77333
rect 30104 77324 30156 77376
rect 10880 77222 10932 77274
rect 10944 77222 10996 77274
rect 11008 77222 11060 77274
rect 11072 77222 11124 77274
rect 11136 77222 11188 77274
rect 20811 77222 20863 77274
rect 20875 77222 20927 77274
rect 20939 77222 20991 77274
rect 21003 77222 21055 77274
rect 21067 77222 21119 77274
rect 28540 77163 28592 77172
rect 28540 77129 28549 77163
rect 28549 77129 28583 77163
rect 28583 77129 28592 77163
rect 28540 77120 28592 77129
rect 29276 77163 29328 77172
rect 29276 77129 29285 77163
rect 29285 77129 29319 77163
rect 29319 77129 29328 77163
rect 29276 77120 29328 77129
rect 2780 76984 2832 77036
rect 28356 77027 28408 77036
rect 28356 76993 28365 77027
rect 28365 76993 28399 77027
rect 28399 76993 28408 77027
rect 28356 76984 28408 76993
rect 29092 77027 29144 77036
rect 29092 76993 29101 77027
rect 29101 76993 29135 77027
rect 29135 76993 29144 77027
rect 29092 76984 29144 76993
rect 1400 76959 1452 76968
rect 1400 76925 1409 76959
rect 1409 76925 1443 76959
rect 1443 76925 1452 76959
rect 1400 76916 1452 76925
rect 13728 76916 13780 76968
rect 29000 76916 29052 76968
rect 8300 76848 8352 76900
rect 30012 76823 30064 76832
rect 30012 76789 30021 76823
rect 30021 76789 30055 76823
rect 30055 76789 30064 76823
rect 30012 76780 30064 76789
rect 5915 76678 5967 76730
rect 5979 76678 6031 76730
rect 6043 76678 6095 76730
rect 6107 76678 6159 76730
rect 6171 76678 6223 76730
rect 15846 76678 15898 76730
rect 15910 76678 15962 76730
rect 15974 76678 16026 76730
rect 16038 76678 16090 76730
rect 16102 76678 16154 76730
rect 25776 76678 25828 76730
rect 25840 76678 25892 76730
rect 25904 76678 25956 76730
rect 25968 76678 26020 76730
rect 26032 76678 26084 76730
rect 28816 76576 28868 76628
rect 1308 76440 1360 76492
rect 2872 76415 2924 76424
rect 2872 76381 2881 76415
rect 2881 76381 2915 76415
rect 2915 76381 2924 76415
rect 2872 76372 2924 76381
rect 26332 76372 26384 76424
rect 29736 76372 29788 76424
rect 10784 76304 10836 76356
rect 14648 76236 14700 76288
rect 19984 76236 20036 76288
rect 21180 76236 21232 76288
rect 30196 76236 30248 76288
rect 10880 76134 10932 76186
rect 10944 76134 10996 76186
rect 11008 76134 11060 76186
rect 11072 76134 11124 76186
rect 11136 76134 11188 76186
rect 20811 76134 20863 76186
rect 20875 76134 20927 76186
rect 20939 76134 20991 76186
rect 21003 76134 21055 76186
rect 21067 76134 21119 76186
rect 14556 76032 14608 76084
rect 29276 76075 29328 76084
rect 29276 76041 29285 76075
rect 29285 76041 29319 76075
rect 29319 76041 29328 76075
rect 29276 76032 29328 76041
rect 14648 76007 14700 76016
rect 14648 75973 14657 76007
rect 14657 75973 14691 76007
rect 14691 75973 14700 76007
rect 14648 75964 14700 75973
rect 15292 75964 15344 76016
rect 1584 75939 1636 75948
rect 1584 75905 1593 75939
rect 1593 75905 1627 75939
rect 1627 75905 1636 75939
rect 1584 75896 1636 75905
rect 14464 75939 14516 75948
rect 14464 75905 14473 75939
rect 14473 75905 14507 75939
rect 14507 75905 14516 75939
rect 14464 75896 14516 75905
rect 15752 75896 15804 75948
rect 16764 75896 16816 75948
rect 19064 75939 19116 75948
rect 19064 75905 19073 75939
rect 19073 75905 19107 75939
rect 19107 75905 19116 75939
rect 19064 75896 19116 75905
rect 19984 75939 20036 75948
rect 19984 75905 19993 75939
rect 19993 75905 20027 75939
rect 20027 75905 20036 75939
rect 19984 75896 20036 75905
rect 20168 75939 20220 75948
rect 20168 75905 20177 75939
rect 20177 75905 20211 75939
rect 20211 75905 20220 75939
rect 30104 75964 30156 76016
rect 20168 75896 20220 75905
rect 29828 75939 29880 75948
rect 29828 75905 29837 75939
rect 29837 75905 29871 75939
rect 29871 75905 29880 75939
rect 29828 75896 29880 75905
rect 21548 75828 21600 75880
rect 19892 75760 19944 75812
rect 15200 75692 15252 75744
rect 17040 75735 17092 75744
rect 17040 75701 17049 75735
rect 17049 75701 17083 75735
rect 17083 75701 17092 75735
rect 17040 75692 17092 75701
rect 19616 75692 19668 75744
rect 19708 75735 19760 75744
rect 19708 75701 19717 75735
rect 19717 75701 19751 75735
rect 19751 75701 19760 75735
rect 30012 75735 30064 75744
rect 19708 75692 19760 75701
rect 30012 75701 30021 75735
rect 30021 75701 30055 75735
rect 30055 75701 30064 75735
rect 30012 75692 30064 75701
rect 5915 75590 5967 75642
rect 5979 75590 6031 75642
rect 6043 75590 6095 75642
rect 6107 75590 6159 75642
rect 6171 75590 6223 75642
rect 15846 75590 15898 75642
rect 15910 75590 15962 75642
rect 15974 75590 16026 75642
rect 16038 75590 16090 75642
rect 16102 75590 16154 75642
rect 25776 75590 25828 75642
rect 25840 75590 25892 75642
rect 25904 75590 25956 75642
rect 25968 75590 26020 75642
rect 26032 75590 26084 75642
rect 21180 75531 21232 75540
rect 21180 75497 21189 75531
rect 21189 75497 21223 75531
rect 21223 75497 21232 75531
rect 21180 75488 21232 75497
rect 22376 75420 22428 75472
rect 15200 75395 15252 75404
rect 15200 75361 15209 75395
rect 15209 75361 15243 75395
rect 15243 75361 15252 75395
rect 15200 75352 15252 75361
rect 17040 75352 17092 75404
rect 19616 75352 19668 75404
rect 1584 75327 1636 75336
rect 1584 75293 1593 75327
rect 1593 75293 1627 75327
rect 1627 75293 1636 75327
rect 1584 75284 1636 75293
rect 14556 75327 14608 75336
rect 14556 75293 14565 75327
rect 14565 75293 14599 75327
rect 14599 75293 14608 75327
rect 14556 75284 14608 75293
rect 19708 75284 19760 75336
rect 29920 75284 29972 75336
rect 14464 75216 14516 75268
rect 16672 75216 16724 75268
rect 16856 75216 16908 75268
rect 19892 75216 19944 75268
rect 21272 75216 21324 75268
rect 14648 75148 14700 75200
rect 16948 75148 17000 75200
rect 17040 75148 17092 75200
rect 21180 75148 21232 75200
rect 24952 75148 25004 75200
rect 30196 75148 30248 75200
rect 10880 75046 10932 75098
rect 10944 75046 10996 75098
rect 11008 75046 11060 75098
rect 11072 75046 11124 75098
rect 11136 75046 11188 75098
rect 20811 75046 20863 75098
rect 20875 75046 20927 75098
rect 20939 75046 20991 75098
rect 21003 75046 21055 75098
rect 21067 75046 21119 75098
rect 15292 74944 15344 74996
rect 21456 74944 21508 74996
rect 14648 74919 14700 74928
rect 14648 74885 14657 74919
rect 14657 74885 14691 74919
rect 14691 74885 14700 74919
rect 14648 74876 14700 74885
rect 17224 74919 17276 74928
rect 17224 74885 17233 74919
rect 17233 74885 17267 74919
rect 17267 74885 17276 74919
rect 17224 74876 17276 74885
rect 20168 74876 20220 74928
rect 20720 74876 20772 74928
rect 1584 74851 1636 74860
rect 1584 74817 1593 74851
rect 1593 74817 1627 74851
rect 1627 74817 1636 74851
rect 1584 74808 1636 74817
rect 14556 74808 14608 74860
rect 16488 74808 16540 74860
rect 17960 74808 18012 74860
rect 21272 74851 21324 74860
rect 16580 74740 16632 74792
rect 18236 74783 18288 74792
rect 18236 74749 18245 74783
rect 18245 74749 18279 74783
rect 18279 74749 18288 74783
rect 18236 74740 18288 74749
rect 16764 74715 16816 74724
rect 16764 74681 16773 74715
rect 16773 74681 16807 74715
rect 16807 74681 16816 74715
rect 16764 74672 16816 74681
rect 21272 74817 21281 74851
rect 21281 74817 21315 74851
rect 21315 74817 21324 74851
rect 21272 74808 21324 74817
rect 21364 74808 21416 74860
rect 27436 74808 27488 74860
rect 21548 74740 21600 74792
rect 21824 74783 21876 74792
rect 21824 74749 21833 74783
rect 21833 74749 21867 74783
rect 21867 74749 21876 74783
rect 21824 74740 21876 74749
rect 20076 74604 20128 74656
rect 21272 74604 21324 74656
rect 22560 74604 22612 74656
rect 22836 74604 22888 74656
rect 30012 74647 30064 74656
rect 30012 74613 30021 74647
rect 30021 74613 30055 74647
rect 30055 74613 30064 74647
rect 30012 74604 30064 74613
rect 5915 74502 5967 74554
rect 5979 74502 6031 74554
rect 6043 74502 6095 74554
rect 6107 74502 6159 74554
rect 6171 74502 6223 74554
rect 15846 74502 15898 74554
rect 15910 74502 15962 74554
rect 15974 74502 16026 74554
rect 16038 74502 16090 74554
rect 16102 74502 16154 74554
rect 25776 74502 25828 74554
rect 25840 74502 25892 74554
rect 25904 74502 25956 74554
rect 25968 74502 26020 74554
rect 26032 74502 26084 74554
rect 15752 74400 15804 74452
rect 18236 74400 18288 74452
rect 16488 74307 16540 74316
rect 16488 74273 16497 74307
rect 16497 74273 16531 74307
rect 16531 74273 16540 74307
rect 16488 74264 16540 74273
rect 19064 74332 19116 74384
rect 18420 74264 18472 74316
rect 19892 74400 19944 74452
rect 21824 74400 21876 74452
rect 20444 74239 20496 74248
rect 20444 74205 20453 74239
rect 20453 74205 20487 74239
rect 20487 74205 20496 74239
rect 20444 74196 20496 74205
rect 21180 74239 21232 74248
rect 21180 74205 21189 74239
rect 21189 74205 21223 74239
rect 21223 74205 21232 74239
rect 21180 74196 21232 74205
rect 21272 74196 21324 74248
rect 26240 74196 26292 74248
rect 14556 74171 14608 74180
rect 14556 74137 14565 74171
rect 14565 74137 14599 74171
rect 14599 74137 14608 74171
rect 14556 74128 14608 74137
rect 14740 74171 14792 74180
rect 14740 74137 14749 74171
rect 14749 74137 14783 74171
rect 14783 74137 14792 74171
rect 14740 74128 14792 74137
rect 16580 74171 16632 74180
rect 16580 74137 16589 74171
rect 16589 74137 16623 74171
rect 16623 74137 16632 74171
rect 16580 74128 16632 74137
rect 19524 74128 19576 74180
rect 19892 74171 19944 74180
rect 19892 74137 19901 74171
rect 19901 74137 19935 74171
rect 19935 74137 19944 74171
rect 19892 74128 19944 74137
rect 17224 74060 17276 74112
rect 19708 74060 19760 74112
rect 22652 74060 22704 74112
rect 30196 74060 30248 74112
rect 10880 73958 10932 74010
rect 10944 73958 10996 74010
rect 11008 73958 11060 74010
rect 11072 73958 11124 74010
rect 11136 73958 11188 74010
rect 20811 73958 20863 74010
rect 20875 73958 20927 74010
rect 20939 73958 20991 74010
rect 21003 73958 21055 74010
rect 21067 73958 21119 74010
rect 14556 73856 14608 73908
rect 16672 73899 16724 73908
rect 16672 73865 16681 73899
rect 16681 73865 16715 73899
rect 16715 73865 16724 73899
rect 16672 73856 16724 73865
rect 17960 73899 18012 73908
rect 17960 73865 17969 73899
rect 17969 73865 18003 73899
rect 18003 73865 18012 73899
rect 17960 73856 18012 73865
rect 19708 73899 19760 73908
rect 19708 73865 19717 73899
rect 19717 73865 19751 73899
rect 19751 73865 19760 73899
rect 19708 73856 19760 73865
rect 21364 73856 21416 73908
rect 1584 73763 1636 73772
rect 1584 73729 1593 73763
rect 1593 73729 1627 73763
rect 1627 73729 1636 73763
rect 1584 73720 1636 73729
rect 13544 73720 13596 73772
rect 16948 73763 17000 73772
rect 16948 73729 16957 73763
rect 16957 73729 16991 73763
rect 16991 73729 17000 73763
rect 16948 73720 17000 73729
rect 17868 73788 17920 73840
rect 19524 73831 19576 73840
rect 17500 73720 17552 73772
rect 18236 73763 18288 73772
rect 18236 73729 18245 73763
rect 18245 73729 18279 73763
rect 18279 73729 18288 73763
rect 18236 73720 18288 73729
rect 19524 73797 19533 73831
rect 19533 73797 19567 73831
rect 19567 73797 19576 73831
rect 19524 73788 19576 73797
rect 14740 73584 14792 73636
rect 17316 73584 17368 73636
rect 18420 73584 18472 73636
rect 19892 73652 19944 73704
rect 20444 73584 20496 73636
rect 18236 73516 18288 73568
rect 20076 73516 20128 73568
rect 21088 73763 21140 73772
rect 21088 73729 21097 73763
rect 21097 73729 21131 73763
rect 21131 73729 21140 73763
rect 21088 73720 21140 73729
rect 21456 73720 21508 73772
rect 27344 73720 27396 73772
rect 21364 73652 21416 73704
rect 21548 73652 21600 73704
rect 22836 73516 22888 73568
rect 30012 73559 30064 73568
rect 30012 73525 30021 73559
rect 30021 73525 30055 73559
rect 30055 73525 30064 73559
rect 30012 73516 30064 73525
rect 5915 73414 5967 73466
rect 5979 73414 6031 73466
rect 6043 73414 6095 73466
rect 6107 73414 6159 73466
rect 6171 73414 6223 73466
rect 15846 73414 15898 73466
rect 15910 73414 15962 73466
rect 15974 73414 16026 73466
rect 16038 73414 16090 73466
rect 16102 73414 16154 73466
rect 25776 73414 25828 73466
rect 25840 73414 25892 73466
rect 25904 73414 25956 73466
rect 25968 73414 26020 73466
rect 26032 73414 26084 73466
rect 17500 73312 17552 73364
rect 19524 73312 19576 73364
rect 19708 73312 19760 73364
rect 21180 73312 21232 73364
rect 16948 73244 17000 73296
rect 1584 73151 1636 73160
rect 1584 73117 1593 73151
rect 1593 73117 1627 73151
rect 1627 73117 1636 73151
rect 1584 73108 1636 73117
rect 9588 73040 9640 73092
rect 10232 72972 10284 73024
rect 15844 73151 15896 73160
rect 15844 73117 15853 73151
rect 15853 73117 15887 73151
rect 15887 73117 15896 73151
rect 15844 73108 15896 73117
rect 17316 73176 17368 73228
rect 14648 73083 14700 73092
rect 14648 73049 14657 73083
rect 14657 73049 14691 73083
rect 14691 73049 14700 73083
rect 14648 73040 14700 73049
rect 14740 73040 14792 73092
rect 14924 73040 14976 73092
rect 16856 73040 16908 73092
rect 17408 73151 17460 73160
rect 17408 73117 17417 73151
rect 17417 73117 17451 73151
rect 17451 73117 17460 73151
rect 20536 73151 20588 73160
rect 17408 73108 17460 73117
rect 17040 72972 17092 73024
rect 19708 73083 19760 73092
rect 17868 72972 17920 73024
rect 19708 73049 19717 73083
rect 19717 73049 19751 73083
rect 19751 73049 19760 73083
rect 19708 73040 19760 73049
rect 20536 73117 20545 73151
rect 20545 73117 20579 73151
rect 20579 73117 20588 73151
rect 20536 73108 20588 73117
rect 26792 73108 26844 73160
rect 26148 73040 26200 73092
rect 20720 72972 20772 73024
rect 30012 73015 30064 73024
rect 30012 72981 30021 73015
rect 30021 72981 30055 73015
rect 30055 72981 30064 73015
rect 30012 72972 30064 72981
rect 10880 72870 10932 72922
rect 10944 72870 10996 72922
rect 11008 72870 11060 72922
rect 11072 72870 11124 72922
rect 11136 72870 11188 72922
rect 20811 72870 20863 72922
rect 20875 72870 20927 72922
rect 20939 72870 20991 72922
rect 21003 72870 21055 72922
rect 21067 72870 21119 72922
rect 10232 72700 10284 72752
rect 16488 72700 16540 72752
rect 1584 72675 1636 72684
rect 1584 72641 1593 72675
rect 1593 72641 1627 72675
rect 1627 72641 1636 72675
rect 1584 72632 1636 72641
rect 14648 72675 14700 72684
rect 14648 72641 14657 72675
rect 14657 72641 14691 72675
rect 14691 72641 14700 72675
rect 14648 72632 14700 72641
rect 14924 72632 14976 72684
rect 17132 72675 17184 72684
rect 17132 72641 17141 72675
rect 17141 72641 17175 72675
rect 17175 72641 17184 72675
rect 17132 72632 17184 72641
rect 29644 72632 29696 72684
rect 18236 72564 18288 72616
rect 17960 72496 18012 72548
rect 14832 72428 14884 72480
rect 17224 72471 17276 72480
rect 17224 72437 17233 72471
rect 17233 72437 17267 72471
rect 17267 72437 17276 72471
rect 17224 72428 17276 72437
rect 30012 72471 30064 72480
rect 30012 72437 30021 72471
rect 30021 72437 30055 72471
rect 30055 72437 30064 72471
rect 30012 72428 30064 72437
rect 5915 72326 5967 72378
rect 5979 72326 6031 72378
rect 6043 72326 6095 72378
rect 6107 72326 6159 72378
rect 6171 72326 6223 72378
rect 15846 72326 15898 72378
rect 15910 72326 15962 72378
rect 15974 72326 16026 72378
rect 16038 72326 16090 72378
rect 16102 72326 16154 72378
rect 25776 72326 25828 72378
rect 25840 72326 25892 72378
rect 25904 72326 25956 72378
rect 25968 72326 26020 72378
rect 26032 72326 26084 72378
rect 14648 72224 14700 72276
rect 14740 72156 14792 72208
rect 1584 72063 1636 72072
rect 1584 72029 1593 72063
rect 1593 72029 1627 72063
rect 1627 72029 1636 72063
rect 1584 72020 1636 72029
rect 13544 72063 13596 72072
rect 13544 72029 13553 72063
rect 13553 72029 13587 72063
rect 13587 72029 13596 72063
rect 13544 72020 13596 72029
rect 14648 72063 14700 72072
rect 14648 72029 14657 72063
rect 14657 72029 14691 72063
rect 14691 72029 14700 72063
rect 14648 72020 14700 72029
rect 14832 72063 14884 72072
rect 14832 72029 14841 72063
rect 14841 72029 14875 72063
rect 14875 72029 14884 72063
rect 14832 72020 14884 72029
rect 18144 72224 18196 72276
rect 17868 72088 17920 72140
rect 17316 72063 17368 72072
rect 17316 72029 17325 72063
rect 17325 72029 17359 72063
rect 17359 72029 17368 72063
rect 17316 72020 17368 72029
rect 30196 72020 30248 72072
rect 16948 71884 17000 71936
rect 30012 71927 30064 71936
rect 30012 71893 30021 71927
rect 30021 71893 30055 71927
rect 30055 71893 30064 71927
rect 30012 71884 30064 71893
rect 10880 71782 10932 71834
rect 10944 71782 10996 71834
rect 11008 71782 11060 71834
rect 11072 71782 11124 71834
rect 11136 71782 11188 71834
rect 20811 71782 20863 71834
rect 20875 71782 20927 71834
rect 20939 71782 20991 71834
rect 21003 71782 21055 71834
rect 21067 71782 21119 71834
rect 17316 71680 17368 71732
rect 8300 71612 8352 71664
rect 12808 71587 12860 71596
rect 12808 71553 12817 71587
rect 12817 71553 12851 71587
rect 12851 71553 12860 71587
rect 12808 71544 12860 71553
rect 17500 71544 17552 71596
rect 21272 71612 21324 71664
rect 17960 71587 18012 71596
rect 17960 71553 17969 71587
rect 17969 71553 18003 71587
rect 18003 71553 18012 71587
rect 17960 71544 18012 71553
rect 21456 71544 21508 71596
rect 30840 71544 30892 71596
rect 17868 71476 17920 71528
rect 18420 71476 18472 71528
rect 19340 71476 19392 71528
rect 22468 71408 22520 71460
rect 17960 71340 18012 71392
rect 19800 71340 19852 71392
rect 21364 71340 21416 71392
rect 30012 71383 30064 71392
rect 30012 71349 30021 71383
rect 30021 71349 30055 71383
rect 30055 71349 30064 71383
rect 30012 71340 30064 71349
rect 5915 71238 5967 71290
rect 5979 71238 6031 71290
rect 6043 71238 6095 71290
rect 6107 71238 6159 71290
rect 6171 71238 6223 71290
rect 15846 71238 15898 71290
rect 15910 71238 15962 71290
rect 15974 71238 16026 71290
rect 16038 71238 16090 71290
rect 16102 71238 16154 71290
rect 25776 71238 25828 71290
rect 25840 71238 25892 71290
rect 25904 71238 25956 71290
rect 25968 71238 26020 71290
rect 26032 71238 26084 71290
rect 16396 71136 16448 71188
rect 18236 71179 18288 71188
rect 18236 71145 18245 71179
rect 18245 71145 18279 71179
rect 18279 71145 18288 71179
rect 18236 71136 18288 71145
rect 20720 71136 20772 71188
rect 19524 71068 19576 71120
rect 1492 71000 1544 71052
rect 1400 70975 1452 70984
rect 1400 70941 1409 70975
rect 1409 70941 1443 70975
rect 1443 70941 1452 70975
rect 1400 70932 1452 70941
rect 9588 70932 9640 70984
rect 16488 71000 16540 71052
rect 11796 70932 11848 70984
rect 12808 70907 12860 70916
rect 12808 70873 12817 70907
rect 12817 70873 12851 70907
rect 12851 70873 12860 70907
rect 12808 70864 12860 70873
rect 16580 70932 16632 70984
rect 17408 70932 17460 70984
rect 30288 70932 30340 70984
rect 14648 70907 14700 70916
rect 14648 70873 14657 70907
rect 14657 70873 14691 70907
rect 14691 70873 14700 70907
rect 14648 70864 14700 70873
rect 18420 70864 18472 70916
rect 19616 70907 19668 70916
rect 19616 70873 19625 70907
rect 19625 70873 19659 70907
rect 19659 70873 19668 70907
rect 19616 70864 19668 70873
rect 15568 70796 15620 70848
rect 17224 70796 17276 70848
rect 30012 70839 30064 70848
rect 30012 70805 30021 70839
rect 30021 70805 30055 70839
rect 30055 70805 30064 70839
rect 30012 70796 30064 70805
rect 10880 70694 10932 70746
rect 10944 70694 10996 70746
rect 11008 70694 11060 70746
rect 11072 70694 11124 70746
rect 11136 70694 11188 70746
rect 20811 70694 20863 70746
rect 20875 70694 20927 70746
rect 20939 70694 20991 70746
rect 21003 70694 21055 70746
rect 21067 70694 21119 70746
rect 1492 70592 1544 70644
rect 12808 70592 12860 70644
rect 11704 70524 11756 70576
rect 15476 70524 15528 70576
rect 1584 70499 1636 70508
rect 1584 70465 1593 70499
rect 1593 70465 1627 70499
rect 1627 70465 1636 70499
rect 1584 70456 1636 70465
rect 12808 70499 12860 70508
rect 12808 70465 12817 70499
rect 12817 70465 12851 70499
rect 12851 70465 12860 70499
rect 12808 70456 12860 70465
rect 13728 70456 13780 70508
rect 15568 70499 15620 70508
rect 13544 70388 13596 70440
rect 14832 70388 14884 70440
rect 15568 70465 15577 70499
rect 15577 70465 15611 70499
rect 15611 70465 15620 70499
rect 15568 70456 15620 70465
rect 18144 70592 18196 70644
rect 18328 70592 18380 70644
rect 19708 70592 19760 70644
rect 19984 70635 20036 70644
rect 19984 70601 19993 70635
rect 19993 70601 20027 70635
rect 20027 70601 20036 70635
rect 19984 70592 20036 70601
rect 22376 70524 22428 70576
rect 16948 70456 17000 70508
rect 19432 70456 19484 70508
rect 19524 70456 19576 70508
rect 19708 70456 19760 70508
rect 20812 70456 20864 70508
rect 22008 70456 22060 70508
rect 16764 70388 16816 70440
rect 21364 70388 21416 70440
rect 22284 70499 22336 70508
rect 22284 70465 22298 70499
rect 22298 70465 22332 70499
rect 22332 70465 22336 70499
rect 22284 70456 22336 70465
rect 29184 70456 29236 70508
rect 15752 70295 15804 70304
rect 15752 70261 15761 70295
rect 15761 70261 15795 70295
rect 15795 70261 15804 70295
rect 15752 70252 15804 70261
rect 21088 70295 21140 70304
rect 21088 70261 21097 70295
rect 21097 70261 21131 70295
rect 21131 70261 21140 70295
rect 21088 70252 21140 70261
rect 21824 70295 21876 70304
rect 21824 70261 21833 70295
rect 21833 70261 21867 70295
rect 21867 70261 21876 70295
rect 21824 70252 21876 70261
rect 30012 70295 30064 70304
rect 30012 70261 30021 70295
rect 30021 70261 30055 70295
rect 30055 70261 30064 70295
rect 30012 70252 30064 70261
rect 5915 70150 5967 70202
rect 5979 70150 6031 70202
rect 6043 70150 6095 70202
rect 6107 70150 6159 70202
rect 6171 70150 6223 70202
rect 15846 70150 15898 70202
rect 15910 70150 15962 70202
rect 15974 70150 16026 70202
rect 16038 70150 16090 70202
rect 16102 70150 16154 70202
rect 25776 70150 25828 70202
rect 25840 70150 25892 70202
rect 25904 70150 25956 70202
rect 25968 70150 26020 70202
rect 26032 70150 26084 70202
rect 18512 70048 18564 70100
rect 20812 70048 20864 70100
rect 22008 70048 22060 70100
rect 24216 70048 24268 70100
rect 29092 69980 29144 70032
rect 1584 69887 1636 69896
rect 1584 69853 1593 69887
rect 1593 69853 1627 69887
rect 1627 69853 1636 69887
rect 1584 69844 1636 69853
rect 10784 69844 10836 69896
rect 12808 69887 12860 69896
rect 12808 69853 12817 69887
rect 12817 69853 12851 69887
rect 12851 69853 12860 69887
rect 12808 69844 12860 69853
rect 15752 69844 15804 69896
rect 21088 69844 21140 69896
rect 22284 69887 22336 69896
rect 22284 69853 22293 69887
rect 22293 69853 22327 69887
rect 22327 69853 22336 69887
rect 22284 69844 22336 69853
rect 14648 69776 14700 69828
rect 18052 69776 18104 69828
rect 19524 69776 19576 69828
rect 19800 69819 19852 69828
rect 19800 69785 19809 69819
rect 19809 69785 19843 69819
rect 19843 69785 19852 69819
rect 19800 69776 19852 69785
rect 19892 69819 19944 69828
rect 19892 69785 19901 69819
rect 19901 69785 19935 69819
rect 19935 69785 19944 69819
rect 19892 69776 19944 69785
rect 21824 69776 21876 69828
rect 21916 69776 21968 69828
rect 9956 69708 10008 69760
rect 16212 69708 16264 69760
rect 17132 69708 17184 69760
rect 17408 69708 17460 69760
rect 22100 69708 22152 69760
rect 25504 69708 25556 69760
rect 29000 69708 29052 69760
rect 30656 69844 30708 69896
rect 30012 69751 30064 69760
rect 30012 69717 30021 69751
rect 30021 69717 30055 69751
rect 30055 69717 30064 69751
rect 30012 69708 30064 69717
rect 10880 69606 10932 69658
rect 10944 69606 10996 69658
rect 11008 69606 11060 69658
rect 11072 69606 11124 69658
rect 11136 69606 11188 69658
rect 20811 69606 20863 69658
rect 20875 69606 20927 69658
rect 20939 69606 20991 69658
rect 21003 69606 21055 69658
rect 21067 69606 21119 69658
rect 21916 69504 21968 69556
rect 29184 69504 29236 69556
rect 29828 69504 29880 69556
rect 9956 69436 10008 69488
rect 17960 69436 18012 69488
rect 20628 69436 20680 69488
rect 1584 69411 1636 69420
rect 1584 69377 1593 69411
rect 1593 69377 1627 69411
rect 1627 69377 1636 69411
rect 1584 69368 1636 69377
rect 12624 69368 12676 69420
rect 14004 69368 14056 69420
rect 17316 69368 17368 69420
rect 13912 69343 13964 69352
rect 13912 69309 13921 69343
rect 13921 69309 13955 69343
rect 13955 69309 13964 69343
rect 13912 69300 13964 69309
rect 16672 69300 16724 69352
rect 20444 69368 20496 69420
rect 21456 69368 21508 69420
rect 22100 69411 22152 69420
rect 22100 69377 22109 69411
rect 22109 69377 22143 69411
rect 22143 69377 22152 69411
rect 22100 69368 22152 69377
rect 22376 69436 22428 69488
rect 29552 69436 29604 69488
rect 29736 69436 29788 69488
rect 22468 69411 22520 69420
rect 18144 69343 18196 69352
rect 18144 69309 18153 69343
rect 18153 69309 18187 69343
rect 18187 69309 18196 69343
rect 18144 69300 18196 69309
rect 19708 69300 19760 69352
rect 20260 69300 20312 69352
rect 22468 69377 22477 69411
rect 22477 69377 22511 69411
rect 22511 69377 22520 69411
rect 22468 69368 22520 69377
rect 28448 69368 28500 69420
rect 29368 69300 29420 69352
rect 22192 69232 22244 69284
rect 29276 69275 29328 69284
rect 29276 69241 29285 69275
rect 29285 69241 29319 69275
rect 29319 69241 29328 69275
rect 29276 69232 29328 69241
rect 11336 69164 11388 69216
rect 14832 69164 14884 69216
rect 16304 69164 16356 69216
rect 19340 69164 19392 69216
rect 19708 69164 19760 69216
rect 29920 69164 29972 69216
rect 5915 69062 5967 69114
rect 5979 69062 6031 69114
rect 6043 69062 6095 69114
rect 6107 69062 6159 69114
rect 6171 69062 6223 69114
rect 15846 69062 15898 69114
rect 15910 69062 15962 69114
rect 15974 69062 16026 69114
rect 16038 69062 16090 69114
rect 16102 69062 16154 69114
rect 25776 69062 25828 69114
rect 25840 69062 25892 69114
rect 25904 69062 25956 69114
rect 25968 69062 26020 69114
rect 26032 69062 26084 69114
rect 14648 69003 14700 69012
rect 14648 68969 14657 69003
rect 14657 68969 14691 69003
rect 14691 68969 14700 69003
rect 14648 68960 14700 68969
rect 16764 68960 16816 69012
rect 20536 68960 20588 69012
rect 22284 68960 22336 69012
rect 1584 68799 1636 68808
rect 1584 68765 1593 68799
rect 1593 68765 1627 68799
rect 1627 68765 1636 68799
rect 1584 68756 1636 68765
rect 12624 68799 12676 68808
rect 12624 68765 12633 68799
rect 12633 68765 12667 68799
rect 12667 68765 12676 68799
rect 12624 68756 12676 68765
rect 16212 68892 16264 68944
rect 24768 68892 24820 68944
rect 14832 68824 14884 68876
rect 12808 68731 12860 68740
rect 12808 68697 12817 68731
rect 12817 68697 12851 68731
rect 12851 68697 12860 68731
rect 12808 68688 12860 68697
rect 14188 68688 14240 68740
rect 15200 68756 15252 68808
rect 17500 68824 17552 68876
rect 20352 68824 20404 68876
rect 19984 68756 20036 68808
rect 20076 68756 20128 68808
rect 27252 68756 27304 68808
rect 29276 68756 29328 68808
rect 17316 68731 17368 68740
rect 17316 68697 17325 68731
rect 17325 68697 17359 68731
rect 17359 68697 17368 68731
rect 17316 68688 17368 68697
rect 18604 68731 18656 68740
rect 18604 68697 18613 68731
rect 18613 68697 18647 68731
rect 18647 68697 18656 68731
rect 18604 68688 18656 68697
rect 19800 68688 19852 68740
rect 20444 68731 20496 68740
rect 20444 68697 20453 68731
rect 20453 68697 20487 68731
rect 20487 68697 20496 68731
rect 20444 68688 20496 68697
rect 20536 68731 20588 68740
rect 20536 68697 20545 68731
rect 20545 68697 20579 68731
rect 20579 68697 20588 68731
rect 20536 68688 20588 68697
rect 1400 68663 1452 68672
rect 1400 68629 1409 68663
rect 1409 68629 1443 68663
rect 1443 68629 1452 68663
rect 1400 68620 1452 68629
rect 14464 68620 14516 68672
rect 20628 68620 20680 68672
rect 28908 68663 28960 68672
rect 28908 68629 28917 68663
rect 28917 68629 28951 68663
rect 28951 68629 28960 68663
rect 28908 68620 28960 68629
rect 30012 68663 30064 68672
rect 30012 68629 30021 68663
rect 30021 68629 30055 68663
rect 30055 68629 30064 68663
rect 30012 68620 30064 68629
rect 10880 68518 10932 68570
rect 10944 68518 10996 68570
rect 11008 68518 11060 68570
rect 11072 68518 11124 68570
rect 11136 68518 11188 68570
rect 20811 68518 20863 68570
rect 20875 68518 20927 68570
rect 20939 68518 20991 68570
rect 21003 68518 21055 68570
rect 21067 68518 21119 68570
rect 1400 68416 1452 68468
rect 12808 68416 12860 68468
rect 13912 68416 13964 68468
rect 13820 68280 13872 68332
rect 16304 68416 16356 68468
rect 20444 68416 20496 68468
rect 29460 68416 29512 68468
rect 15200 68348 15252 68400
rect 18236 68348 18288 68400
rect 19524 68391 19576 68400
rect 19524 68357 19533 68391
rect 19533 68357 19567 68391
rect 19567 68357 19576 68391
rect 19524 68348 19576 68357
rect 20352 68391 20404 68400
rect 20352 68357 20361 68391
rect 20361 68357 20395 68391
rect 20395 68357 20404 68391
rect 20352 68348 20404 68357
rect 14464 68323 14516 68332
rect 14464 68289 14473 68323
rect 14473 68289 14507 68323
rect 14507 68289 14516 68323
rect 14464 68280 14516 68289
rect 20720 68280 20772 68332
rect 26424 68280 26476 68332
rect 14924 68212 14976 68264
rect 14004 68144 14056 68196
rect 14188 68144 14240 68196
rect 20076 68187 20128 68196
rect 20076 68153 20085 68187
rect 20085 68153 20119 68187
rect 20119 68153 20128 68187
rect 20076 68144 20128 68153
rect 20536 68212 20588 68264
rect 21180 68212 21232 68264
rect 27068 68212 27120 68264
rect 27528 68280 27580 68332
rect 22468 68144 22520 68196
rect 26516 68144 26568 68196
rect 17316 68076 17368 68128
rect 30472 68280 30524 68332
rect 29920 68076 29972 68128
rect 5915 67974 5967 68026
rect 5979 67974 6031 68026
rect 6043 67974 6095 68026
rect 6107 67974 6159 68026
rect 6171 67974 6223 68026
rect 15846 67974 15898 68026
rect 15910 67974 15962 68026
rect 15974 67974 16026 68026
rect 16038 67974 16090 68026
rect 16102 67974 16154 68026
rect 25776 67974 25828 68026
rect 25840 67974 25892 68026
rect 25904 67974 25956 68026
rect 25968 67974 26020 68026
rect 26032 67974 26084 68026
rect 18144 67872 18196 67924
rect 26240 67915 26292 67924
rect 26240 67881 26249 67915
rect 26249 67881 26283 67915
rect 26283 67881 26292 67915
rect 26240 67872 26292 67881
rect 27436 67872 27488 67924
rect 11244 67804 11296 67856
rect 21272 67847 21324 67856
rect 21272 67813 21281 67847
rect 21281 67813 21315 67847
rect 21315 67813 21324 67847
rect 21272 67804 21324 67813
rect 26056 67804 26108 67856
rect 26608 67804 26660 67856
rect 27068 67804 27120 67856
rect 27620 67804 27672 67856
rect 28908 67847 28960 67856
rect 28908 67813 28917 67847
rect 28917 67813 28951 67847
rect 28951 67813 28960 67847
rect 28908 67804 28960 67813
rect 30012 67847 30064 67856
rect 30012 67813 30021 67847
rect 30021 67813 30055 67847
rect 30055 67813 30064 67847
rect 30012 67804 30064 67813
rect 1584 67711 1636 67720
rect 1584 67677 1593 67711
rect 1593 67677 1627 67711
rect 1627 67677 1636 67711
rect 1584 67668 1636 67677
rect 11336 67668 11388 67720
rect 16672 67711 16724 67720
rect 16672 67677 16681 67711
rect 16681 67677 16715 67711
rect 16715 67677 16724 67711
rect 16672 67668 16724 67677
rect 17408 67711 17460 67720
rect 17408 67677 17417 67711
rect 17417 67677 17451 67711
rect 17451 67677 17460 67711
rect 17408 67668 17460 67677
rect 18696 67668 18748 67720
rect 25136 67668 25188 67720
rect 25412 67668 25464 67720
rect 12624 67600 12676 67652
rect 17592 67643 17644 67652
rect 17592 67609 17601 67643
rect 17601 67609 17635 67643
rect 17635 67609 17644 67643
rect 17592 67600 17644 67609
rect 19984 67643 20036 67652
rect 19984 67609 19993 67643
rect 19993 67609 20027 67643
rect 20027 67609 20036 67643
rect 19984 67600 20036 67609
rect 24952 67600 25004 67652
rect 25228 67643 25280 67652
rect 25228 67609 25237 67643
rect 25237 67609 25271 67643
rect 25271 67609 25280 67643
rect 25228 67600 25280 67609
rect 26700 67711 26752 67720
rect 26700 67677 26709 67711
rect 26709 67677 26743 67711
rect 26743 67677 26752 67711
rect 26700 67668 26752 67677
rect 26884 67711 26936 67720
rect 26884 67677 26893 67711
rect 26893 67677 26927 67711
rect 26927 67677 26936 67711
rect 26884 67668 26936 67677
rect 27068 67668 27120 67720
rect 27620 67711 27672 67720
rect 27620 67677 27629 67711
rect 27629 67677 27663 67711
rect 27663 67677 27672 67711
rect 27620 67668 27672 67677
rect 13084 67575 13136 67584
rect 13084 67541 13093 67575
rect 13093 67541 13127 67575
rect 13127 67541 13136 67575
rect 13084 67532 13136 67541
rect 15200 67532 15252 67584
rect 17684 67532 17736 67584
rect 25596 67532 25648 67584
rect 26148 67532 26200 67584
rect 27620 67532 27672 67584
rect 27804 67711 27856 67720
rect 27804 67677 27813 67711
rect 27813 67677 27847 67711
rect 27847 67677 27856 67711
rect 27804 67668 27856 67677
rect 29000 67668 29052 67720
rect 29460 67668 29512 67720
rect 27804 67532 27856 67584
rect 10880 67430 10932 67482
rect 10944 67430 10996 67482
rect 11008 67430 11060 67482
rect 11072 67430 11124 67482
rect 11136 67430 11188 67482
rect 20811 67430 20863 67482
rect 20875 67430 20927 67482
rect 20939 67430 20991 67482
rect 21003 67430 21055 67482
rect 21067 67430 21119 67482
rect 18604 67328 18656 67380
rect 26884 67328 26936 67380
rect 11244 67260 11296 67312
rect 13084 67260 13136 67312
rect 1584 67235 1636 67244
rect 1584 67201 1593 67235
rect 1593 67201 1627 67235
rect 1627 67201 1636 67235
rect 1584 67192 1636 67201
rect 12624 67235 12676 67244
rect 12624 67201 12633 67235
rect 12633 67201 12667 67235
rect 12667 67201 12676 67235
rect 12624 67192 12676 67201
rect 14924 67192 14976 67244
rect 19524 67260 19576 67312
rect 14188 67124 14240 67176
rect 14556 67056 14608 67108
rect 15200 67056 15252 67108
rect 19708 67192 19760 67244
rect 23572 67192 23624 67244
rect 25136 67192 25188 67244
rect 17040 67124 17092 67176
rect 18696 67099 18748 67108
rect 18696 67065 18705 67099
rect 18705 67065 18739 67099
rect 18739 67065 18748 67099
rect 18696 67056 18748 67065
rect 19892 67124 19944 67176
rect 20076 67124 20128 67176
rect 25412 67192 25464 67244
rect 26056 67192 26108 67244
rect 26240 67235 26292 67244
rect 26240 67201 26249 67235
rect 26249 67201 26283 67235
rect 26283 67201 26292 67235
rect 27620 67328 27672 67380
rect 27804 67328 27856 67380
rect 27896 67260 27948 67312
rect 26240 67192 26292 67201
rect 27620 67235 27672 67244
rect 25044 67056 25096 67108
rect 11244 66988 11296 67040
rect 14740 66988 14792 67040
rect 15384 66988 15436 67040
rect 23940 66988 23992 67040
rect 24860 66988 24912 67040
rect 25504 67124 25556 67176
rect 27068 67124 27120 67176
rect 27620 67201 27629 67235
rect 27629 67201 27663 67235
rect 27663 67201 27672 67235
rect 27620 67192 27672 67201
rect 28264 67192 28316 67244
rect 26884 67056 26936 67108
rect 27436 67056 27488 67108
rect 29092 67056 29144 67108
rect 28908 66988 28960 67040
rect 29828 66988 29880 67040
rect 5915 66886 5967 66938
rect 5979 66886 6031 66938
rect 6043 66886 6095 66938
rect 6107 66886 6159 66938
rect 6171 66886 6223 66938
rect 15846 66886 15898 66938
rect 15910 66886 15962 66938
rect 15974 66886 16026 66938
rect 16038 66886 16090 66938
rect 16102 66886 16154 66938
rect 25776 66886 25828 66938
rect 25840 66886 25892 66938
rect 25904 66886 25956 66938
rect 25968 66886 26020 66938
rect 26032 66886 26084 66938
rect 14924 66784 14976 66836
rect 18420 66827 18472 66836
rect 18420 66793 18429 66827
rect 18429 66793 18463 66827
rect 18463 66793 18472 66827
rect 18420 66784 18472 66793
rect 19616 66784 19668 66836
rect 22560 66784 22612 66836
rect 23572 66784 23624 66836
rect 26976 66784 27028 66836
rect 28816 66784 28868 66836
rect 29092 66784 29144 66836
rect 23296 66716 23348 66768
rect 26516 66716 26568 66768
rect 14188 66648 14240 66700
rect 1584 66623 1636 66632
rect 1584 66589 1593 66623
rect 1593 66589 1627 66623
rect 1627 66589 1636 66623
rect 1584 66580 1636 66589
rect 16396 66648 16448 66700
rect 14556 66623 14608 66632
rect 14556 66589 14565 66623
rect 14565 66589 14599 66623
rect 14599 66589 14608 66623
rect 14740 66623 14792 66632
rect 14556 66580 14608 66589
rect 14740 66589 14749 66623
rect 14749 66589 14783 66623
rect 14783 66589 14792 66623
rect 14740 66580 14792 66589
rect 15292 66623 15344 66632
rect 15292 66589 15301 66623
rect 15301 66589 15335 66623
rect 15335 66589 15344 66623
rect 15292 66580 15344 66589
rect 15384 66580 15436 66632
rect 14832 66512 14884 66564
rect 11336 66444 11388 66496
rect 14096 66487 14148 66496
rect 14096 66453 14105 66487
rect 14105 66453 14139 66487
rect 14139 66453 14148 66487
rect 14096 66444 14148 66453
rect 17132 66487 17184 66496
rect 17132 66453 17141 66487
rect 17141 66453 17175 66487
rect 17175 66453 17184 66487
rect 17132 66444 17184 66453
rect 17684 66580 17736 66632
rect 18328 66648 18380 66700
rect 18604 66580 18656 66632
rect 17868 66512 17920 66564
rect 20168 66648 20220 66700
rect 22836 66648 22888 66700
rect 20536 66623 20588 66632
rect 20536 66589 20545 66623
rect 20545 66589 20579 66623
rect 20579 66589 20588 66623
rect 20536 66580 20588 66589
rect 22560 66623 22612 66632
rect 22560 66589 22569 66623
rect 22569 66589 22603 66623
rect 22603 66589 22612 66623
rect 22560 66580 22612 66589
rect 23572 66580 23624 66632
rect 25228 66580 25280 66632
rect 24216 66512 24268 66564
rect 18420 66444 18472 66496
rect 20720 66487 20772 66496
rect 20720 66453 20729 66487
rect 20729 66453 20763 66487
rect 20763 66453 20772 66487
rect 20720 66444 20772 66453
rect 23388 66444 23440 66496
rect 23664 66487 23716 66496
rect 23664 66453 23673 66487
rect 23673 66453 23707 66487
rect 23707 66453 23716 66487
rect 23664 66444 23716 66453
rect 24676 66444 24728 66496
rect 25136 66512 25188 66564
rect 25412 66512 25464 66564
rect 26148 66580 26200 66632
rect 27252 66648 27304 66700
rect 26976 66580 27028 66632
rect 27620 66648 27672 66700
rect 27804 66691 27856 66700
rect 27804 66657 27813 66691
rect 27813 66657 27847 66691
rect 27847 66657 27856 66691
rect 27804 66648 27856 66657
rect 28816 66580 28868 66632
rect 27804 66512 27856 66564
rect 26976 66444 27028 66496
rect 10880 66342 10932 66394
rect 10944 66342 10996 66394
rect 11008 66342 11060 66394
rect 11072 66342 11124 66394
rect 11136 66342 11188 66394
rect 20811 66342 20863 66394
rect 20875 66342 20927 66394
rect 20939 66342 20991 66394
rect 21003 66342 21055 66394
rect 21067 66342 21119 66394
rect 27620 66240 27672 66292
rect 29460 66240 29512 66292
rect 11244 66172 11296 66224
rect 14096 66172 14148 66224
rect 17132 66172 17184 66224
rect 22376 66172 22428 66224
rect 23020 66172 23072 66224
rect 30104 66215 30156 66224
rect 30104 66181 30113 66215
rect 30113 66181 30147 66215
rect 30147 66181 30156 66215
rect 30104 66172 30156 66181
rect 1584 66147 1636 66156
rect 1584 66113 1593 66147
rect 1593 66113 1627 66147
rect 1627 66113 1636 66147
rect 1584 66104 1636 66113
rect 12624 66147 12676 66156
rect 12624 66113 12633 66147
rect 12633 66113 12667 66147
rect 12667 66113 12676 66147
rect 12624 66104 12676 66113
rect 16856 66104 16908 66156
rect 18696 66104 18748 66156
rect 21916 66104 21968 66156
rect 22560 66104 22612 66156
rect 23296 66147 23348 66156
rect 23296 66113 23305 66147
rect 23305 66113 23339 66147
rect 23339 66113 23348 66147
rect 23296 66104 23348 66113
rect 23572 66104 23624 66156
rect 25228 66147 25280 66156
rect 25228 66113 25237 66147
rect 25237 66113 25271 66147
rect 25271 66113 25280 66147
rect 25228 66104 25280 66113
rect 25412 66147 25464 66156
rect 25412 66113 25421 66147
rect 25421 66113 25455 66147
rect 25455 66113 25464 66147
rect 25412 66104 25464 66113
rect 26148 66104 26200 66156
rect 27988 66104 28040 66156
rect 28632 66147 28684 66156
rect 28632 66113 28641 66147
rect 28641 66113 28675 66147
rect 28675 66113 28684 66147
rect 28632 66104 28684 66113
rect 28724 66104 28776 66156
rect 13728 66079 13780 66088
rect 13728 66045 13737 66079
rect 13737 66045 13771 66079
rect 13771 66045 13780 66079
rect 13728 66036 13780 66045
rect 22376 66036 22428 66088
rect 28908 66036 28960 66088
rect 20628 65968 20680 66020
rect 11428 65900 11480 65952
rect 12992 65943 13044 65952
rect 12992 65909 13001 65943
rect 13001 65909 13035 65943
rect 13035 65909 13044 65943
rect 12992 65900 13044 65909
rect 14832 65900 14884 65952
rect 18420 65943 18472 65952
rect 18420 65909 18429 65943
rect 18429 65909 18463 65943
rect 18463 65909 18472 65943
rect 21824 65943 21876 65952
rect 18420 65900 18472 65909
rect 21824 65909 21833 65943
rect 21833 65909 21867 65943
rect 21867 65909 21876 65943
rect 21824 65900 21876 65909
rect 23480 65900 23532 65952
rect 24676 65900 24728 65952
rect 28080 65943 28132 65952
rect 28080 65909 28089 65943
rect 28089 65909 28123 65943
rect 28123 65909 28132 65943
rect 28080 65900 28132 65909
rect 28172 65900 28224 65952
rect 29552 65968 29604 66020
rect 30104 66036 30156 66088
rect 30380 65968 30432 66020
rect 29920 65900 29972 65952
rect 5915 65798 5967 65850
rect 5979 65798 6031 65850
rect 6043 65798 6095 65850
rect 6107 65798 6159 65850
rect 6171 65798 6223 65850
rect 15846 65798 15898 65850
rect 15910 65798 15962 65850
rect 15974 65798 16026 65850
rect 16038 65798 16090 65850
rect 16102 65798 16154 65850
rect 25776 65798 25828 65850
rect 25840 65798 25892 65850
rect 25904 65798 25956 65850
rect 25968 65798 26020 65850
rect 26032 65798 26084 65850
rect 12624 65696 12676 65748
rect 15292 65696 15344 65748
rect 16856 65739 16908 65748
rect 16856 65705 16865 65739
rect 16865 65705 16899 65739
rect 16899 65705 16908 65739
rect 16856 65696 16908 65705
rect 18052 65696 18104 65748
rect 19432 65739 19484 65748
rect 19432 65705 19441 65739
rect 19441 65705 19475 65739
rect 19475 65705 19484 65739
rect 19432 65696 19484 65705
rect 20536 65696 20588 65748
rect 27344 65696 27396 65748
rect 27804 65696 27856 65748
rect 17316 65603 17368 65612
rect 17316 65569 17325 65603
rect 17325 65569 17359 65603
rect 17359 65569 17368 65603
rect 17316 65560 17368 65569
rect 17500 65560 17552 65612
rect 20812 65628 20864 65680
rect 21180 65628 21232 65680
rect 24308 65628 24360 65680
rect 20720 65560 20772 65612
rect 25228 65603 25280 65612
rect 25228 65569 25237 65603
rect 25237 65569 25271 65603
rect 25271 65569 25280 65603
rect 25228 65560 25280 65569
rect 1584 65535 1636 65544
rect 1584 65501 1593 65535
rect 1593 65501 1627 65535
rect 1627 65501 1636 65535
rect 1584 65492 1636 65501
rect 12900 65535 12952 65544
rect 12900 65501 12909 65535
rect 12909 65501 12943 65535
rect 12943 65501 12952 65535
rect 12900 65492 12952 65501
rect 15292 65535 15344 65544
rect 15292 65501 15301 65535
rect 15301 65501 15335 65535
rect 15335 65501 15344 65535
rect 15292 65492 15344 65501
rect 19340 65492 19392 65544
rect 24584 65492 24636 65544
rect 27620 65492 27672 65544
rect 20260 65467 20312 65476
rect 20260 65433 20269 65467
rect 20269 65433 20303 65467
rect 20303 65433 20312 65467
rect 20260 65424 20312 65433
rect 21180 65424 21232 65476
rect 27896 65535 27948 65544
rect 27896 65501 27905 65535
rect 27905 65501 27939 65535
rect 27939 65501 27948 65535
rect 29920 65628 29972 65680
rect 31852 65628 31904 65680
rect 27896 65492 27948 65501
rect 29920 65492 29972 65544
rect 28448 65424 28500 65476
rect 11244 65356 11296 65408
rect 17592 65356 17644 65408
rect 20444 65399 20496 65408
rect 20444 65365 20453 65399
rect 20453 65365 20487 65399
rect 20487 65365 20496 65399
rect 20444 65356 20496 65365
rect 22744 65399 22796 65408
rect 22744 65365 22753 65399
rect 22753 65365 22787 65399
rect 22787 65365 22796 65399
rect 22744 65356 22796 65365
rect 28356 65356 28408 65408
rect 30564 65356 30616 65408
rect 10880 65254 10932 65306
rect 10944 65254 10996 65306
rect 11008 65254 11060 65306
rect 11072 65254 11124 65306
rect 11136 65254 11188 65306
rect 20811 65254 20863 65306
rect 20875 65254 20927 65306
rect 20939 65254 20991 65306
rect 21003 65254 21055 65306
rect 21067 65254 21119 65306
rect 13728 65152 13780 65204
rect 15292 65152 15344 65204
rect 17592 65152 17644 65204
rect 18696 65195 18748 65204
rect 18696 65161 18705 65195
rect 18705 65161 18739 65195
rect 18739 65161 18748 65195
rect 18696 65152 18748 65161
rect 17500 65127 17552 65136
rect 17500 65093 17509 65127
rect 17509 65093 17543 65127
rect 17543 65093 17552 65127
rect 17500 65084 17552 65093
rect 21272 65152 21324 65204
rect 21916 65152 21968 65204
rect 23204 65195 23256 65204
rect 23204 65161 23213 65195
rect 23213 65161 23247 65195
rect 23247 65161 23256 65195
rect 23204 65152 23256 65161
rect 27896 65152 27948 65204
rect 20444 65127 20496 65136
rect 20444 65093 20453 65127
rect 20453 65093 20487 65127
rect 20487 65093 20496 65127
rect 20444 65084 20496 65093
rect 20720 65084 20772 65136
rect 21824 65084 21876 65136
rect 12900 65059 12952 65068
rect 12900 65025 12909 65059
rect 12909 65025 12943 65059
rect 12943 65025 12952 65059
rect 12900 65016 12952 65025
rect 14004 65016 14056 65068
rect 15568 65016 15620 65068
rect 17132 65016 17184 65068
rect 18604 65016 18656 65068
rect 20260 65059 20312 65068
rect 20260 65025 20269 65059
rect 20269 65025 20303 65059
rect 20303 65025 20312 65059
rect 20260 65016 20312 65025
rect 14556 64948 14608 65000
rect 25504 65016 25556 65068
rect 23480 64948 23532 65000
rect 23756 64948 23808 65000
rect 28356 65016 28408 65068
rect 26148 64880 26200 64932
rect 28080 64948 28132 65000
rect 28908 64948 28960 65000
rect 30012 65016 30064 65068
rect 30380 65016 30432 65068
rect 29828 64948 29880 65000
rect 28356 64880 28408 64932
rect 12716 64855 12768 64864
rect 12716 64821 12725 64855
rect 12725 64821 12759 64855
rect 12759 64821 12768 64855
rect 12716 64812 12768 64821
rect 15476 64812 15528 64864
rect 21548 64812 21600 64864
rect 23388 64812 23440 64864
rect 30748 64812 30800 64864
rect 5915 64710 5967 64762
rect 5979 64710 6031 64762
rect 6043 64710 6095 64762
rect 6107 64710 6159 64762
rect 6171 64710 6223 64762
rect 15846 64710 15898 64762
rect 15910 64710 15962 64762
rect 15974 64710 16026 64762
rect 16038 64710 16090 64762
rect 16102 64710 16154 64762
rect 25776 64710 25828 64762
rect 25840 64710 25892 64762
rect 25904 64710 25956 64762
rect 25968 64710 26020 64762
rect 26032 64710 26084 64762
rect 19984 64608 20036 64660
rect 20076 64651 20128 64660
rect 20076 64617 20085 64651
rect 20085 64617 20119 64651
rect 20119 64617 20128 64651
rect 21180 64651 21232 64660
rect 20076 64608 20128 64617
rect 21180 64617 21189 64651
rect 21189 64617 21223 64651
rect 21223 64617 21232 64651
rect 21180 64608 21232 64617
rect 24860 64608 24912 64660
rect 25228 64608 25280 64660
rect 26332 64608 26384 64660
rect 21640 64540 21692 64592
rect 22376 64540 22428 64592
rect 31300 64608 31352 64660
rect 20352 64472 20404 64524
rect 1584 64447 1636 64456
rect 1584 64413 1593 64447
rect 1593 64413 1627 64447
rect 1627 64413 1636 64447
rect 1584 64404 1636 64413
rect 11244 64404 11296 64456
rect 19340 64404 19392 64456
rect 12716 64379 12768 64388
rect 12716 64345 12725 64379
rect 12725 64345 12759 64379
rect 12759 64345 12768 64379
rect 12716 64336 12768 64345
rect 20536 64336 20588 64388
rect 12164 64268 12216 64320
rect 15108 64268 15160 64320
rect 21640 64447 21692 64456
rect 21640 64413 21649 64447
rect 21649 64413 21683 64447
rect 21683 64413 21692 64447
rect 24400 64472 24452 64524
rect 21640 64404 21692 64413
rect 21916 64336 21968 64388
rect 22744 64404 22796 64456
rect 23480 64404 23532 64456
rect 24952 64404 25004 64456
rect 25136 64447 25188 64456
rect 25136 64413 25145 64447
rect 25145 64413 25179 64447
rect 25179 64413 25188 64447
rect 25136 64404 25188 64413
rect 25504 64404 25556 64456
rect 26148 64447 26200 64456
rect 26148 64413 26157 64447
rect 26157 64413 26191 64447
rect 26191 64413 26200 64447
rect 26148 64404 26200 64413
rect 26332 64404 26384 64456
rect 27068 64472 27120 64524
rect 27620 64472 27672 64524
rect 24492 64336 24544 64388
rect 24768 64336 24820 64388
rect 26516 64336 26568 64388
rect 24124 64268 24176 64320
rect 24676 64311 24728 64320
rect 24676 64277 24685 64311
rect 24685 64277 24719 64311
rect 24719 64277 24728 64311
rect 24676 64268 24728 64277
rect 25228 64268 25280 64320
rect 26976 64447 27028 64456
rect 26976 64413 26985 64447
rect 26985 64413 27019 64447
rect 27019 64413 27028 64447
rect 26976 64404 27028 64413
rect 27804 64447 27856 64456
rect 27804 64413 27813 64447
rect 27813 64413 27847 64447
rect 27847 64413 27856 64447
rect 27804 64404 27856 64413
rect 27896 64404 27948 64456
rect 31116 64404 31168 64456
rect 28908 64336 28960 64388
rect 28356 64268 28408 64320
rect 28632 64268 28684 64320
rect 29092 64268 29144 64320
rect 29828 64336 29880 64388
rect 30380 64336 30432 64388
rect 10880 64166 10932 64218
rect 10944 64166 10996 64218
rect 11008 64166 11060 64218
rect 11072 64166 11124 64218
rect 11136 64166 11188 64218
rect 20811 64166 20863 64218
rect 20875 64166 20927 64218
rect 20939 64166 20991 64218
rect 21003 64166 21055 64218
rect 21067 64166 21119 64218
rect 11336 64064 11388 64116
rect 12164 64039 12216 64048
rect 12164 64005 12173 64039
rect 12173 64005 12207 64039
rect 12207 64005 12216 64039
rect 12164 63996 12216 64005
rect 14648 63996 14700 64048
rect 20628 64064 20680 64116
rect 25504 64064 25556 64116
rect 25688 64064 25740 64116
rect 26792 64064 26844 64116
rect 20260 63996 20312 64048
rect 20720 64039 20772 64048
rect 20720 64005 20729 64039
rect 20729 64005 20763 64039
rect 20763 64005 20772 64039
rect 20720 63996 20772 64005
rect 24676 63996 24728 64048
rect 1584 63971 1636 63980
rect 1584 63937 1593 63971
rect 1593 63937 1627 63971
rect 1627 63937 1636 63971
rect 1584 63928 1636 63937
rect 12716 63928 12768 63980
rect 15568 63928 15620 63980
rect 17132 63971 17184 63980
rect 17132 63937 17141 63971
rect 17141 63937 17175 63971
rect 17175 63937 17184 63971
rect 17132 63928 17184 63937
rect 20536 63971 20588 63980
rect 20536 63937 20545 63971
rect 20545 63937 20579 63971
rect 20579 63937 20588 63971
rect 20536 63928 20588 63937
rect 22928 63928 22980 63980
rect 23204 63928 23256 63980
rect 23480 63928 23532 63980
rect 25136 63928 25188 63980
rect 27068 63928 27120 63980
rect 27528 63996 27580 64048
rect 27712 64064 27764 64116
rect 29460 64064 29512 64116
rect 28172 63971 28224 63980
rect 14556 63903 14608 63912
rect 14004 63835 14056 63844
rect 14004 63801 14013 63835
rect 14013 63801 14047 63835
rect 14047 63801 14056 63835
rect 14004 63792 14056 63801
rect 14556 63869 14565 63903
rect 14565 63869 14599 63903
rect 14599 63869 14608 63903
rect 14556 63860 14608 63869
rect 24032 63860 24084 63912
rect 25412 63860 25464 63912
rect 25688 63860 25740 63912
rect 28172 63937 28181 63971
rect 28181 63937 28215 63971
rect 28215 63937 28224 63971
rect 28172 63928 28224 63937
rect 28356 63971 28408 63980
rect 28356 63937 28365 63971
rect 28365 63937 28399 63971
rect 28399 63937 28408 63971
rect 29092 63996 29144 64048
rect 28356 63928 28408 63937
rect 28080 63860 28132 63912
rect 29460 63928 29512 63980
rect 30012 63928 30064 63980
rect 17960 63792 18012 63844
rect 27712 63792 27764 63844
rect 11336 63724 11388 63776
rect 13912 63724 13964 63776
rect 24124 63724 24176 63776
rect 28264 63792 28316 63844
rect 28816 63792 28868 63844
rect 30748 63860 30800 63912
rect 31668 63860 31720 63912
rect 5915 63622 5967 63674
rect 5979 63622 6031 63674
rect 6043 63622 6095 63674
rect 6107 63622 6159 63674
rect 6171 63622 6223 63674
rect 15846 63622 15898 63674
rect 15910 63622 15962 63674
rect 15974 63622 16026 63674
rect 16038 63622 16090 63674
rect 16102 63622 16154 63674
rect 25776 63622 25828 63674
rect 25840 63622 25892 63674
rect 25904 63622 25956 63674
rect 25968 63622 26020 63674
rect 26032 63622 26084 63674
rect 23388 63520 23440 63572
rect 23664 63520 23716 63572
rect 27712 63520 27764 63572
rect 13820 63452 13872 63504
rect 15568 63495 15620 63504
rect 15568 63461 15577 63495
rect 15577 63461 15611 63495
rect 15611 63461 15620 63495
rect 15568 63452 15620 63461
rect 17776 63452 17828 63504
rect 20352 63452 20404 63504
rect 23572 63452 23624 63504
rect 28080 63452 28132 63504
rect 28264 63452 28316 63504
rect 1584 63359 1636 63368
rect 1584 63325 1593 63359
rect 1593 63325 1627 63359
rect 1627 63325 1636 63359
rect 1584 63316 1636 63325
rect 11428 63248 11480 63300
rect 13820 63316 13872 63368
rect 14188 63316 14240 63368
rect 20260 63427 20312 63436
rect 20260 63393 20269 63427
rect 20269 63393 20303 63427
rect 20303 63393 20312 63427
rect 20260 63384 20312 63393
rect 20720 63384 20772 63436
rect 23664 63384 23716 63436
rect 24584 63427 24636 63436
rect 24584 63393 24593 63427
rect 24593 63393 24627 63427
rect 24627 63393 24636 63427
rect 24584 63384 24636 63393
rect 28540 63520 28592 63572
rect 28540 63427 28592 63436
rect 15568 63316 15620 63368
rect 23848 63316 23900 63368
rect 24952 63316 25004 63368
rect 25412 63316 25464 63368
rect 12716 63248 12768 63300
rect 14556 63248 14608 63300
rect 15384 63291 15436 63300
rect 15384 63257 15393 63291
rect 15393 63257 15427 63291
rect 15427 63257 15436 63291
rect 15384 63248 15436 63257
rect 16580 63291 16632 63300
rect 16580 63257 16589 63291
rect 16589 63257 16623 63291
rect 16623 63257 16632 63291
rect 16580 63248 16632 63257
rect 11244 63180 11296 63232
rect 14648 63223 14700 63232
rect 14648 63189 14657 63223
rect 14657 63189 14691 63223
rect 14691 63189 14700 63223
rect 14648 63180 14700 63189
rect 15016 63180 15068 63232
rect 23940 63248 23992 63300
rect 24584 63248 24636 63300
rect 27712 63316 27764 63368
rect 27620 63248 27672 63300
rect 21272 63180 21324 63232
rect 25412 63180 25464 63232
rect 26148 63180 26200 63232
rect 26792 63180 26844 63232
rect 28540 63393 28543 63427
rect 28543 63393 28577 63427
rect 28577 63393 28592 63427
rect 28540 63384 28592 63393
rect 28264 63359 28316 63368
rect 28264 63325 28273 63359
rect 28273 63325 28307 63359
rect 28307 63325 28316 63359
rect 28264 63316 28316 63325
rect 28356 63316 28408 63368
rect 30564 63384 30616 63436
rect 28540 63248 28592 63300
rect 29092 63316 29144 63368
rect 29828 63359 29880 63368
rect 29828 63325 29837 63359
rect 29837 63325 29871 63359
rect 29871 63325 29880 63359
rect 29828 63316 29880 63325
rect 29276 63248 29328 63300
rect 29736 63248 29788 63300
rect 30380 63248 30432 63300
rect 30564 63248 30616 63300
rect 29552 63180 29604 63232
rect 10880 63078 10932 63130
rect 10944 63078 10996 63130
rect 11008 63078 11060 63130
rect 11072 63078 11124 63130
rect 11136 63078 11188 63130
rect 20811 63078 20863 63130
rect 20875 63078 20927 63130
rect 20939 63078 20991 63130
rect 21003 63078 21055 63130
rect 21067 63078 21119 63130
rect 11336 62908 11388 62960
rect 17868 62976 17920 63028
rect 1584 62883 1636 62892
rect 1584 62849 1593 62883
rect 1593 62849 1627 62883
rect 1627 62849 1636 62883
rect 1584 62840 1636 62849
rect 12716 62840 12768 62892
rect 17408 62840 17460 62892
rect 17224 62772 17276 62824
rect 17868 62883 17920 62892
rect 17868 62849 17877 62883
rect 17877 62849 17911 62883
rect 17911 62849 17920 62883
rect 17868 62840 17920 62849
rect 19432 62840 19484 62892
rect 20352 62883 20404 62892
rect 20352 62849 20361 62883
rect 20361 62849 20395 62883
rect 20395 62849 20404 62883
rect 20352 62840 20404 62849
rect 23848 62840 23900 62892
rect 18420 62772 18472 62824
rect 24584 62772 24636 62824
rect 26976 62976 27028 63028
rect 28632 62976 28684 63028
rect 29184 62976 29236 63028
rect 27620 62840 27672 62892
rect 28908 62908 28960 62960
rect 15200 62704 15252 62756
rect 17316 62704 17368 62756
rect 26516 62772 26568 62824
rect 28540 62840 28592 62892
rect 28632 62772 28684 62824
rect 11336 62636 11388 62688
rect 15108 62636 15160 62688
rect 16488 62636 16540 62688
rect 17408 62636 17460 62688
rect 19984 62636 20036 62688
rect 21088 62636 21140 62688
rect 24032 62636 24084 62688
rect 27160 62679 27212 62688
rect 27160 62645 27169 62679
rect 27169 62645 27203 62679
rect 27203 62645 27212 62679
rect 27160 62636 27212 62645
rect 27344 62636 27396 62688
rect 28080 62704 28132 62756
rect 28540 62704 28592 62756
rect 29368 62883 29420 62892
rect 29368 62849 29377 62883
rect 29377 62849 29411 62883
rect 29411 62849 29420 62883
rect 29368 62840 29420 62849
rect 29184 62772 29236 62824
rect 30012 62840 30064 62892
rect 5915 62534 5967 62586
rect 5979 62534 6031 62586
rect 6043 62534 6095 62586
rect 6107 62534 6159 62586
rect 6171 62534 6223 62586
rect 15846 62534 15898 62586
rect 15910 62534 15962 62586
rect 15974 62534 16026 62586
rect 16038 62534 16090 62586
rect 16102 62534 16154 62586
rect 25776 62534 25828 62586
rect 25840 62534 25892 62586
rect 25904 62534 25956 62586
rect 25968 62534 26020 62586
rect 26032 62534 26084 62586
rect 18328 62432 18380 62484
rect 24400 62432 24452 62484
rect 28356 62432 28408 62484
rect 29460 62432 29512 62484
rect 16028 62364 16080 62416
rect 16028 62228 16080 62280
rect 16212 62271 16264 62280
rect 16212 62237 16221 62271
rect 16221 62237 16255 62271
rect 16255 62237 16264 62271
rect 16212 62228 16264 62237
rect 16856 62296 16908 62348
rect 21088 62339 21140 62348
rect 21088 62305 21097 62339
rect 21097 62305 21131 62339
rect 21131 62305 21140 62339
rect 21088 62296 21140 62305
rect 22100 62296 22152 62348
rect 24952 62364 25004 62416
rect 16488 62271 16540 62280
rect 16488 62237 16497 62271
rect 16497 62237 16531 62271
rect 16531 62237 16540 62271
rect 17316 62271 17368 62280
rect 16488 62228 16540 62237
rect 17316 62237 17325 62271
rect 17325 62237 17359 62271
rect 17359 62237 17368 62271
rect 17316 62228 17368 62237
rect 17408 62228 17460 62280
rect 23480 62271 23532 62280
rect 23480 62237 23489 62271
rect 23489 62237 23523 62271
rect 23523 62237 23532 62271
rect 23480 62228 23532 62237
rect 26148 62296 26200 62348
rect 24860 62271 24912 62280
rect 24860 62237 24869 62271
rect 24869 62237 24903 62271
rect 24903 62237 24912 62271
rect 24860 62228 24912 62237
rect 25228 62228 25280 62280
rect 26976 62228 27028 62280
rect 27252 62271 27304 62280
rect 27252 62237 27261 62271
rect 27261 62237 27295 62271
rect 27295 62237 27304 62271
rect 27252 62228 27304 62237
rect 27712 62296 27764 62348
rect 28632 62296 28684 62348
rect 29276 62296 29328 62348
rect 29460 62296 29512 62348
rect 27436 62228 27488 62280
rect 16764 62160 16816 62212
rect 21824 62160 21876 62212
rect 28632 62203 28684 62212
rect 14648 62092 14700 62144
rect 16672 62092 16724 62144
rect 17500 62092 17552 62144
rect 18696 62135 18748 62144
rect 18696 62101 18705 62135
rect 18705 62101 18739 62135
rect 18739 62101 18748 62135
rect 18696 62092 18748 62101
rect 18880 62092 18932 62144
rect 28632 62169 28641 62203
rect 28641 62169 28675 62203
rect 28675 62169 28684 62203
rect 28632 62160 28684 62169
rect 29092 62228 29144 62280
rect 30012 62271 30064 62280
rect 30012 62237 30021 62271
rect 30021 62237 30055 62271
rect 30055 62237 30064 62271
rect 30012 62228 30064 62237
rect 25964 62092 26016 62144
rect 26424 62092 26476 62144
rect 27896 62092 27948 62144
rect 10880 61990 10932 62042
rect 10944 61990 10996 62042
rect 11008 61990 11060 62042
rect 11072 61990 11124 62042
rect 11136 61990 11188 62042
rect 20811 61990 20863 62042
rect 20875 61990 20927 62042
rect 20939 61990 20991 62042
rect 21003 61990 21055 62042
rect 21067 61990 21119 62042
rect 14096 61888 14148 61940
rect 11244 61820 11296 61872
rect 1584 61795 1636 61804
rect 1584 61761 1593 61795
rect 1593 61761 1627 61795
rect 1627 61761 1636 61795
rect 1584 61752 1636 61761
rect 12532 61795 12584 61804
rect 12532 61761 12541 61795
rect 12541 61761 12575 61795
rect 12575 61761 12584 61795
rect 12532 61752 12584 61761
rect 15200 61795 15252 61804
rect 15200 61761 15209 61795
rect 15209 61761 15243 61795
rect 15243 61761 15252 61795
rect 15200 61752 15252 61761
rect 16856 61888 16908 61940
rect 21824 61931 21876 61940
rect 21824 61897 21833 61931
rect 21833 61897 21867 61931
rect 21867 61897 21876 61931
rect 21824 61888 21876 61897
rect 24768 61888 24820 61940
rect 25044 61931 25096 61940
rect 25044 61897 25053 61931
rect 25053 61897 25087 61931
rect 25087 61897 25096 61931
rect 25044 61888 25096 61897
rect 25688 61931 25740 61940
rect 25688 61897 25697 61931
rect 25697 61897 25731 61931
rect 25731 61897 25740 61931
rect 25688 61888 25740 61897
rect 15568 61795 15620 61804
rect 15568 61761 15577 61795
rect 15577 61761 15611 61795
rect 15611 61761 15620 61795
rect 15568 61752 15620 61761
rect 16580 61752 16632 61804
rect 19708 61820 19760 61872
rect 21180 61820 21232 61872
rect 18788 61795 18840 61804
rect 18788 61761 18822 61795
rect 18822 61761 18840 61795
rect 22100 61795 22152 61804
rect 18788 61752 18840 61761
rect 22100 61761 22109 61795
rect 22109 61761 22143 61795
rect 22143 61761 22152 61795
rect 22100 61752 22152 61761
rect 22376 61820 22428 61872
rect 22468 61795 22520 61804
rect 16212 61684 16264 61736
rect 17224 61684 17276 61736
rect 17500 61684 17552 61736
rect 18512 61727 18564 61736
rect 18512 61693 18521 61727
rect 18521 61693 18555 61727
rect 18555 61693 18564 61727
rect 18512 61684 18564 61693
rect 22008 61684 22060 61736
rect 22468 61761 22477 61795
rect 22477 61761 22511 61795
rect 22511 61761 22520 61795
rect 22468 61752 22520 61761
rect 23848 61752 23900 61804
rect 24124 61795 24176 61804
rect 24124 61761 24133 61795
rect 24133 61761 24167 61795
rect 24167 61761 24176 61795
rect 24124 61752 24176 61761
rect 24492 61752 24544 61804
rect 24860 61795 24912 61804
rect 24860 61761 24869 61795
rect 24869 61761 24903 61795
rect 24903 61761 24912 61795
rect 25964 61820 26016 61872
rect 24860 61752 24912 61761
rect 25228 61752 25280 61804
rect 25688 61752 25740 61804
rect 26332 61752 26384 61804
rect 26976 61752 27028 61804
rect 27344 61761 27353 61788
rect 27353 61761 27387 61788
rect 27387 61761 27396 61788
rect 27344 61736 27396 61761
rect 27528 61752 27580 61804
rect 30656 61820 30708 61872
rect 28356 61752 28408 61804
rect 28724 61752 28776 61804
rect 29184 61795 29236 61804
rect 29184 61761 29193 61795
rect 29193 61761 29227 61795
rect 29227 61761 29236 61795
rect 29184 61752 29236 61761
rect 7564 61548 7616 61600
rect 14740 61548 14792 61600
rect 14924 61591 14976 61600
rect 14924 61557 14933 61591
rect 14933 61557 14967 61591
rect 14967 61557 14976 61591
rect 14924 61548 14976 61557
rect 19156 61548 19208 61600
rect 22836 61548 22888 61600
rect 23480 61548 23532 61600
rect 27896 61616 27948 61668
rect 24952 61548 25004 61600
rect 25044 61548 25096 61600
rect 25412 61548 25464 61600
rect 27436 61548 27488 61600
rect 28724 61616 28776 61668
rect 28816 61548 28868 61600
rect 5915 61446 5967 61498
rect 5979 61446 6031 61498
rect 6043 61446 6095 61498
rect 6107 61446 6159 61498
rect 6171 61446 6223 61498
rect 15846 61446 15898 61498
rect 15910 61446 15962 61498
rect 15974 61446 16026 61498
rect 16038 61446 16090 61498
rect 16102 61446 16154 61498
rect 25776 61446 25828 61498
rect 25840 61446 25892 61498
rect 25904 61446 25956 61498
rect 25968 61446 26020 61498
rect 26032 61446 26084 61498
rect 15384 61344 15436 61396
rect 16396 61387 16448 61396
rect 16396 61353 16405 61387
rect 16405 61353 16439 61387
rect 16439 61353 16448 61387
rect 16396 61344 16448 61353
rect 18512 61344 18564 61396
rect 24676 61344 24728 61396
rect 25412 61344 25464 61396
rect 20168 61276 20220 61328
rect 27436 61344 27488 61396
rect 29736 61344 29788 61396
rect 28816 61276 28868 61328
rect 29092 61276 29144 61328
rect 29276 61276 29328 61328
rect 29368 61276 29420 61328
rect 7564 61208 7616 61260
rect 1584 61183 1636 61192
rect 1584 61149 1593 61183
rect 1593 61149 1627 61183
rect 1627 61149 1636 61183
rect 1584 61140 1636 61149
rect 12900 61183 12952 61192
rect 12900 61149 12909 61183
rect 12909 61149 12943 61183
rect 12943 61149 12952 61183
rect 12900 61140 12952 61149
rect 13452 61140 13504 61192
rect 15200 61208 15252 61260
rect 15660 61208 15712 61260
rect 16856 61208 16908 61260
rect 17408 61140 17460 61192
rect 18328 61208 18380 61260
rect 23940 61208 23992 61260
rect 24860 61208 24912 61260
rect 17960 61183 18012 61192
rect 17960 61149 17969 61183
rect 17969 61149 18003 61183
rect 18003 61149 18012 61183
rect 18512 61183 18564 61192
rect 17960 61140 18012 61149
rect 18512 61149 18521 61183
rect 18521 61149 18555 61183
rect 18555 61149 18564 61183
rect 18512 61140 18564 61149
rect 19708 61183 19760 61192
rect 19708 61149 19717 61183
rect 19717 61149 19751 61183
rect 19751 61149 19760 61183
rect 19708 61140 19760 61149
rect 20260 61140 20312 61192
rect 22376 61140 22428 61192
rect 23480 61183 23532 61192
rect 23480 61149 23489 61183
rect 23489 61149 23523 61183
rect 23523 61149 23532 61183
rect 23480 61140 23532 61149
rect 25228 61140 25280 61192
rect 25688 61140 25740 61192
rect 25964 61140 26016 61192
rect 26332 61183 26384 61192
rect 26332 61149 26341 61183
rect 26341 61149 26375 61183
rect 26375 61149 26384 61183
rect 26332 61140 26384 61149
rect 26976 61140 27028 61192
rect 11244 61004 11296 61056
rect 12532 61004 12584 61056
rect 16212 61072 16264 61124
rect 17500 61072 17552 61124
rect 24860 61072 24912 61124
rect 25596 61072 25648 61124
rect 25780 61072 25832 61124
rect 28632 61208 28684 61260
rect 27896 61183 27948 61192
rect 27896 61149 27905 61183
rect 27905 61149 27939 61183
rect 27939 61149 27948 61183
rect 27896 61140 27948 61149
rect 28448 61140 28500 61192
rect 28816 61140 28868 61192
rect 29092 61140 29144 61192
rect 30012 61183 30064 61192
rect 30012 61149 30021 61183
rect 30021 61149 30055 61183
rect 30055 61149 30064 61183
rect 30012 61140 30064 61149
rect 16948 61004 17000 61056
rect 19708 61004 19760 61056
rect 23480 61004 23532 61056
rect 24584 61004 24636 61056
rect 25320 61004 25372 61056
rect 25504 61004 25556 61056
rect 25688 61004 25740 61056
rect 26240 61047 26292 61056
rect 26240 61013 26249 61047
rect 26249 61013 26283 61047
rect 26283 61013 26292 61047
rect 26240 61004 26292 61013
rect 29092 61004 29144 61056
rect 30104 61004 30156 61056
rect 10880 60902 10932 60954
rect 10944 60902 10996 60954
rect 11008 60902 11060 60954
rect 11072 60902 11124 60954
rect 11136 60902 11188 60954
rect 20811 60902 20863 60954
rect 20875 60902 20927 60954
rect 20939 60902 20991 60954
rect 21003 60902 21055 60954
rect 21067 60902 21119 60954
rect 12532 60775 12584 60784
rect 12532 60741 12541 60775
rect 12541 60741 12575 60775
rect 12575 60741 12584 60775
rect 12532 60732 12584 60741
rect 1584 60707 1636 60716
rect 1584 60673 1593 60707
rect 1593 60673 1627 60707
rect 1627 60673 1636 60707
rect 1584 60664 1636 60673
rect 11336 60596 11388 60648
rect 13636 60707 13688 60716
rect 13636 60673 13645 60707
rect 13645 60673 13679 60707
rect 13679 60673 13688 60707
rect 13636 60664 13688 60673
rect 16120 60800 16172 60852
rect 18328 60843 18380 60852
rect 18328 60809 18337 60843
rect 18337 60809 18371 60843
rect 18371 60809 18380 60843
rect 18328 60800 18380 60809
rect 18788 60800 18840 60852
rect 17868 60732 17920 60784
rect 18972 60732 19024 60784
rect 14004 60707 14056 60716
rect 14004 60673 14013 60707
rect 14013 60673 14047 60707
rect 14047 60673 14056 60707
rect 14004 60664 14056 60673
rect 14004 60528 14056 60580
rect 12716 60460 12768 60512
rect 12900 60503 12952 60512
rect 12900 60469 12909 60503
rect 12909 60469 12943 60503
rect 12943 60469 12952 60503
rect 12900 60460 12952 60469
rect 16672 60664 16724 60716
rect 19064 60664 19116 60716
rect 19708 60800 19760 60852
rect 24124 60800 24176 60852
rect 24676 60800 24728 60852
rect 25872 60800 25924 60852
rect 14280 60596 14332 60648
rect 16856 60596 16908 60648
rect 18420 60596 18472 60648
rect 19616 60664 19668 60716
rect 20812 60664 20864 60716
rect 22008 60732 22060 60784
rect 22652 60732 22704 60784
rect 27528 60800 27580 60852
rect 27804 60800 27856 60852
rect 21180 60664 21232 60716
rect 21548 60664 21600 60716
rect 22836 60707 22888 60716
rect 22836 60673 22845 60707
rect 22845 60673 22879 60707
rect 22879 60673 22888 60707
rect 22836 60664 22888 60673
rect 23112 60664 23164 60716
rect 24952 60664 25004 60716
rect 25228 60664 25280 60716
rect 25320 60664 25372 60716
rect 25780 60670 25832 60722
rect 19800 60596 19852 60648
rect 14740 60460 14792 60512
rect 15752 60460 15804 60512
rect 18696 60528 18748 60580
rect 25504 60596 25556 60648
rect 27068 60664 27120 60716
rect 27436 60707 27488 60716
rect 24400 60528 24452 60580
rect 26792 60596 26844 60648
rect 27436 60673 27445 60707
rect 27445 60673 27479 60707
rect 27479 60673 27488 60707
rect 27436 60664 27488 60673
rect 28632 60800 28684 60852
rect 29460 60732 29512 60784
rect 29736 60775 29788 60784
rect 29736 60741 29745 60775
rect 29745 60741 29779 60775
rect 29779 60741 29788 60775
rect 29736 60732 29788 60741
rect 28908 60707 28960 60716
rect 19616 60460 19668 60512
rect 20628 60503 20680 60512
rect 20628 60469 20637 60503
rect 20637 60469 20671 60503
rect 20671 60469 20680 60503
rect 20628 60460 20680 60469
rect 22100 60460 22152 60512
rect 23572 60460 23624 60512
rect 26148 60528 26200 60580
rect 26332 60528 26384 60580
rect 27068 60528 27120 60580
rect 28908 60673 28917 60707
rect 28917 60673 28951 60707
rect 28951 60673 28960 60707
rect 28908 60664 28960 60673
rect 29092 60664 29144 60716
rect 29368 60596 29420 60648
rect 29460 60596 29512 60648
rect 30932 60596 30984 60648
rect 27344 60460 27396 60512
rect 28356 60460 28408 60512
rect 29736 60460 29788 60512
rect 29828 60503 29880 60512
rect 29828 60469 29837 60503
rect 29837 60469 29871 60503
rect 29871 60469 29880 60503
rect 29828 60460 29880 60469
rect 5915 60358 5967 60410
rect 5979 60358 6031 60410
rect 6043 60358 6095 60410
rect 6107 60358 6159 60410
rect 6171 60358 6223 60410
rect 15846 60358 15898 60410
rect 15910 60358 15962 60410
rect 15974 60358 16026 60410
rect 16038 60358 16090 60410
rect 16102 60358 16154 60410
rect 25776 60358 25828 60410
rect 25840 60358 25892 60410
rect 25904 60358 25956 60410
rect 25968 60358 26020 60410
rect 26032 60358 26084 60410
rect 13636 60256 13688 60308
rect 15752 60256 15804 60308
rect 17316 60256 17368 60308
rect 21732 60256 21784 60308
rect 22376 60299 22428 60308
rect 14096 60188 14148 60240
rect 19340 60120 19392 60172
rect 20352 60120 20404 60172
rect 20536 60120 20588 60172
rect 22376 60265 22385 60299
rect 22385 60265 22419 60299
rect 22419 60265 22428 60299
rect 22376 60256 22428 60265
rect 23940 60256 23992 60308
rect 25320 60256 25372 60308
rect 26608 60256 26660 60308
rect 26700 60256 26752 60308
rect 23480 60188 23532 60240
rect 27160 60188 27212 60240
rect 25872 60120 25924 60172
rect 1584 60095 1636 60104
rect 1584 60061 1593 60095
rect 1593 60061 1627 60095
rect 1627 60061 1636 60095
rect 1584 60052 1636 60061
rect 11244 60052 11296 60104
rect 12532 60095 12584 60104
rect 12532 60061 12541 60095
rect 12541 60061 12575 60095
rect 12575 60061 12584 60095
rect 17684 60095 17736 60104
rect 12532 60052 12584 60061
rect 17684 60061 17693 60095
rect 17693 60061 17727 60095
rect 17727 60061 17736 60095
rect 17684 60052 17736 60061
rect 19616 60095 19668 60104
rect 14464 60027 14516 60036
rect 14464 59993 14473 60027
rect 14473 59993 14507 60027
rect 14507 59993 14516 60027
rect 14464 59984 14516 59993
rect 14648 60027 14700 60036
rect 14648 59993 14657 60027
rect 14657 59993 14691 60027
rect 14691 59993 14700 60027
rect 14648 59984 14700 59993
rect 14740 60027 14792 60036
rect 14740 59993 14749 60027
rect 14749 59993 14783 60027
rect 14783 59993 14792 60027
rect 15476 60027 15528 60036
rect 14740 59984 14792 59993
rect 15476 59993 15485 60027
rect 15485 59993 15519 60027
rect 15519 59993 15528 60027
rect 15476 59984 15528 59993
rect 15752 59984 15804 60036
rect 18972 59984 19024 60036
rect 19616 60061 19625 60095
rect 19625 60061 19659 60095
rect 19659 60061 19668 60095
rect 19616 60052 19668 60061
rect 19800 60052 19852 60104
rect 19892 60095 19944 60104
rect 19892 60061 19901 60095
rect 19901 60061 19935 60095
rect 19935 60061 19944 60095
rect 19892 60052 19944 60061
rect 23204 60052 23256 60104
rect 25780 60095 25832 60104
rect 25780 60061 25789 60095
rect 25789 60061 25823 60095
rect 25823 60061 25832 60095
rect 25780 60052 25832 60061
rect 26332 60052 26384 60104
rect 26608 60052 26660 60104
rect 27160 60052 27212 60104
rect 27804 60095 27856 60104
rect 27804 60061 27813 60095
rect 27813 60061 27847 60095
rect 27847 60061 27856 60095
rect 27804 60052 27856 60061
rect 28356 60095 28408 60104
rect 20536 59984 20588 60036
rect 20628 59984 20680 60036
rect 21456 59984 21508 60036
rect 21916 59984 21968 60036
rect 28080 59984 28132 60036
rect 28356 60061 28365 60095
rect 28365 60061 28399 60095
rect 28399 60061 28408 60095
rect 28356 60052 28408 60061
rect 29920 60052 29972 60104
rect 11336 59916 11388 59968
rect 16672 59916 16724 59968
rect 19156 59916 19208 59968
rect 23296 59959 23348 59968
rect 23296 59925 23305 59959
rect 23305 59925 23339 59959
rect 23339 59925 23348 59959
rect 23296 59916 23348 59925
rect 26608 59916 26660 59968
rect 26792 59916 26844 59968
rect 28356 59916 28408 59968
rect 28632 59916 28684 59968
rect 29460 59916 29512 59968
rect 10880 59814 10932 59866
rect 10944 59814 10996 59866
rect 11008 59814 11060 59866
rect 11072 59814 11124 59866
rect 11136 59814 11188 59866
rect 20811 59814 20863 59866
rect 20875 59814 20927 59866
rect 20939 59814 20991 59866
rect 21003 59814 21055 59866
rect 21067 59814 21119 59866
rect 13544 59755 13596 59764
rect 13544 59721 13553 59755
rect 13553 59721 13587 59755
rect 13587 59721 13596 59755
rect 13544 59712 13596 59721
rect 14280 59755 14332 59764
rect 14280 59721 14289 59755
rect 14289 59721 14323 59755
rect 14323 59721 14332 59755
rect 14280 59712 14332 59721
rect 16856 59755 16908 59764
rect 16856 59721 16865 59755
rect 16865 59721 16899 59755
rect 16899 59721 16908 59755
rect 16856 59712 16908 59721
rect 12532 59687 12584 59696
rect 12532 59653 12541 59687
rect 12541 59653 12575 59687
rect 12575 59653 12584 59687
rect 12532 59644 12584 59653
rect 12716 59687 12768 59696
rect 12716 59653 12725 59687
rect 12725 59653 12759 59687
rect 12759 59653 12768 59687
rect 12716 59644 12768 59653
rect 16304 59644 16356 59696
rect 19156 59644 19208 59696
rect 1584 59619 1636 59628
rect 1584 59585 1593 59619
rect 1593 59585 1627 59619
rect 1627 59585 1636 59619
rect 1584 59576 1636 59585
rect 13452 59619 13504 59628
rect 13452 59585 13461 59619
rect 13461 59585 13495 59619
rect 13495 59585 13504 59619
rect 13452 59576 13504 59585
rect 14096 59619 14148 59628
rect 14096 59585 14105 59619
rect 14105 59585 14139 59619
rect 14139 59585 14148 59619
rect 14096 59576 14148 59585
rect 16764 59576 16816 59628
rect 19064 59576 19116 59628
rect 12900 59508 12952 59560
rect 19892 59576 19944 59628
rect 23112 59619 23164 59628
rect 23112 59585 23121 59619
rect 23121 59585 23155 59619
rect 23155 59585 23164 59619
rect 23112 59576 23164 59585
rect 23940 59576 23992 59628
rect 23020 59508 23072 59560
rect 23480 59508 23532 59560
rect 11244 59372 11296 59424
rect 18880 59440 18932 59492
rect 20536 59440 20588 59492
rect 25872 59712 25924 59764
rect 26884 59712 26936 59764
rect 25228 59644 25280 59696
rect 26332 59576 26384 59628
rect 27160 59576 27212 59628
rect 27344 59576 27396 59628
rect 27712 59619 27764 59628
rect 27712 59585 27721 59619
rect 27721 59585 27755 59619
rect 27755 59585 27764 59619
rect 27712 59576 27764 59585
rect 31024 59644 31076 59696
rect 28080 59619 28132 59628
rect 26884 59508 26936 59560
rect 28080 59585 28089 59619
rect 28089 59585 28123 59619
rect 28123 59585 28132 59619
rect 28080 59576 28132 59585
rect 29828 59576 29880 59628
rect 28724 59508 28776 59560
rect 25228 59440 25280 59492
rect 25780 59440 25832 59492
rect 26976 59440 27028 59492
rect 14832 59372 14884 59424
rect 21732 59372 21784 59424
rect 23204 59372 23256 59424
rect 27344 59372 27396 59424
rect 30748 59440 30800 59492
rect 5915 59270 5967 59322
rect 5979 59270 6031 59322
rect 6043 59270 6095 59322
rect 6107 59270 6159 59322
rect 6171 59270 6223 59322
rect 15846 59270 15898 59322
rect 15910 59270 15962 59322
rect 15974 59270 16026 59322
rect 16038 59270 16090 59322
rect 16102 59270 16154 59322
rect 25776 59270 25828 59322
rect 25840 59270 25892 59322
rect 25904 59270 25956 59322
rect 25968 59270 26020 59322
rect 26032 59270 26084 59322
rect 18604 59168 18656 59220
rect 20260 59168 20312 59220
rect 20536 59168 20588 59220
rect 21364 59168 21416 59220
rect 23388 59168 23440 59220
rect 21824 59100 21876 59152
rect 28632 59168 28684 59220
rect 29736 59168 29788 59220
rect 30380 59168 30432 59220
rect 30656 59100 30708 59152
rect 27436 59032 27488 59084
rect 11336 58964 11388 59016
rect 13544 58964 13596 59016
rect 16396 58964 16448 59016
rect 20536 58964 20588 59016
rect 13176 58939 13228 58948
rect 13176 58905 13185 58939
rect 13185 58905 13219 58939
rect 13219 58905 13228 58939
rect 29368 58964 29420 59016
rect 13176 58896 13228 58905
rect 18328 58896 18380 58948
rect 20168 58896 20220 58948
rect 23848 58896 23900 58948
rect 24400 58896 24452 58948
rect 27436 58896 27488 58948
rect 28632 58939 28684 58948
rect 28632 58905 28641 58939
rect 28641 58905 28675 58939
rect 28675 58905 28684 58939
rect 28632 58896 28684 58905
rect 29736 58939 29788 58948
rect 29736 58905 29745 58939
rect 29745 58905 29779 58939
rect 29779 58905 29788 58939
rect 29736 58896 29788 58905
rect 30104 58939 30156 58948
rect 30104 58905 30113 58939
rect 30113 58905 30147 58939
rect 30147 58905 30156 58939
rect 30104 58896 30156 58905
rect 14464 58828 14516 58880
rect 17224 58828 17276 58880
rect 10880 58726 10932 58778
rect 10944 58726 10996 58778
rect 11008 58726 11060 58778
rect 11072 58726 11124 58778
rect 11136 58726 11188 58778
rect 20811 58726 20863 58778
rect 20875 58726 20927 58778
rect 20939 58726 20991 58778
rect 21003 58726 21055 58778
rect 21067 58726 21119 58778
rect 19156 58624 19208 58676
rect 27620 58624 27672 58676
rect 27712 58624 27764 58676
rect 11244 58556 11296 58608
rect 16672 58556 16724 58608
rect 17592 58556 17644 58608
rect 19248 58556 19300 58608
rect 21180 58556 21232 58608
rect 21640 58556 21692 58608
rect 26332 58556 26384 58608
rect 1400 58531 1452 58540
rect 1400 58497 1409 58531
rect 1409 58497 1443 58531
rect 1443 58497 1452 58531
rect 1400 58488 1452 58497
rect 13176 58531 13228 58540
rect 13176 58497 13185 58531
rect 13185 58497 13219 58531
rect 13219 58497 13228 58531
rect 13176 58488 13228 58497
rect 19524 58531 19576 58540
rect 17224 58463 17276 58472
rect 17224 58429 17233 58463
rect 17233 58429 17267 58463
rect 17267 58429 17276 58463
rect 17224 58420 17276 58429
rect 17316 58463 17368 58472
rect 17316 58429 17325 58463
rect 17325 58429 17359 58463
rect 17359 58429 17368 58463
rect 19524 58497 19533 58531
rect 19533 58497 19567 58531
rect 19567 58497 19576 58531
rect 19524 58488 19576 58497
rect 20076 58488 20128 58540
rect 20352 58488 20404 58540
rect 23664 58488 23716 58540
rect 24400 58488 24452 58540
rect 26976 58488 27028 58540
rect 27344 58488 27396 58540
rect 28632 58624 28684 58676
rect 30012 58624 30064 58676
rect 29092 58556 29144 58608
rect 17316 58420 17368 58429
rect 21180 58420 21232 58472
rect 1584 58395 1636 58404
rect 1584 58361 1593 58395
rect 1593 58361 1627 58395
rect 1627 58361 1636 58395
rect 1584 58352 1636 58361
rect 16488 58352 16540 58404
rect 16764 58395 16816 58404
rect 16764 58361 16773 58395
rect 16773 58361 16807 58395
rect 16807 58361 16816 58395
rect 16764 58352 16816 58361
rect 26332 58352 26384 58404
rect 28632 58531 28684 58540
rect 13544 58327 13596 58336
rect 13544 58293 13553 58327
rect 13553 58293 13587 58327
rect 13587 58293 13596 58327
rect 13544 58284 13596 58293
rect 26976 58284 27028 58336
rect 28632 58497 28641 58531
rect 28641 58497 28675 58531
rect 28675 58497 28684 58531
rect 28632 58488 28684 58497
rect 29368 58531 29420 58540
rect 29368 58497 29377 58531
rect 29377 58497 29411 58531
rect 29411 58497 29420 58531
rect 29368 58488 29420 58497
rect 30656 58556 30708 58608
rect 31208 58556 31260 58608
rect 30012 58488 30064 58540
rect 30380 58488 30432 58540
rect 31484 58420 31536 58472
rect 30380 58352 30432 58404
rect 29828 58284 29880 58336
rect 30104 58284 30156 58336
rect 5915 58182 5967 58234
rect 5979 58182 6031 58234
rect 6043 58182 6095 58234
rect 6107 58182 6159 58234
rect 6171 58182 6223 58234
rect 15846 58182 15898 58234
rect 15910 58182 15962 58234
rect 15974 58182 16026 58234
rect 16038 58182 16090 58234
rect 16102 58182 16154 58234
rect 25776 58182 25828 58234
rect 25840 58182 25892 58234
rect 25904 58182 25956 58234
rect 25968 58182 26020 58234
rect 26032 58182 26084 58234
rect 18512 58080 18564 58132
rect 13544 58012 13596 58064
rect 21548 58012 21600 58064
rect 25872 58012 25924 58064
rect 27160 58012 27212 58064
rect 15108 57944 15160 57996
rect 17868 57944 17920 57996
rect 23020 57944 23072 57996
rect 23664 57944 23716 57996
rect 2136 57876 2188 57928
rect 13820 57876 13872 57928
rect 17224 57876 17276 57928
rect 27160 57876 27212 57928
rect 15292 57851 15344 57860
rect 15292 57817 15301 57851
rect 15301 57817 15335 57851
rect 15335 57817 15344 57851
rect 15292 57808 15344 57817
rect 16304 57851 16356 57860
rect 16304 57817 16313 57851
rect 16313 57817 16347 57851
rect 16347 57817 16356 57851
rect 16304 57808 16356 57817
rect 17316 57808 17368 57860
rect 17868 57808 17920 57860
rect 18236 57808 18288 57860
rect 26976 57808 27028 57860
rect 27344 57808 27396 57860
rect 1584 57783 1636 57792
rect 1584 57749 1593 57783
rect 1593 57749 1627 57783
rect 1627 57749 1636 57783
rect 1584 57740 1636 57749
rect 12992 57740 13044 57792
rect 14188 57740 14240 57792
rect 15568 57740 15620 57792
rect 16488 57783 16540 57792
rect 16488 57749 16497 57783
rect 16497 57749 16531 57783
rect 16531 57749 16540 57783
rect 16488 57740 16540 57749
rect 17592 57740 17644 57792
rect 20444 57740 20496 57792
rect 26700 57740 26752 57792
rect 27436 57740 27488 57792
rect 28356 57876 28408 57928
rect 28172 57740 28224 57792
rect 29368 58080 29420 58132
rect 29092 57876 29144 57928
rect 29368 57876 29420 57928
rect 29092 57740 29144 57792
rect 29184 57740 29236 57792
rect 30104 57740 30156 57792
rect 10880 57638 10932 57690
rect 10944 57638 10996 57690
rect 11008 57638 11060 57690
rect 11072 57638 11124 57690
rect 11136 57638 11188 57690
rect 20811 57638 20863 57690
rect 20875 57638 20927 57690
rect 20939 57638 20991 57690
rect 21003 57638 21055 57690
rect 21067 57638 21119 57690
rect 1400 57536 1452 57588
rect 15292 57536 15344 57588
rect 20536 57536 20588 57588
rect 25412 57536 25464 57588
rect 29736 57536 29788 57588
rect 14924 57511 14976 57520
rect 14924 57477 14958 57511
rect 14958 57477 14976 57511
rect 14924 57468 14976 57477
rect 20260 57468 20312 57520
rect 1860 57400 1912 57452
rect 2688 57400 2740 57452
rect 13636 57400 13688 57452
rect 14096 57400 14148 57452
rect 14188 57443 14240 57452
rect 14188 57409 14197 57443
rect 14197 57409 14231 57443
rect 14231 57409 14240 57443
rect 14188 57400 14240 57409
rect 17960 57400 18012 57452
rect 19340 57400 19392 57452
rect 19616 57443 19668 57452
rect 19616 57409 19625 57443
rect 19625 57409 19659 57443
rect 19659 57409 19668 57443
rect 19616 57400 19668 57409
rect 19800 57400 19852 57452
rect 19892 57443 19944 57452
rect 19892 57409 19901 57443
rect 19901 57409 19935 57443
rect 19935 57409 19944 57443
rect 20628 57443 20680 57452
rect 19892 57400 19944 57409
rect 20628 57409 20637 57443
rect 20637 57409 20671 57443
rect 20671 57409 20680 57443
rect 20628 57400 20680 57409
rect 13820 57264 13872 57316
rect 20812 57443 20864 57452
rect 20812 57409 20821 57443
rect 20821 57409 20855 57443
rect 20855 57409 20864 57443
rect 21088 57468 21140 57520
rect 20812 57400 20864 57409
rect 26608 57468 26660 57520
rect 23112 57400 23164 57452
rect 23940 57443 23992 57452
rect 23940 57409 23949 57443
rect 23949 57409 23983 57443
rect 23983 57409 23992 57443
rect 23940 57400 23992 57409
rect 26056 57443 26108 57452
rect 26056 57409 26065 57443
rect 26065 57409 26099 57443
rect 26099 57409 26108 57443
rect 26056 57400 26108 57409
rect 26332 57443 26384 57452
rect 26332 57409 26341 57443
rect 26341 57409 26375 57443
rect 26375 57409 26384 57443
rect 26332 57400 26384 57409
rect 1584 57239 1636 57248
rect 1584 57205 1593 57239
rect 1593 57205 1627 57239
rect 1627 57205 1636 57239
rect 1584 57196 1636 57205
rect 14188 57196 14240 57248
rect 21732 57332 21784 57384
rect 25872 57332 25924 57384
rect 20720 57264 20772 57316
rect 21272 57264 21324 57316
rect 26976 57443 27028 57452
rect 26976 57409 26985 57443
rect 26985 57409 27019 57443
rect 27019 57409 27028 57443
rect 26976 57400 27028 57409
rect 27344 57332 27396 57384
rect 29184 57332 29236 57384
rect 29736 57443 29788 57452
rect 29736 57409 29745 57443
rect 29745 57409 29779 57443
rect 29779 57409 29788 57443
rect 29736 57400 29788 57409
rect 29736 57264 29788 57316
rect 15384 57196 15436 57248
rect 15660 57196 15712 57248
rect 18328 57239 18380 57248
rect 18328 57205 18337 57239
rect 18337 57205 18371 57239
rect 18371 57205 18380 57239
rect 18328 57196 18380 57205
rect 18420 57196 18472 57248
rect 20352 57239 20404 57248
rect 20352 57205 20361 57239
rect 20361 57205 20395 57239
rect 20395 57205 20404 57239
rect 20352 57196 20404 57205
rect 21548 57196 21600 57248
rect 23020 57196 23072 57248
rect 24124 57196 24176 57248
rect 24400 57196 24452 57248
rect 28172 57196 28224 57248
rect 30656 57196 30708 57248
rect 5915 57094 5967 57146
rect 5979 57094 6031 57146
rect 6043 57094 6095 57146
rect 6107 57094 6159 57146
rect 6171 57094 6223 57146
rect 15846 57094 15898 57146
rect 15910 57094 15962 57146
rect 15974 57094 16026 57146
rect 16038 57094 16090 57146
rect 16102 57094 16154 57146
rect 25776 57094 25828 57146
rect 25840 57094 25892 57146
rect 25904 57094 25956 57146
rect 25968 57094 26020 57146
rect 26032 57094 26084 57146
rect 2136 57035 2188 57044
rect 2136 57001 2145 57035
rect 2145 57001 2179 57035
rect 2179 57001 2188 57035
rect 2136 56992 2188 57001
rect 13636 56992 13688 57044
rect 16212 57035 16264 57044
rect 16212 57001 16221 57035
rect 16221 57001 16255 57035
rect 16255 57001 16264 57035
rect 16212 56992 16264 57001
rect 17684 56992 17736 57044
rect 21088 56992 21140 57044
rect 21548 56992 21600 57044
rect 21364 56924 21416 56976
rect 22560 56924 22612 56976
rect 17224 56899 17276 56908
rect 17224 56865 17233 56899
rect 17233 56865 17267 56899
rect 17267 56865 17276 56899
rect 17224 56856 17276 56865
rect 17500 56856 17552 56908
rect 17868 56899 17920 56908
rect 17868 56865 17877 56899
rect 17877 56865 17911 56899
rect 17911 56865 17920 56899
rect 17868 56856 17920 56865
rect 1400 56831 1452 56840
rect 1400 56797 1409 56831
rect 1409 56797 1443 56831
rect 1443 56797 1452 56831
rect 1400 56788 1452 56797
rect 2596 56788 2648 56840
rect 14004 56788 14056 56840
rect 14188 56788 14240 56840
rect 17684 56788 17736 56840
rect 19248 56831 19300 56840
rect 17316 56763 17368 56772
rect 17316 56729 17325 56763
rect 17325 56729 17359 56763
rect 17359 56729 17368 56763
rect 17316 56720 17368 56729
rect 19248 56797 19257 56831
rect 19257 56797 19291 56831
rect 19291 56797 19300 56831
rect 19248 56788 19300 56797
rect 20352 56788 20404 56840
rect 21272 56788 21324 56840
rect 21548 56831 21600 56840
rect 21548 56797 21557 56831
rect 21557 56797 21591 56831
rect 21591 56797 21600 56831
rect 21548 56788 21600 56797
rect 21824 56788 21876 56840
rect 19800 56720 19852 56772
rect 20260 56720 20312 56772
rect 20444 56720 20496 56772
rect 1584 56695 1636 56704
rect 1584 56661 1593 56695
rect 1593 56661 1627 56695
rect 1627 56661 1636 56695
rect 1584 56652 1636 56661
rect 17592 56652 17644 56704
rect 20628 56695 20680 56704
rect 20628 56661 20637 56695
rect 20637 56661 20671 56695
rect 20671 56661 20680 56695
rect 20628 56652 20680 56661
rect 21824 56652 21876 56704
rect 22100 56652 22152 56704
rect 23664 56992 23716 57044
rect 23480 56924 23532 56976
rect 24492 56924 24544 56976
rect 25596 56992 25648 57044
rect 24952 56856 25004 56908
rect 25596 56856 25648 56908
rect 23020 56788 23072 56840
rect 24124 56788 24176 56840
rect 24584 56831 24636 56840
rect 24584 56797 24593 56831
rect 24593 56797 24627 56831
rect 24627 56797 24636 56831
rect 24584 56788 24636 56797
rect 25228 56788 25280 56840
rect 25964 56788 26016 56840
rect 26332 56992 26384 57044
rect 27344 56924 27396 56976
rect 26240 56788 26292 56840
rect 23388 56763 23440 56772
rect 23388 56729 23397 56763
rect 23397 56729 23431 56763
rect 23431 56729 23440 56763
rect 23388 56720 23440 56729
rect 24400 56763 24452 56772
rect 24400 56729 24409 56763
rect 24409 56729 24443 56763
rect 24443 56729 24452 56763
rect 24400 56720 24452 56729
rect 24952 56763 25004 56772
rect 24952 56729 24961 56763
rect 24961 56729 24995 56763
rect 24995 56729 25004 56763
rect 24952 56720 25004 56729
rect 22468 56652 22520 56704
rect 22744 56652 22796 56704
rect 24492 56652 24544 56704
rect 25228 56652 25280 56704
rect 25872 56652 25924 56704
rect 26056 56652 26108 56704
rect 27436 56856 27488 56908
rect 29092 56992 29144 57044
rect 27344 56831 27396 56840
rect 27344 56797 27353 56831
rect 27353 56797 27387 56831
rect 27387 56797 27396 56831
rect 27344 56788 27396 56797
rect 29092 56856 29144 56908
rect 30564 56992 30616 57044
rect 28724 56788 28776 56840
rect 29736 56831 29788 56840
rect 29736 56797 29745 56831
rect 29745 56797 29779 56831
rect 29779 56797 29788 56831
rect 29736 56788 29788 56797
rect 30012 56720 30064 56772
rect 28172 56652 28224 56704
rect 10880 56550 10932 56602
rect 10944 56550 10996 56602
rect 11008 56550 11060 56602
rect 11072 56550 11124 56602
rect 11136 56550 11188 56602
rect 20811 56550 20863 56602
rect 20875 56550 20927 56602
rect 20939 56550 20991 56602
rect 21003 56550 21055 56602
rect 21067 56550 21119 56602
rect 1860 56448 1912 56500
rect 15384 56491 15436 56500
rect 15384 56457 15393 56491
rect 15393 56457 15427 56491
rect 15427 56457 15436 56491
rect 15384 56448 15436 56457
rect 22468 56448 22520 56500
rect 23020 56448 23072 56500
rect 23572 56448 23624 56500
rect 24400 56491 24452 56500
rect 24400 56457 24409 56491
rect 24409 56457 24443 56491
rect 24443 56457 24452 56491
rect 24400 56448 24452 56457
rect 16488 56380 16540 56432
rect 18420 56380 18472 56432
rect 2136 56312 2188 56364
rect 2320 56355 2372 56364
rect 2320 56321 2329 56355
rect 2329 56321 2363 56355
rect 2363 56321 2372 56355
rect 2320 56312 2372 56321
rect 14740 56312 14792 56364
rect 15568 56312 15620 56364
rect 17592 56312 17644 56364
rect 19064 56312 19116 56364
rect 22744 56380 22796 56432
rect 24216 56380 24268 56432
rect 25044 56448 25096 56500
rect 25412 56448 25464 56500
rect 25688 56448 25740 56500
rect 25872 56448 25924 56500
rect 22100 56355 22152 56364
rect 22100 56321 22134 56355
rect 22134 56321 22152 56355
rect 22100 56312 22152 56321
rect 23296 56312 23348 56364
rect 24124 56312 24176 56364
rect 24400 56312 24452 56364
rect 25964 56355 26016 56364
rect 25964 56321 25973 56355
rect 25973 56321 26007 56355
rect 26007 56321 26016 56355
rect 25964 56312 26016 56321
rect 14464 56287 14516 56296
rect 14464 56253 14473 56287
rect 14473 56253 14507 56287
rect 14507 56253 14516 56287
rect 14464 56244 14516 56253
rect 26240 56355 26292 56364
rect 26240 56321 26249 56355
rect 26249 56321 26283 56355
rect 26283 56321 26292 56355
rect 26240 56312 26292 56321
rect 28724 56355 28776 56364
rect 14004 56219 14056 56228
rect 14004 56185 14013 56219
rect 14013 56185 14047 56219
rect 14047 56185 14056 56219
rect 14004 56176 14056 56185
rect 1584 56151 1636 56160
rect 1584 56117 1593 56151
rect 1593 56117 1627 56151
rect 1627 56117 1636 56151
rect 1584 56108 1636 56117
rect 14096 56108 14148 56160
rect 18052 56108 18104 56160
rect 19340 56108 19392 56160
rect 20168 56151 20220 56160
rect 20168 56117 20177 56151
rect 20177 56117 20211 56151
rect 20211 56117 20220 56151
rect 20168 56108 20220 56117
rect 21548 56108 21600 56160
rect 27160 56244 27212 56296
rect 28724 56321 28733 56355
rect 28733 56321 28767 56355
rect 28767 56321 28776 56355
rect 28724 56312 28776 56321
rect 29184 56448 29236 56500
rect 29736 56448 29788 56500
rect 29920 56448 29972 56500
rect 29092 56380 29144 56432
rect 30012 56312 30064 56364
rect 29092 56244 29144 56296
rect 24124 56219 24176 56228
rect 24124 56185 24133 56219
rect 24133 56185 24167 56219
rect 24167 56185 24176 56219
rect 24124 56176 24176 56185
rect 27344 56176 27396 56228
rect 30748 56176 30800 56228
rect 31576 56176 31628 56228
rect 24216 56108 24268 56160
rect 26608 56108 26660 56160
rect 5915 56006 5967 56058
rect 5979 56006 6031 56058
rect 6043 56006 6095 56058
rect 6107 56006 6159 56058
rect 6171 56006 6223 56058
rect 15846 56006 15898 56058
rect 15910 56006 15962 56058
rect 15974 56006 16026 56058
rect 16038 56006 16090 56058
rect 16102 56006 16154 56058
rect 25776 56006 25828 56058
rect 25840 56006 25892 56058
rect 25904 56006 25956 56058
rect 25968 56006 26020 56058
rect 26032 56006 26084 56058
rect 1400 55904 1452 55956
rect 2688 55904 2740 55956
rect 15384 55904 15436 55956
rect 21180 55904 21232 55956
rect 21272 55904 21324 55956
rect 24400 55947 24452 55956
rect 2320 55836 2372 55888
rect 15200 55836 15252 55888
rect 16304 55836 16356 55888
rect 21824 55836 21876 55888
rect 16212 55811 16264 55820
rect 16212 55777 16221 55811
rect 16221 55777 16255 55811
rect 16255 55777 16264 55811
rect 16212 55768 16264 55777
rect 24400 55913 24409 55947
rect 24409 55913 24443 55947
rect 24443 55913 24452 55947
rect 24400 55904 24452 55913
rect 24492 55904 24544 55956
rect 24584 55904 24636 55956
rect 25688 55904 25740 55956
rect 30748 55904 30800 55956
rect 31392 55904 31444 55956
rect 1860 55743 1912 55752
rect 1860 55709 1869 55743
rect 1869 55709 1903 55743
rect 1903 55709 1912 55743
rect 1860 55700 1912 55709
rect 18696 55700 18748 55752
rect 24400 55768 24452 55820
rect 22468 55700 22520 55752
rect 23112 55700 23164 55752
rect 24584 55743 24636 55752
rect 24584 55709 24593 55743
rect 24593 55709 24627 55743
rect 24627 55709 24636 55743
rect 24584 55700 24636 55709
rect 16580 55632 16632 55684
rect 16948 55675 17000 55684
rect 16948 55641 16957 55675
rect 16957 55641 16991 55675
rect 16991 55641 17000 55675
rect 16948 55632 17000 55641
rect 19616 55675 19668 55684
rect 19616 55641 19625 55675
rect 19625 55641 19659 55675
rect 19659 55641 19668 55675
rect 19616 55632 19668 55641
rect 17776 55564 17828 55616
rect 18236 55607 18288 55616
rect 18236 55573 18245 55607
rect 18245 55573 18279 55607
rect 18279 55573 18288 55607
rect 18236 55564 18288 55573
rect 21916 55564 21968 55616
rect 24492 55632 24544 55684
rect 30564 55836 30616 55888
rect 31300 55836 31352 55888
rect 25964 55768 26016 55820
rect 27436 55768 27488 55820
rect 28908 55768 28960 55820
rect 30656 55768 30708 55820
rect 31668 55768 31720 55820
rect 25504 55675 25556 55684
rect 25504 55641 25513 55675
rect 25513 55641 25547 55675
rect 25547 55641 25556 55675
rect 25504 55632 25556 55641
rect 25688 55675 25740 55684
rect 25688 55641 25697 55675
rect 25697 55641 25731 55675
rect 25731 55641 25740 55675
rect 25688 55632 25740 55641
rect 22560 55564 22612 55616
rect 22744 55564 22796 55616
rect 24216 55564 24268 55616
rect 25044 55564 25096 55616
rect 25320 55564 25372 55616
rect 28448 55743 28500 55752
rect 28448 55709 28457 55743
rect 28457 55709 28491 55743
rect 28491 55709 28500 55743
rect 28448 55700 28500 55709
rect 25964 55632 26016 55684
rect 27160 55632 27212 55684
rect 29736 55675 29788 55684
rect 29736 55641 29745 55675
rect 29745 55641 29779 55675
rect 29779 55641 29788 55675
rect 29736 55632 29788 55641
rect 30932 55632 30984 55684
rect 31760 55632 31812 55684
rect 26516 55564 26568 55616
rect 26792 55564 26844 55616
rect 28632 55564 28684 55616
rect 29368 55564 29420 55616
rect 10880 55462 10932 55514
rect 10944 55462 10996 55514
rect 11008 55462 11060 55514
rect 11072 55462 11124 55514
rect 11136 55462 11188 55514
rect 20811 55462 20863 55514
rect 20875 55462 20927 55514
rect 20939 55462 20991 55514
rect 21003 55462 21055 55514
rect 21067 55462 21119 55514
rect 2136 55403 2188 55412
rect 2136 55369 2145 55403
rect 2145 55369 2179 55403
rect 2179 55369 2188 55403
rect 2136 55360 2188 55369
rect 16580 55360 16632 55412
rect 17316 55403 17368 55412
rect 17316 55369 17325 55403
rect 17325 55369 17359 55403
rect 17359 55369 17368 55403
rect 17316 55360 17368 55369
rect 17960 55360 18012 55412
rect 18880 55360 18932 55412
rect 16212 55292 16264 55344
rect 1400 55267 1452 55276
rect 1400 55233 1409 55267
rect 1409 55233 1443 55267
rect 1443 55233 1452 55267
rect 1400 55224 1452 55233
rect 4804 55224 4856 55276
rect 18328 55292 18380 55344
rect 17224 55267 17276 55276
rect 17224 55233 17233 55267
rect 17233 55233 17267 55267
rect 17267 55233 17276 55267
rect 17224 55224 17276 55233
rect 17684 55224 17736 55276
rect 19800 55267 19852 55276
rect 19800 55233 19809 55267
rect 19809 55233 19843 55267
rect 19843 55233 19852 55267
rect 19800 55224 19852 55233
rect 20720 55360 20772 55412
rect 23112 55360 23164 55412
rect 23664 55360 23716 55412
rect 24952 55360 25004 55412
rect 25780 55403 25832 55412
rect 25780 55369 25789 55403
rect 25789 55369 25823 55403
rect 25823 55369 25832 55403
rect 25780 55360 25832 55369
rect 27528 55360 27580 55412
rect 19708 55156 19760 55208
rect 21272 55224 21324 55276
rect 23296 55224 23348 55276
rect 25412 55292 25464 55344
rect 25872 55335 25924 55344
rect 25872 55301 25881 55335
rect 25881 55301 25915 55335
rect 25915 55301 25924 55335
rect 25872 55292 25924 55301
rect 26424 55292 26476 55344
rect 24584 55224 24636 55276
rect 29184 55360 29236 55412
rect 30288 55360 30340 55412
rect 28448 55292 28500 55344
rect 20260 55156 20312 55208
rect 20628 55156 20680 55208
rect 23204 55156 23256 55208
rect 24492 55199 24544 55208
rect 1584 55131 1636 55140
rect 1584 55097 1593 55131
rect 1593 55097 1627 55131
rect 1627 55097 1636 55131
rect 1584 55088 1636 55097
rect 23664 55088 23716 55140
rect 14648 55020 14700 55072
rect 18788 55020 18840 55072
rect 19800 55020 19852 55072
rect 23204 55063 23256 55072
rect 23204 55029 23213 55063
rect 23213 55029 23247 55063
rect 23247 55029 23256 55063
rect 23204 55020 23256 55029
rect 23572 55020 23624 55072
rect 24492 55165 24501 55199
rect 24501 55165 24535 55199
rect 24535 55165 24544 55199
rect 24492 55156 24544 55165
rect 24216 55088 24268 55140
rect 25044 55156 25096 55208
rect 25320 55156 25372 55208
rect 25228 55088 25280 55140
rect 25320 55020 25372 55072
rect 27344 55088 27396 55140
rect 26240 55020 26292 55072
rect 28632 55224 28684 55276
rect 28172 55088 28224 55140
rect 28632 55020 28684 55072
rect 28816 55224 28868 55276
rect 30932 55292 30984 55344
rect 30012 55224 30064 55276
rect 31668 55156 31720 55208
rect 30840 55088 30892 55140
rect 30012 55020 30064 55072
rect 5915 54918 5967 54970
rect 5979 54918 6031 54970
rect 6043 54918 6095 54970
rect 6107 54918 6159 54970
rect 6171 54918 6223 54970
rect 15846 54918 15898 54970
rect 15910 54918 15962 54970
rect 15974 54918 16026 54970
rect 16038 54918 16090 54970
rect 16102 54918 16154 54970
rect 25776 54918 25828 54970
rect 25840 54918 25892 54970
rect 25904 54918 25956 54970
rect 25968 54918 26020 54970
rect 26032 54918 26084 54970
rect 15476 54816 15528 54868
rect 13360 54748 13412 54800
rect 21824 54816 21876 54868
rect 23664 54816 23716 54868
rect 24584 54816 24636 54868
rect 26148 54816 26200 54868
rect 26976 54816 27028 54868
rect 28632 54816 28684 54868
rect 30380 54816 30432 54868
rect 31208 54816 31260 54868
rect 17408 54748 17460 54800
rect 22652 54748 22704 54800
rect 26056 54748 26108 54800
rect 27436 54748 27488 54800
rect 2136 54612 2188 54664
rect 2596 54544 2648 54596
rect 20444 54680 20496 54732
rect 23664 54680 23716 54732
rect 24032 54680 24084 54732
rect 26976 54680 27028 54732
rect 30932 54680 30984 54732
rect 16304 54655 16356 54664
rect 16304 54621 16313 54655
rect 16313 54621 16347 54655
rect 16347 54621 16356 54655
rect 16304 54612 16356 54621
rect 17040 54544 17092 54596
rect 22100 54587 22152 54596
rect 22100 54553 22109 54587
rect 22109 54553 22143 54587
rect 22143 54553 22152 54587
rect 26240 54612 26292 54664
rect 29736 54655 29788 54664
rect 22100 54544 22152 54553
rect 27344 54544 27396 54596
rect 27620 54544 27672 54596
rect 28632 54587 28684 54596
rect 28632 54553 28641 54587
rect 28641 54553 28675 54587
rect 28675 54553 28684 54587
rect 28632 54544 28684 54553
rect 29736 54621 29745 54655
rect 29745 54621 29779 54655
rect 29779 54621 29788 54655
rect 29736 54612 29788 54621
rect 30380 54612 30432 54664
rect 31300 54612 31352 54664
rect 30288 54544 30340 54596
rect 1584 54519 1636 54528
rect 1584 54485 1593 54519
rect 1593 54485 1627 54519
rect 1627 54485 1636 54519
rect 1584 54476 1636 54485
rect 16672 54476 16724 54528
rect 22284 54476 22336 54528
rect 23388 54519 23440 54528
rect 23388 54485 23397 54519
rect 23397 54485 23431 54519
rect 23431 54485 23440 54519
rect 23388 54476 23440 54485
rect 24216 54476 24268 54528
rect 26148 54476 26200 54528
rect 28172 54476 28224 54528
rect 31300 54476 31352 54528
rect 10880 54374 10932 54426
rect 10944 54374 10996 54426
rect 11008 54374 11060 54426
rect 11072 54374 11124 54426
rect 11136 54374 11188 54426
rect 20811 54374 20863 54426
rect 20875 54374 20927 54426
rect 20939 54374 20991 54426
rect 21003 54374 21055 54426
rect 21067 54374 21119 54426
rect 1400 54272 1452 54324
rect 17408 54272 17460 54324
rect 19892 54272 19944 54324
rect 25320 54272 25372 54324
rect 27344 54272 27396 54324
rect 16856 54204 16908 54256
rect 19340 54204 19392 54256
rect 1400 54179 1452 54188
rect 1400 54145 1409 54179
rect 1409 54145 1443 54179
rect 1443 54145 1452 54179
rect 1400 54136 1452 54145
rect 7564 54136 7616 54188
rect 16672 54179 16724 54188
rect 16672 54145 16681 54179
rect 16681 54145 16715 54179
rect 16715 54145 16724 54179
rect 16672 54136 16724 54145
rect 19800 54136 19852 54188
rect 22836 54204 22888 54256
rect 29368 54272 29420 54324
rect 29460 54272 29512 54324
rect 23296 54179 23348 54188
rect 23296 54145 23305 54179
rect 23305 54145 23339 54179
rect 23339 54145 23348 54179
rect 23296 54136 23348 54145
rect 25228 54179 25280 54188
rect 25228 54145 25237 54179
rect 25237 54145 25271 54179
rect 25271 54145 25280 54179
rect 25228 54136 25280 54145
rect 27436 54136 27488 54188
rect 19708 54111 19760 54120
rect 19708 54077 19717 54111
rect 19717 54077 19751 54111
rect 19751 54077 19760 54111
rect 19708 54068 19760 54077
rect 25044 54068 25096 54120
rect 27620 54068 27672 54120
rect 29368 54179 29420 54188
rect 29368 54145 29377 54179
rect 29377 54145 29411 54179
rect 29411 54145 29420 54179
rect 29368 54136 29420 54145
rect 30196 54272 30248 54324
rect 30012 54136 30064 54188
rect 31392 54068 31444 54120
rect 29092 54000 29144 54052
rect 30288 54000 30340 54052
rect 1584 53975 1636 53984
rect 1584 53941 1593 53975
rect 1593 53941 1627 53975
rect 1627 53941 1636 53975
rect 1584 53932 1636 53941
rect 24032 53932 24084 53984
rect 24492 53932 24544 53984
rect 27160 53932 27212 53984
rect 29644 53932 29696 53984
rect 30196 53932 30248 53984
rect 5915 53830 5967 53882
rect 5979 53830 6031 53882
rect 6043 53830 6095 53882
rect 6107 53830 6159 53882
rect 6171 53830 6223 53882
rect 15846 53830 15898 53882
rect 15910 53830 15962 53882
rect 15974 53830 16026 53882
rect 16038 53830 16090 53882
rect 16102 53830 16154 53882
rect 25776 53830 25828 53882
rect 25840 53830 25892 53882
rect 25904 53830 25956 53882
rect 25968 53830 26020 53882
rect 26032 53830 26084 53882
rect 2136 53771 2188 53780
rect 2136 53737 2145 53771
rect 2145 53737 2179 53771
rect 2179 53737 2188 53771
rect 2136 53728 2188 53737
rect 18052 53771 18104 53780
rect 18052 53737 18061 53771
rect 18061 53737 18095 53771
rect 18095 53737 18104 53771
rect 18052 53728 18104 53737
rect 18696 53771 18748 53780
rect 18696 53737 18705 53771
rect 18705 53737 18739 53771
rect 18739 53737 18748 53771
rect 18696 53728 18748 53737
rect 19432 53771 19484 53780
rect 19432 53737 19441 53771
rect 19441 53737 19475 53771
rect 19475 53737 19484 53771
rect 19432 53728 19484 53737
rect 29644 53728 29696 53780
rect 31024 53728 31076 53780
rect 22192 53660 22244 53712
rect 19340 53592 19392 53644
rect 19800 53592 19852 53644
rect 23112 53592 23164 53644
rect 24400 53592 24452 53644
rect 25872 53592 25924 53644
rect 2228 53524 2280 53576
rect 6276 53524 6328 53576
rect 17868 53567 17920 53576
rect 17868 53533 17877 53567
rect 17877 53533 17911 53567
rect 17911 53533 17920 53567
rect 17868 53524 17920 53533
rect 19984 53567 20036 53576
rect 19984 53533 19993 53567
rect 19993 53533 20027 53567
rect 20027 53533 20036 53567
rect 19984 53524 20036 53533
rect 22376 53567 22428 53576
rect 22376 53533 22385 53567
rect 22385 53533 22419 53567
rect 22419 53533 22428 53567
rect 22376 53524 22428 53533
rect 21180 53456 21232 53508
rect 22560 53456 22612 53508
rect 23112 53456 23164 53508
rect 26148 53524 26200 53576
rect 26976 53567 27028 53576
rect 26976 53533 26985 53567
rect 26985 53533 27019 53567
rect 27019 53533 27028 53567
rect 27988 53567 28040 53576
rect 26976 53524 27028 53533
rect 27988 53533 27997 53567
rect 27997 53533 28031 53567
rect 28031 53533 28040 53567
rect 27988 53524 28040 53533
rect 28724 53567 28776 53576
rect 28724 53533 28733 53567
rect 28733 53533 28767 53567
rect 28767 53533 28776 53567
rect 28724 53524 28776 53533
rect 29736 53567 29788 53576
rect 29736 53533 29745 53567
rect 29745 53533 29779 53567
rect 29779 53533 29788 53567
rect 29736 53524 29788 53533
rect 1584 53431 1636 53440
rect 1584 53397 1593 53431
rect 1593 53397 1627 53431
rect 1627 53397 1636 53431
rect 1584 53388 1636 53397
rect 21272 53431 21324 53440
rect 21272 53397 21281 53431
rect 21281 53397 21315 53431
rect 21315 53397 21324 53431
rect 21272 53388 21324 53397
rect 22468 53431 22520 53440
rect 22468 53397 22477 53431
rect 22477 53397 22511 53431
rect 22511 53397 22520 53431
rect 22468 53388 22520 53397
rect 25964 53431 26016 53440
rect 25964 53397 25973 53431
rect 25973 53397 26007 53431
rect 26007 53397 26016 53431
rect 25964 53388 26016 53397
rect 26516 53431 26568 53440
rect 26516 53397 26525 53431
rect 26525 53397 26559 53431
rect 26559 53397 26568 53431
rect 26516 53388 26568 53397
rect 27712 53388 27764 53440
rect 28172 53431 28224 53440
rect 28172 53397 28181 53431
rect 28181 53397 28215 53431
rect 28215 53397 28224 53431
rect 28172 53388 28224 53397
rect 29092 53388 29144 53440
rect 29736 53388 29788 53440
rect 10880 53286 10932 53338
rect 10944 53286 10996 53338
rect 11008 53286 11060 53338
rect 11072 53286 11124 53338
rect 11136 53286 11188 53338
rect 20811 53286 20863 53338
rect 20875 53286 20927 53338
rect 20939 53286 20991 53338
rect 21003 53286 21055 53338
rect 21067 53286 21119 53338
rect 1400 53184 1452 53236
rect 2228 53184 2280 53236
rect 17776 53227 17828 53236
rect 1952 53048 2004 53100
rect 14188 53091 14240 53100
rect 14188 53057 14222 53091
rect 14222 53057 14240 53091
rect 14188 53048 14240 53057
rect 13912 53023 13964 53032
rect 13912 52989 13921 53023
rect 13921 52989 13955 53023
rect 13955 52989 13964 53023
rect 13912 52980 13964 52989
rect 17776 53193 17785 53227
rect 17785 53193 17819 53227
rect 17819 53193 17828 53227
rect 17776 53184 17828 53193
rect 19248 53184 19300 53236
rect 19708 53184 19760 53236
rect 22100 53184 22152 53236
rect 27896 53184 27948 53236
rect 28172 53184 28224 53236
rect 29276 53227 29328 53236
rect 18236 53116 18288 53168
rect 20168 53116 20220 53168
rect 20720 53116 20772 53168
rect 25320 53116 25372 53168
rect 26516 53116 26568 53168
rect 18328 53091 18380 53100
rect 18328 53057 18337 53091
rect 18337 53057 18371 53091
rect 18371 53057 18380 53091
rect 18328 53048 18380 53057
rect 19156 53048 19208 53100
rect 21824 53048 21876 53100
rect 22100 53048 22152 53100
rect 22376 53048 22428 53100
rect 23664 53048 23716 53100
rect 26148 53091 26200 53100
rect 26148 53057 26157 53091
rect 26157 53057 26191 53091
rect 26191 53057 26200 53091
rect 26148 53048 26200 53057
rect 23296 52980 23348 53032
rect 27344 53048 27396 53100
rect 27620 53048 27672 53100
rect 19248 52955 19300 52964
rect 19248 52921 19257 52955
rect 19257 52921 19291 52955
rect 19291 52921 19300 52955
rect 19248 52912 19300 52921
rect 21916 52912 21968 52964
rect 26976 52980 27028 53032
rect 25872 52912 25924 52964
rect 27712 52912 27764 52964
rect 27896 53091 27948 53100
rect 27896 53057 27905 53091
rect 27905 53057 27939 53091
rect 27939 53057 27948 53091
rect 28448 53116 28500 53168
rect 27896 53048 27948 53057
rect 28632 53048 28684 53100
rect 29276 53193 29285 53227
rect 29285 53193 29319 53227
rect 29319 53193 29328 53227
rect 29276 53184 29328 53193
rect 29644 53048 29696 53100
rect 30012 53048 30064 53100
rect 29736 52980 29788 53032
rect 30932 52980 30984 53032
rect 29276 52912 29328 52964
rect 14280 52844 14332 52896
rect 19800 52844 19852 52896
rect 20628 52844 20680 52896
rect 23664 52887 23716 52896
rect 23664 52853 23673 52887
rect 23673 52853 23707 52887
rect 23707 52853 23716 52887
rect 23664 52844 23716 52853
rect 26332 52844 26384 52896
rect 28632 52844 28684 52896
rect 29828 52844 29880 52896
rect 31668 52844 31720 52896
rect 5915 52742 5967 52794
rect 5979 52742 6031 52794
rect 6043 52742 6095 52794
rect 6107 52742 6159 52794
rect 6171 52742 6223 52794
rect 15846 52742 15898 52794
rect 15910 52742 15962 52794
rect 15974 52742 16026 52794
rect 16038 52742 16090 52794
rect 16102 52742 16154 52794
rect 25776 52742 25828 52794
rect 25840 52742 25892 52794
rect 25904 52742 25956 52794
rect 25968 52742 26020 52794
rect 26032 52742 26084 52794
rect 13360 52683 13412 52692
rect 13360 52649 13369 52683
rect 13369 52649 13403 52683
rect 13403 52649 13412 52683
rect 13360 52640 13412 52649
rect 13544 52640 13596 52692
rect 13912 52640 13964 52692
rect 17868 52640 17920 52692
rect 18328 52640 18380 52692
rect 20536 52640 20588 52692
rect 23296 52683 23348 52692
rect 23296 52649 23305 52683
rect 23305 52649 23339 52683
rect 23339 52649 23348 52683
rect 23296 52640 23348 52649
rect 26608 52640 26660 52692
rect 1492 52572 1544 52624
rect 2044 52615 2096 52624
rect 2044 52581 2053 52615
rect 2053 52581 2087 52615
rect 2087 52581 2096 52615
rect 2044 52572 2096 52581
rect 14188 52572 14240 52624
rect 18512 52572 18564 52624
rect 21732 52572 21784 52624
rect 2872 52504 2924 52556
rect 1584 52479 1636 52488
rect 1584 52445 1593 52479
rect 1593 52445 1627 52479
rect 1627 52445 1636 52479
rect 1584 52436 1636 52445
rect 2228 52479 2280 52488
rect 2228 52445 2237 52479
rect 2237 52445 2271 52479
rect 2271 52445 2280 52479
rect 2228 52436 2280 52445
rect 11796 52479 11848 52488
rect 11796 52445 11805 52479
rect 11805 52445 11839 52479
rect 11839 52445 11848 52479
rect 11796 52436 11848 52445
rect 11888 52436 11940 52488
rect 14280 52436 14332 52488
rect 20628 52504 20680 52556
rect 21916 52547 21968 52556
rect 21916 52513 21925 52547
rect 21925 52513 21959 52547
rect 21959 52513 21968 52547
rect 21916 52504 21968 52513
rect 23756 52504 23808 52556
rect 24308 52504 24360 52556
rect 27528 52572 27580 52624
rect 14832 52436 14884 52488
rect 18052 52436 18104 52488
rect 18328 52436 18380 52488
rect 14924 52368 14976 52420
rect 14372 52300 14424 52352
rect 17776 52368 17828 52420
rect 19892 52411 19944 52420
rect 19892 52377 19901 52411
rect 19901 52377 19935 52411
rect 19935 52377 19944 52411
rect 19892 52368 19944 52377
rect 20720 52436 20772 52488
rect 26148 52436 26200 52488
rect 26976 52436 27028 52488
rect 27344 52436 27396 52488
rect 29184 52640 29236 52692
rect 29460 52640 29512 52692
rect 30012 52640 30064 52692
rect 27988 52504 28040 52556
rect 28632 52572 28684 52624
rect 30840 52572 30892 52624
rect 22192 52411 22244 52420
rect 22192 52377 22226 52411
rect 22226 52377 22244 52411
rect 19800 52343 19852 52352
rect 19800 52309 19809 52343
rect 19809 52309 19843 52343
rect 19843 52309 19852 52343
rect 19800 52300 19852 52309
rect 20444 52300 20496 52352
rect 22192 52368 22244 52377
rect 23940 52368 23992 52420
rect 24308 52368 24360 52420
rect 27988 52368 28040 52420
rect 23020 52300 23072 52352
rect 25964 52300 26016 52352
rect 26700 52300 26752 52352
rect 26884 52300 26936 52352
rect 27436 52300 27488 52352
rect 28448 52479 28500 52488
rect 28448 52445 28457 52479
rect 28457 52445 28491 52479
rect 28491 52445 28500 52479
rect 28448 52436 28500 52445
rect 28632 52479 28684 52488
rect 28632 52445 28641 52479
rect 28641 52445 28675 52479
rect 28675 52445 28684 52479
rect 28632 52436 28684 52445
rect 28908 52504 28960 52556
rect 29000 52504 29052 52556
rect 29276 52504 29328 52556
rect 29736 52411 29788 52420
rect 29736 52377 29745 52411
rect 29745 52377 29779 52411
rect 29779 52377 29788 52411
rect 29736 52368 29788 52377
rect 29000 52343 29052 52352
rect 29000 52309 29009 52343
rect 29009 52309 29043 52343
rect 29043 52309 29052 52343
rect 29000 52300 29052 52309
rect 29552 52300 29604 52352
rect 10880 52198 10932 52250
rect 10944 52198 10996 52250
rect 11008 52198 11060 52250
rect 11072 52198 11124 52250
rect 11136 52198 11188 52250
rect 20811 52198 20863 52250
rect 20875 52198 20927 52250
rect 20939 52198 20991 52250
rect 21003 52198 21055 52250
rect 21067 52198 21119 52250
rect 2228 52096 2280 52148
rect 11796 52096 11848 52148
rect 14004 52028 14056 52080
rect 14648 52028 14700 52080
rect 16948 52096 17000 52148
rect 18052 52071 18104 52080
rect 18052 52037 18061 52071
rect 18061 52037 18095 52071
rect 18095 52037 18104 52071
rect 18052 52028 18104 52037
rect 19800 52096 19852 52148
rect 22468 52096 22520 52148
rect 23020 52096 23072 52148
rect 23572 52096 23624 52148
rect 24400 52096 24452 52148
rect 25964 52139 26016 52148
rect 25964 52105 25973 52139
rect 25973 52105 26007 52139
rect 26007 52105 26016 52139
rect 25964 52096 26016 52105
rect 27436 52096 27488 52148
rect 28724 52096 28776 52148
rect 29368 52096 29420 52148
rect 25688 52028 25740 52080
rect 26608 52028 26660 52080
rect 11612 51960 11664 52012
rect 14464 51960 14516 52012
rect 17040 52003 17092 52012
rect 17040 51969 17049 52003
rect 17049 51969 17083 52003
rect 17083 51969 17092 52003
rect 17040 51960 17092 51969
rect 17960 51960 18012 52012
rect 20720 51960 20772 52012
rect 22928 51960 22980 52012
rect 25596 51960 25648 52012
rect 27344 52003 27396 52012
rect 27344 51969 27353 52003
rect 27353 51969 27387 52003
rect 27387 51969 27396 52003
rect 27344 51960 27396 51969
rect 28448 52028 28500 52080
rect 27712 52003 27764 52012
rect 12624 51935 12676 51944
rect 12624 51901 12633 51935
rect 12633 51901 12667 51935
rect 12667 51901 12676 51935
rect 12624 51892 12676 51901
rect 12900 51935 12952 51944
rect 12900 51901 12909 51935
rect 12909 51901 12943 51935
rect 12943 51901 12952 51935
rect 12900 51892 12952 51901
rect 14740 51935 14792 51944
rect 14740 51901 14749 51935
rect 14749 51901 14783 51935
rect 14783 51901 14792 51935
rect 14740 51892 14792 51901
rect 18328 51935 18380 51944
rect 18328 51901 18337 51935
rect 18337 51901 18371 51935
rect 18371 51901 18380 51935
rect 18328 51892 18380 51901
rect 21732 51892 21784 51944
rect 22560 51892 22612 51944
rect 24400 51892 24452 51944
rect 26608 51892 26660 51944
rect 27712 51969 27721 52003
rect 27721 51969 27755 52003
rect 27755 51969 27764 52003
rect 27712 51960 27764 51969
rect 19156 51824 19208 51876
rect 15752 51756 15804 51808
rect 24216 51824 24268 51876
rect 25412 51824 25464 51876
rect 26976 51824 27028 51876
rect 29184 51960 29236 52012
rect 29644 52028 29696 52080
rect 30012 52028 30064 52080
rect 30472 52028 30524 52080
rect 23848 51756 23900 51808
rect 28908 51892 28960 51944
rect 29276 51892 29328 51944
rect 29644 51935 29696 51944
rect 29644 51901 29653 51935
rect 29653 51901 29687 51935
rect 29687 51901 29696 51935
rect 29644 51892 29696 51901
rect 29092 51756 29144 51808
rect 29460 51756 29512 51808
rect 5915 51654 5967 51706
rect 5979 51654 6031 51706
rect 6043 51654 6095 51706
rect 6107 51654 6159 51706
rect 6171 51654 6223 51706
rect 15846 51654 15898 51706
rect 15910 51654 15962 51706
rect 15974 51654 16026 51706
rect 16038 51654 16090 51706
rect 16102 51654 16154 51706
rect 25776 51654 25828 51706
rect 25840 51654 25892 51706
rect 25904 51654 25956 51706
rect 25968 51654 26020 51706
rect 26032 51654 26084 51706
rect 12624 51552 12676 51604
rect 14464 51595 14516 51604
rect 14464 51561 14473 51595
rect 14473 51561 14507 51595
rect 14507 51561 14516 51595
rect 14464 51552 14516 51561
rect 14740 51552 14792 51604
rect 17960 51595 18012 51604
rect 17960 51561 17969 51595
rect 17969 51561 18003 51595
rect 18003 51561 18012 51595
rect 17960 51552 18012 51561
rect 19340 51595 19392 51604
rect 19340 51561 19349 51595
rect 19349 51561 19383 51595
rect 19383 51561 19392 51595
rect 19340 51552 19392 51561
rect 19524 51552 19576 51604
rect 22192 51552 22244 51604
rect 27620 51552 27672 51604
rect 29644 51552 29696 51604
rect 25320 51484 25372 51536
rect 25964 51484 26016 51536
rect 29460 51484 29512 51536
rect 30472 51484 30524 51536
rect 1400 51348 1452 51400
rect 2228 51391 2280 51400
rect 2228 51357 2237 51391
rect 2237 51357 2271 51391
rect 2271 51357 2280 51391
rect 2228 51348 2280 51357
rect 14648 51348 14700 51400
rect 15752 51416 15804 51468
rect 18328 51416 18380 51468
rect 19892 51459 19944 51468
rect 19892 51425 19901 51459
rect 19901 51425 19935 51459
rect 19935 51425 19944 51459
rect 19892 51416 19944 51425
rect 14372 51280 14424 51332
rect 14924 51391 14976 51400
rect 14924 51357 14933 51391
rect 14933 51357 14967 51391
rect 14967 51357 14976 51391
rect 14924 51348 14976 51357
rect 1768 51212 1820 51264
rect 2044 51255 2096 51264
rect 2044 51221 2053 51255
rect 2053 51221 2087 51255
rect 2087 51221 2096 51255
rect 2044 51212 2096 51221
rect 12624 51212 12676 51264
rect 15384 51348 15436 51400
rect 17684 51348 17736 51400
rect 20628 51348 20680 51400
rect 22468 51391 22520 51400
rect 22468 51357 22477 51391
rect 22477 51357 22511 51391
rect 22511 51357 22520 51391
rect 22468 51348 22520 51357
rect 23296 51416 23348 51468
rect 24032 51416 24084 51468
rect 24400 51416 24452 51468
rect 22652 51348 22704 51400
rect 22836 51391 22888 51400
rect 22836 51357 22845 51391
rect 22845 51357 22879 51391
rect 22879 51357 22888 51391
rect 24584 51391 24636 51400
rect 22836 51348 22888 51357
rect 24584 51357 24593 51391
rect 24593 51357 24627 51391
rect 24627 51357 24636 51391
rect 24584 51348 24636 51357
rect 26148 51416 26200 51468
rect 29368 51416 29420 51468
rect 17224 51280 17276 51332
rect 19800 51323 19852 51332
rect 19800 51289 19809 51323
rect 19809 51289 19843 51323
rect 19843 51289 19852 51323
rect 19800 51280 19852 51289
rect 24400 51323 24452 51332
rect 24400 51289 24409 51323
rect 24409 51289 24443 51323
rect 24443 51289 24452 51323
rect 24400 51280 24452 51289
rect 20628 51212 20680 51264
rect 21364 51212 21416 51264
rect 23388 51212 23440 51264
rect 24492 51212 24544 51264
rect 24952 51323 25004 51332
rect 24952 51289 24961 51323
rect 24961 51289 24995 51323
rect 24995 51289 25004 51323
rect 24952 51280 25004 51289
rect 24768 51255 24820 51264
rect 24768 51221 24777 51255
rect 24777 51221 24811 51255
rect 24811 51221 24820 51255
rect 25320 51348 25372 51400
rect 28724 51391 28776 51400
rect 25596 51280 25648 51332
rect 26056 51280 26108 51332
rect 28724 51357 28733 51391
rect 28733 51357 28767 51391
rect 28767 51357 28776 51391
rect 28724 51348 28776 51357
rect 27620 51280 27672 51332
rect 27804 51280 27856 51332
rect 24768 51212 24820 51221
rect 26332 51212 26384 51264
rect 28908 51255 28960 51264
rect 28908 51221 28917 51255
rect 28917 51221 28951 51255
rect 28951 51221 28960 51255
rect 28908 51212 28960 51221
rect 29092 51212 29144 51264
rect 29920 51280 29972 51332
rect 30288 51212 30340 51264
rect 30472 51212 30524 51264
rect 10880 51110 10932 51162
rect 10944 51110 10996 51162
rect 11008 51110 11060 51162
rect 11072 51110 11124 51162
rect 11136 51110 11188 51162
rect 20811 51110 20863 51162
rect 20875 51110 20927 51162
rect 20939 51110 20991 51162
rect 21003 51110 21055 51162
rect 21067 51110 21119 51162
rect 14924 51008 14976 51060
rect 14372 50940 14424 50992
rect 1584 50915 1636 50924
rect 1584 50881 1593 50915
rect 1593 50881 1627 50915
rect 1627 50881 1636 50915
rect 1584 50872 1636 50881
rect 14924 50915 14976 50924
rect 14924 50881 14933 50915
rect 14933 50881 14967 50915
rect 14967 50881 14976 50915
rect 14924 50872 14976 50881
rect 19708 51008 19760 51060
rect 20352 51008 20404 51060
rect 15108 50915 15160 50924
rect 15108 50881 15117 50915
rect 15117 50881 15151 50915
rect 15151 50881 15160 50915
rect 15108 50872 15160 50881
rect 13728 50804 13780 50856
rect 1860 50736 1912 50788
rect 19432 50940 19484 50992
rect 21272 50940 21324 50992
rect 17316 50915 17368 50924
rect 17316 50881 17325 50915
rect 17325 50881 17359 50915
rect 17359 50881 17368 50915
rect 17316 50872 17368 50881
rect 15476 50804 15528 50856
rect 22376 51008 22428 51060
rect 22468 51008 22520 51060
rect 23940 51008 23992 51060
rect 24216 51008 24268 51060
rect 22100 50983 22152 50992
rect 22100 50949 22109 50983
rect 22109 50949 22143 50983
rect 22143 50949 22152 50983
rect 22100 50940 22152 50949
rect 23296 50940 23348 50992
rect 22284 50872 22336 50924
rect 22192 50804 22244 50856
rect 15568 50736 15620 50788
rect 21916 50736 21968 50788
rect 22008 50736 22060 50788
rect 23480 50872 23532 50924
rect 24492 50872 24544 50924
rect 25780 51008 25832 51060
rect 25964 51008 26016 51060
rect 26424 51008 26476 51060
rect 26056 50940 26108 50992
rect 23388 50804 23440 50856
rect 23756 50736 23808 50788
rect 25504 50872 25556 50924
rect 28816 50872 28868 50924
rect 29552 51008 29604 51060
rect 30840 51008 30892 51060
rect 29644 50940 29696 50992
rect 29828 50940 29880 50992
rect 24860 50804 24912 50856
rect 29000 50804 29052 50856
rect 30932 50804 30984 50856
rect 31852 50804 31904 50856
rect 24952 50736 25004 50788
rect 25780 50736 25832 50788
rect 30104 50736 30156 50788
rect 1676 50668 1728 50720
rect 15752 50668 15804 50720
rect 20168 50711 20220 50720
rect 20168 50677 20177 50711
rect 20177 50677 20211 50711
rect 20211 50677 20220 50711
rect 20168 50668 20220 50677
rect 22100 50668 22152 50720
rect 22744 50668 22796 50720
rect 29092 50711 29144 50720
rect 29092 50677 29101 50711
rect 29101 50677 29135 50711
rect 29135 50677 29144 50711
rect 29092 50668 29144 50677
rect 29828 50711 29880 50720
rect 29828 50677 29837 50711
rect 29837 50677 29871 50711
rect 29871 50677 29880 50711
rect 29828 50668 29880 50677
rect 29920 50668 29972 50720
rect 5915 50566 5967 50618
rect 5979 50566 6031 50618
rect 6043 50566 6095 50618
rect 6107 50566 6159 50618
rect 6171 50566 6223 50618
rect 15846 50566 15898 50618
rect 15910 50566 15962 50618
rect 15974 50566 16026 50618
rect 16038 50566 16090 50618
rect 16102 50566 16154 50618
rect 25776 50566 25828 50618
rect 25840 50566 25892 50618
rect 25904 50566 25956 50618
rect 25968 50566 26020 50618
rect 26032 50566 26084 50618
rect 2688 50507 2740 50516
rect 2688 50473 2697 50507
rect 2697 50473 2731 50507
rect 2731 50473 2740 50507
rect 2688 50464 2740 50473
rect 21456 50464 21508 50516
rect 21732 50507 21784 50516
rect 21732 50473 21741 50507
rect 21741 50473 21775 50507
rect 21775 50473 21784 50507
rect 21732 50464 21784 50473
rect 22376 50464 22428 50516
rect 21640 50396 21692 50448
rect 1492 50260 1544 50312
rect 2044 50260 2096 50312
rect 11888 50260 11940 50312
rect 1492 50124 1544 50176
rect 1860 50192 1912 50244
rect 10508 50192 10560 50244
rect 15476 50260 15528 50312
rect 15660 50260 15712 50312
rect 15844 50303 15896 50312
rect 15844 50269 15878 50303
rect 15878 50269 15896 50303
rect 15844 50260 15896 50269
rect 19708 50303 19760 50312
rect 19708 50269 19717 50303
rect 19717 50269 19751 50303
rect 19751 50269 19760 50303
rect 19708 50260 19760 50269
rect 19984 50260 20036 50312
rect 12256 50192 12308 50244
rect 21088 50260 21140 50312
rect 21640 50260 21692 50312
rect 22468 50303 22520 50312
rect 22468 50269 22477 50303
rect 22477 50269 22511 50303
rect 22511 50269 22520 50303
rect 22468 50260 22520 50269
rect 23020 50396 23072 50448
rect 23020 50260 23072 50312
rect 13084 50124 13136 50176
rect 23940 50396 23992 50448
rect 24768 50464 24820 50516
rect 25228 50464 25280 50516
rect 24584 50396 24636 50448
rect 24952 50396 25004 50448
rect 27896 50396 27948 50448
rect 28172 50396 28224 50448
rect 23756 50328 23808 50380
rect 23756 50236 23808 50288
rect 24032 50260 24084 50312
rect 24676 50260 24728 50312
rect 27988 50303 28040 50312
rect 27988 50269 27997 50303
rect 27997 50269 28031 50303
rect 28031 50269 28040 50303
rect 27988 50260 28040 50269
rect 14924 50124 14976 50176
rect 21548 50124 21600 50176
rect 22652 50124 22704 50176
rect 23664 50167 23716 50176
rect 23664 50133 23673 50167
rect 23673 50133 23707 50167
rect 23707 50133 23716 50167
rect 25228 50192 25280 50244
rect 27896 50192 27948 50244
rect 28540 50192 28592 50244
rect 28724 50192 28776 50244
rect 29000 50235 29052 50244
rect 29000 50201 29009 50235
rect 29009 50201 29043 50235
rect 29043 50201 29052 50235
rect 29000 50192 29052 50201
rect 29736 50235 29788 50244
rect 29736 50201 29745 50235
rect 29745 50201 29779 50235
rect 29779 50201 29788 50235
rect 29736 50192 29788 50201
rect 23664 50124 23716 50133
rect 27252 50124 27304 50176
rect 29828 50167 29880 50176
rect 29828 50133 29837 50167
rect 29837 50133 29871 50167
rect 29871 50133 29880 50167
rect 29828 50124 29880 50133
rect 10880 50022 10932 50074
rect 10944 50022 10996 50074
rect 11008 50022 11060 50074
rect 11072 50022 11124 50074
rect 11136 50022 11188 50074
rect 20811 50022 20863 50074
rect 20875 50022 20927 50074
rect 20939 50022 20991 50074
rect 21003 50022 21055 50074
rect 21067 50022 21119 50074
rect 11888 49963 11940 49972
rect 11888 49929 11897 49963
rect 11897 49929 11931 49963
rect 11931 49929 11940 49963
rect 11888 49920 11940 49929
rect 15660 49963 15712 49972
rect 15660 49929 15669 49963
rect 15669 49929 15703 49963
rect 15703 49929 15712 49963
rect 15660 49920 15712 49929
rect 19984 49963 20036 49972
rect 19984 49929 19993 49963
rect 19993 49929 20027 49963
rect 20027 49929 20036 49963
rect 19984 49920 20036 49929
rect 23020 49963 23072 49972
rect 23020 49929 23029 49963
rect 23029 49929 23063 49963
rect 23063 49929 23072 49963
rect 23020 49920 23072 49929
rect 23756 49963 23808 49972
rect 23756 49929 23765 49963
rect 23765 49929 23799 49963
rect 23799 49929 23808 49963
rect 23756 49920 23808 49929
rect 24768 49920 24820 49972
rect 1492 49852 1544 49904
rect 1768 49895 1820 49904
rect 1768 49861 1777 49895
rect 1777 49861 1811 49895
rect 1811 49861 1820 49895
rect 1768 49852 1820 49861
rect 2780 49784 2832 49836
rect 11704 49827 11756 49836
rect 11704 49793 11713 49827
rect 11713 49793 11747 49827
rect 11747 49793 11756 49827
rect 11704 49784 11756 49793
rect 14280 49784 14332 49836
rect 15476 49827 15528 49836
rect 15476 49793 15485 49827
rect 15485 49793 15519 49827
rect 15519 49793 15528 49827
rect 15476 49784 15528 49793
rect 19524 49784 19576 49836
rect 20352 49784 20404 49836
rect 22376 49827 22428 49836
rect 22376 49793 22385 49827
rect 22385 49793 22419 49827
rect 22419 49793 22428 49827
rect 22376 49784 22428 49793
rect 2504 49716 2556 49768
rect 12532 49716 12584 49768
rect 14188 49716 14240 49768
rect 14556 49716 14608 49768
rect 17132 49716 17184 49768
rect 14096 49648 14148 49700
rect 22008 49648 22060 49700
rect 2136 49580 2188 49632
rect 21548 49580 21600 49632
rect 23480 49716 23532 49768
rect 23756 49716 23808 49768
rect 24584 49784 24636 49836
rect 23296 49648 23348 49700
rect 24492 49716 24544 49768
rect 25228 49852 25280 49904
rect 24768 49784 24820 49836
rect 24768 49648 24820 49700
rect 25780 49920 25832 49972
rect 28540 49852 28592 49904
rect 29092 49852 29144 49904
rect 30932 49920 30984 49972
rect 29828 49852 29880 49904
rect 26332 49784 26384 49836
rect 27252 49784 27304 49836
rect 25228 49580 25280 49632
rect 25872 49716 25924 49768
rect 29000 49784 29052 49836
rect 27436 49648 27488 49700
rect 29736 49716 29788 49768
rect 30012 49759 30064 49768
rect 30012 49725 30021 49759
rect 30021 49725 30055 49759
rect 30055 49725 30064 49759
rect 30012 49716 30064 49725
rect 5915 49478 5967 49530
rect 5979 49478 6031 49530
rect 6043 49478 6095 49530
rect 6107 49478 6159 49530
rect 6171 49478 6223 49530
rect 15846 49478 15898 49530
rect 15910 49478 15962 49530
rect 15974 49478 16026 49530
rect 16038 49478 16090 49530
rect 16102 49478 16154 49530
rect 25776 49478 25828 49530
rect 25840 49478 25892 49530
rect 25904 49478 25956 49530
rect 25968 49478 26020 49530
rect 26032 49478 26084 49530
rect 10968 49376 11020 49428
rect 14096 49376 14148 49428
rect 14280 49419 14332 49428
rect 14280 49385 14289 49419
rect 14289 49385 14323 49419
rect 14323 49385 14332 49419
rect 14280 49376 14332 49385
rect 19708 49376 19760 49428
rect 22376 49376 22428 49428
rect 25504 49376 25556 49428
rect 26700 49419 26752 49428
rect 26700 49385 26709 49419
rect 26709 49385 26743 49419
rect 26743 49385 26752 49419
rect 26700 49376 26752 49385
rect 27620 49419 27672 49428
rect 27620 49385 27629 49419
rect 27629 49385 27663 49419
rect 27663 49385 27672 49419
rect 27620 49376 27672 49385
rect 17776 49308 17828 49360
rect 20628 49308 20680 49360
rect 23388 49308 23440 49360
rect 25228 49308 25280 49360
rect 1492 49172 1544 49224
rect 1676 49172 1728 49224
rect 9956 49215 10008 49224
rect 9956 49181 9965 49215
rect 9965 49181 9999 49215
rect 9999 49181 10008 49215
rect 9956 49172 10008 49181
rect 12072 49240 12124 49292
rect 19800 49240 19852 49292
rect 25780 49240 25832 49292
rect 27160 49308 27212 49360
rect 27436 49308 27488 49360
rect 26700 49240 26752 49292
rect 12624 49172 12676 49224
rect 14096 49215 14148 49224
rect 14096 49181 14105 49215
rect 14105 49181 14139 49215
rect 14139 49181 14148 49215
rect 14096 49172 14148 49181
rect 21732 49172 21784 49224
rect 22284 49215 22336 49224
rect 22284 49181 22293 49215
rect 22293 49181 22327 49215
rect 22327 49181 22336 49215
rect 22284 49172 22336 49181
rect 23296 49172 23348 49224
rect 25228 49172 25280 49224
rect 25872 49172 25924 49224
rect 26424 49172 26476 49224
rect 26516 49172 26568 49224
rect 27436 49172 27488 49224
rect 27896 49240 27948 49292
rect 28172 49240 28224 49292
rect 28724 49172 28776 49224
rect 2320 49104 2372 49156
rect 3240 49104 3292 49156
rect 9588 49104 9640 49156
rect 10968 49104 11020 49156
rect 12348 49104 12400 49156
rect 13176 49147 13228 49156
rect 13176 49113 13185 49147
rect 13185 49113 13219 49147
rect 13219 49113 13228 49147
rect 13176 49104 13228 49113
rect 20352 49104 20404 49156
rect 21272 49104 21324 49156
rect 22468 49104 22520 49156
rect 9864 49036 9916 49088
rect 11428 49036 11480 49088
rect 12164 49036 12216 49088
rect 20076 49079 20128 49088
rect 20076 49045 20085 49079
rect 20085 49045 20119 49079
rect 20119 49045 20128 49079
rect 20076 49036 20128 49045
rect 20720 49036 20772 49088
rect 22928 49036 22980 49088
rect 25504 49036 25556 49088
rect 28172 49104 28224 49156
rect 28356 49104 28408 49156
rect 29736 49147 29788 49156
rect 29736 49113 29745 49147
rect 29745 49113 29779 49147
rect 29779 49113 29788 49147
rect 29736 49104 29788 49113
rect 30932 49104 30984 49156
rect 26424 49036 26476 49088
rect 26976 49036 27028 49088
rect 27528 49036 27580 49088
rect 27620 49036 27672 49088
rect 10880 48934 10932 48986
rect 10944 48934 10996 48986
rect 11008 48934 11060 48986
rect 11072 48934 11124 48986
rect 11136 48934 11188 48986
rect 20811 48934 20863 48986
rect 20875 48934 20927 48986
rect 20939 48934 20991 48986
rect 21003 48934 21055 48986
rect 21067 48934 21119 48986
rect 3240 48875 3292 48884
rect 3240 48841 3249 48875
rect 3249 48841 3283 48875
rect 3283 48841 3292 48875
rect 3240 48832 3292 48841
rect 9956 48832 10008 48884
rect 1492 48764 1544 48816
rect 2136 48764 2188 48816
rect 13728 48832 13780 48884
rect 15200 48832 15252 48884
rect 11980 48764 12032 48816
rect 12164 48764 12216 48816
rect 2320 48696 2372 48748
rect 2596 48739 2648 48748
rect 2596 48705 2605 48739
rect 2605 48705 2639 48739
rect 2639 48705 2648 48739
rect 2596 48696 2648 48705
rect 3424 48739 3476 48748
rect 3424 48705 3433 48739
rect 3433 48705 3467 48739
rect 3467 48705 3476 48739
rect 3424 48696 3476 48705
rect 11428 48696 11480 48748
rect 15752 48696 15804 48748
rect 18512 48764 18564 48816
rect 19800 48807 19852 48816
rect 19800 48773 19809 48807
rect 19809 48773 19843 48807
rect 19843 48773 19852 48807
rect 19800 48764 19852 48773
rect 20168 48764 20220 48816
rect 20720 48807 20772 48816
rect 20720 48773 20729 48807
rect 20729 48773 20763 48807
rect 20763 48773 20772 48807
rect 20720 48764 20772 48773
rect 21548 48764 21600 48816
rect 22376 48764 22428 48816
rect 22928 48832 22980 48884
rect 24492 48832 24544 48884
rect 24584 48832 24636 48884
rect 25688 48875 25740 48884
rect 25688 48841 25697 48875
rect 25697 48841 25731 48875
rect 25731 48841 25740 48875
rect 25688 48832 25740 48841
rect 25872 48832 25924 48884
rect 25964 48832 26016 48884
rect 17776 48739 17828 48748
rect 12072 48671 12124 48680
rect 12072 48637 12081 48671
rect 12081 48637 12115 48671
rect 12115 48637 12124 48671
rect 12072 48628 12124 48637
rect 12164 48671 12216 48680
rect 12164 48637 12173 48671
rect 12173 48637 12207 48671
rect 12207 48637 12216 48671
rect 12164 48628 12216 48637
rect 12348 48628 12400 48680
rect 11612 48603 11664 48612
rect 11612 48569 11621 48603
rect 11621 48569 11655 48603
rect 11655 48569 11664 48603
rect 11612 48560 11664 48569
rect 14740 48603 14792 48612
rect 14740 48569 14749 48603
rect 14749 48569 14783 48603
rect 14783 48569 14792 48603
rect 14740 48560 14792 48569
rect 17776 48705 17785 48739
rect 17785 48705 17819 48739
rect 17819 48705 17828 48739
rect 17776 48696 17828 48705
rect 22100 48696 22152 48748
rect 23296 48696 23348 48748
rect 20352 48628 20404 48680
rect 17592 48560 17644 48612
rect 17776 48560 17828 48612
rect 19524 48603 19576 48612
rect 19524 48569 19533 48603
rect 19533 48569 19567 48603
rect 19567 48569 19576 48603
rect 19524 48560 19576 48569
rect 23480 48628 23532 48680
rect 1952 48535 2004 48544
rect 1952 48501 1961 48535
rect 1961 48501 1995 48535
rect 1995 48501 2004 48535
rect 1952 48492 2004 48501
rect 17408 48492 17460 48544
rect 20628 48492 20680 48544
rect 22100 48492 22152 48544
rect 22928 48560 22980 48612
rect 23020 48492 23072 48544
rect 25504 48764 25556 48816
rect 26976 48832 27028 48884
rect 28264 48832 28316 48884
rect 29000 48832 29052 48884
rect 29552 48764 29604 48816
rect 24768 48696 24820 48748
rect 25228 48696 25280 48748
rect 25780 48628 25832 48680
rect 26148 48628 26200 48680
rect 26424 48696 26476 48748
rect 26884 48696 26936 48748
rect 27160 48696 27212 48748
rect 27528 48696 27580 48748
rect 28264 48696 28316 48748
rect 29092 48696 29144 48748
rect 26700 48628 26752 48680
rect 30012 48671 30064 48680
rect 30012 48637 30021 48671
rect 30021 48637 30055 48671
rect 30055 48637 30064 48671
rect 30012 48628 30064 48637
rect 26516 48492 26568 48544
rect 26884 48492 26936 48544
rect 28264 48492 28316 48544
rect 5915 48390 5967 48442
rect 5979 48390 6031 48442
rect 6043 48390 6095 48442
rect 6107 48390 6159 48442
rect 6171 48390 6223 48442
rect 15846 48390 15898 48442
rect 15910 48390 15962 48442
rect 15974 48390 16026 48442
rect 16038 48390 16090 48442
rect 16102 48390 16154 48442
rect 25776 48390 25828 48442
rect 25840 48390 25892 48442
rect 25904 48390 25956 48442
rect 25968 48390 26020 48442
rect 26032 48390 26084 48442
rect 1492 48288 1544 48340
rect 1952 48288 2004 48340
rect 18512 48331 18564 48340
rect 2872 48220 2924 48272
rect 11704 48220 11756 48272
rect 18512 48297 18521 48331
rect 18521 48297 18555 48331
rect 18555 48297 18564 48331
rect 18512 48288 18564 48297
rect 18972 48288 19024 48340
rect 19524 48220 19576 48272
rect 2412 48084 2464 48136
rect 12072 48084 12124 48136
rect 14280 48084 14332 48136
rect 14372 48084 14424 48136
rect 19432 48152 19484 48204
rect 19800 48152 19852 48204
rect 22468 48220 22520 48272
rect 25320 48220 25372 48272
rect 26240 48288 26292 48340
rect 26424 48288 26476 48340
rect 26516 48288 26568 48340
rect 26148 48220 26200 48272
rect 2320 48059 2372 48068
rect 2320 48025 2329 48059
rect 2329 48025 2363 48059
rect 2363 48025 2372 48059
rect 2320 48016 2372 48025
rect 1768 47948 1820 48000
rect 13360 48059 13412 48068
rect 13360 48025 13369 48059
rect 13369 48025 13403 48059
rect 13403 48025 13412 48059
rect 13360 48016 13412 48025
rect 18512 48084 18564 48136
rect 19248 48127 19300 48136
rect 19248 48093 19257 48127
rect 19257 48093 19291 48127
rect 19291 48093 19300 48127
rect 19248 48084 19300 48093
rect 20352 48127 20404 48136
rect 20352 48093 20361 48127
rect 20361 48093 20395 48127
rect 20395 48093 20404 48127
rect 20352 48084 20404 48093
rect 20720 48084 20772 48136
rect 21732 48084 21784 48136
rect 15108 48016 15160 48068
rect 12164 47948 12216 48000
rect 13912 47948 13964 48000
rect 14924 47948 14976 48000
rect 16212 47991 16264 48000
rect 16212 47957 16221 47991
rect 16221 47957 16255 47991
rect 16255 47957 16264 47991
rect 16212 47948 16264 47957
rect 17408 48059 17460 48068
rect 17408 48025 17442 48059
rect 17442 48025 17460 48059
rect 17408 48016 17460 48025
rect 27896 48220 27948 48272
rect 28356 48220 28408 48272
rect 31116 48220 31168 48272
rect 25320 48084 25372 48136
rect 25688 48084 25740 48136
rect 25228 48016 25280 48068
rect 26056 48084 26108 48136
rect 26700 48084 26752 48136
rect 27528 48127 27580 48136
rect 27528 48093 27537 48127
rect 27537 48093 27571 48127
rect 27571 48093 27580 48127
rect 27528 48084 27580 48093
rect 27896 48084 27948 48136
rect 29000 48127 29052 48136
rect 29000 48093 29009 48127
rect 29009 48093 29043 48127
rect 29043 48093 29052 48127
rect 29000 48084 29052 48093
rect 31116 48084 31168 48136
rect 18420 47948 18472 48000
rect 19432 47991 19484 48000
rect 19432 47957 19441 47991
rect 19441 47957 19475 47991
rect 19475 47957 19484 47991
rect 19432 47948 19484 47957
rect 20352 47948 20404 48000
rect 20536 47948 20588 48000
rect 29000 47948 29052 48000
rect 30288 47948 30340 48000
rect 10880 47846 10932 47898
rect 10944 47846 10996 47898
rect 11008 47846 11060 47898
rect 11072 47846 11124 47898
rect 11136 47846 11188 47898
rect 20811 47846 20863 47898
rect 20875 47846 20927 47898
rect 20939 47846 20991 47898
rect 21003 47846 21055 47898
rect 21067 47846 21119 47898
rect 1768 47744 1820 47796
rect 2596 47744 2648 47796
rect 13912 47787 13964 47796
rect 13912 47753 13921 47787
rect 13921 47753 13955 47787
rect 13955 47753 13964 47787
rect 13912 47744 13964 47753
rect 17684 47744 17736 47796
rect 17868 47744 17920 47796
rect 18512 47787 18564 47796
rect 2504 47676 2556 47728
rect 1584 47651 1636 47660
rect 1584 47617 1593 47651
rect 1593 47617 1627 47651
rect 1627 47617 1636 47651
rect 1584 47608 1636 47617
rect 2228 47651 2280 47660
rect 2228 47617 2237 47651
rect 2237 47617 2271 47651
rect 2271 47617 2280 47651
rect 2228 47608 2280 47617
rect 14740 47676 14792 47728
rect 18512 47753 18521 47787
rect 18521 47753 18555 47787
rect 18555 47753 18564 47787
rect 18512 47744 18564 47753
rect 25964 47787 26016 47796
rect 25964 47753 25973 47787
rect 25973 47753 26007 47787
rect 26007 47753 26016 47787
rect 25964 47744 26016 47753
rect 26056 47676 26108 47728
rect 29000 47676 29052 47728
rect 30012 47719 30064 47728
rect 30012 47685 30021 47719
rect 30021 47685 30055 47719
rect 30055 47685 30064 47719
rect 30012 47676 30064 47685
rect 14464 47608 14516 47660
rect 16764 47608 16816 47660
rect 14556 47540 14608 47592
rect 17316 47608 17368 47660
rect 17480 47651 17532 47660
rect 17480 47617 17509 47651
rect 17509 47617 17532 47651
rect 17480 47608 17532 47617
rect 18328 47651 18380 47660
rect 14096 47472 14148 47524
rect 14648 47515 14700 47524
rect 14648 47481 14657 47515
rect 14657 47481 14691 47515
rect 14691 47481 14700 47515
rect 14648 47472 14700 47481
rect 17592 47472 17644 47524
rect 17684 47472 17736 47524
rect 18328 47617 18337 47651
rect 18337 47617 18371 47651
rect 18371 47617 18380 47651
rect 18328 47608 18380 47617
rect 17960 47540 18012 47592
rect 19984 47608 20036 47660
rect 26148 47651 26200 47660
rect 26148 47617 26157 47651
rect 26157 47617 26191 47651
rect 26191 47617 26200 47651
rect 26148 47608 26200 47617
rect 25228 47540 25280 47592
rect 27252 47540 27304 47592
rect 27528 47540 27580 47592
rect 19800 47472 19852 47524
rect 19156 47447 19208 47456
rect 19156 47413 19165 47447
rect 19165 47413 19199 47447
rect 19199 47413 19208 47447
rect 19156 47404 19208 47413
rect 20720 47404 20772 47456
rect 25504 47404 25556 47456
rect 26424 47404 26476 47456
rect 28356 47404 28408 47456
rect 5915 47302 5967 47354
rect 5979 47302 6031 47354
rect 6043 47302 6095 47354
rect 6107 47302 6159 47354
rect 6171 47302 6223 47354
rect 15846 47302 15898 47354
rect 15910 47302 15962 47354
rect 15974 47302 16026 47354
rect 16038 47302 16090 47354
rect 16102 47302 16154 47354
rect 25776 47302 25828 47354
rect 25840 47302 25892 47354
rect 25904 47302 25956 47354
rect 25968 47302 26020 47354
rect 26032 47302 26084 47354
rect 14372 47200 14424 47252
rect 1584 47039 1636 47048
rect 1584 47005 1593 47039
rect 1593 47005 1627 47039
rect 1627 47005 1636 47039
rect 1584 46996 1636 47005
rect 2412 46996 2464 47048
rect 14372 46996 14424 47048
rect 14648 47039 14700 47048
rect 14648 47005 14657 47039
rect 14657 47005 14691 47039
rect 14691 47005 14700 47039
rect 14648 46996 14700 47005
rect 14924 47039 14976 47048
rect 14924 47005 14958 47039
rect 14958 47005 14976 47039
rect 14924 46996 14976 47005
rect 14740 46928 14792 46980
rect 17500 47200 17552 47252
rect 20536 47200 20588 47252
rect 23480 47243 23532 47252
rect 23480 47209 23489 47243
rect 23489 47209 23523 47243
rect 23523 47209 23532 47243
rect 23480 47200 23532 47209
rect 24032 47200 24084 47252
rect 26608 47200 26660 47252
rect 17040 47132 17092 47184
rect 19248 47132 19300 47184
rect 19616 47132 19668 47184
rect 22560 47132 22612 47184
rect 24768 47132 24820 47184
rect 26056 47132 26108 47184
rect 17316 47107 17368 47116
rect 17316 47073 17325 47107
rect 17325 47073 17359 47107
rect 17359 47073 17368 47107
rect 17316 47064 17368 47073
rect 27252 47132 27304 47184
rect 18144 46996 18196 47048
rect 19340 46996 19392 47048
rect 26148 47064 26200 47116
rect 26608 47064 26660 47116
rect 27160 47064 27212 47116
rect 27896 47064 27948 47116
rect 30748 47064 30800 47116
rect 30932 47064 30984 47116
rect 22284 47039 22336 47048
rect 2228 46860 2280 46912
rect 2320 46860 2372 46912
rect 17224 46928 17276 46980
rect 20536 46928 20588 46980
rect 21180 46928 21232 46980
rect 22284 47005 22293 47039
rect 22293 47005 22327 47039
rect 22327 47005 22336 47039
rect 22284 46996 22336 47005
rect 22560 46996 22612 47048
rect 22744 46996 22796 47048
rect 23112 46996 23164 47048
rect 27528 46996 27580 47048
rect 28724 47039 28776 47048
rect 28724 47005 28733 47039
rect 28733 47005 28767 47039
rect 28767 47005 28776 47039
rect 28724 46996 28776 47005
rect 20076 46903 20128 46912
rect 20076 46869 20085 46903
rect 20085 46869 20119 46903
rect 20119 46869 20128 46903
rect 20076 46860 20128 46869
rect 22376 46903 22428 46912
rect 22376 46869 22385 46903
rect 22385 46869 22419 46903
rect 22419 46869 22428 46903
rect 22376 46860 22428 46869
rect 23020 46860 23072 46912
rect 23388 46860 23440 46912
rect 24768 46928 24820 46980
rect 26148 46928 26200 46980
rect 29736 46971 29788 46980
rect 29736 46937 29745 46971
rect 29745 46937 29779 46971
rect 29779 46937 29788 46971
rect 29736 46928 29788 46937
rect 30748 46928 30800 46980
rect 26516 46860 26568 46912
rect 27528 46860 27580 46912
rect 28356 46860 28408 46912
rect 10880 46758 10932 46810
rect 10944 46758 10996 46810
rect 11008 46758 11060 46810
rect 11072 46758 11124 46810
rect 11136 46758 11188 46810
rect 20811 46758 20863 46810
rect 20875 46758 20927 46810
rect 20939 46758 20991 46810
rect 21003 46758 21055 46810
rect 21067 46758 21119 46810
rect 13176 46699 13228 46708
rect 13176 46665 13185 46699
rect 13185 46665 13219 46699
rect 13219 46665 13228 46699
rect 13176 46656 13228 46665
rect 14188 46656 14240 46708
rect 16488 46656 16540 46708
rect 19064 46699 19116 46708
rect 19064 46665 19073 46699
rect 19073 46665 19107 46699
rect 19107 46665 19116 46699
rect 19064 46656 19116 46665
rect 24952 46656 25004 46708
rect 26516 46656 26568 46708
rect 28724 46656 28776 46708
rect 28908 46656 28960 46708
rect 12808 46588 12860 46640
rect 14464 46631 14516 46640
rect 14464 46597 14473 46631
rect 14473 46597 14507 46631
rect 14507 46597 14516 46631
rect 14464 46588 14516 46597
rect 14740 46588 14792 46640
rect 15568 46588 15620 46640
rect 19432 46588 19484 46640
rect 21272 46631 21324 46640
rect 21272 46597 21281 46631
rect 21281 46597 21315 46631
rect 21315 46597 21324 46631
rect 21272 46588 21324 46597
rect 1400 46520 1452 46572
rect 11888 46563 11940 46572
rect 11888 46529 11897 46563
rect 11897 46529 11931 46563
rect 11931 46529 11940 46563
rect 11888 46520 11940 46529
rect 15660 46520 15712 46572
rect 16212 46520 16264 46572
rect 17960 46563 18012 46572
rect 17960 46529 17969 46563
rect 17969 46529 18003 46563
rect 18003 46529 18012 46563
rect 17960 46520 18012 46529
rect 18880 46563 18932 46572
rect 18880 46529 18889 46563
rect 18889 46529 18923 46563
rect 18923 46529 18932 46563
rect 18880 46520 18932 46529
rect 23388 46588 23440 46640
rect 22376 46520 22428 46572
rect 22744 46520 22796 46572
rect 22928 46520 22980 46572
rect 23112 46520 23164 46572
rect 23480 46563 23532 46572
rect 23480 46529 23489 46563
rect 23489 46529 23523 46563
rect 23523 46529 23532 46563
rect 23480 46520 23532 46529
rect 28816 46520 28868 46572
rect 29736 46563 29788 46572
rect 29736 46529 29745 46563
rect 29745 46529 29779 46563
rect 29779 46529 29788 46563
rect 29736 46520 29788 46529
rect 14556 46452 14608 46504
rect 16304 46452 16356 46504
rect 22468 46452 22520 46504
rect 14832 46384 14884 46436
rect 15476 46427 15528 46436
rect 15476 46393 15485 46427
rect 15485 46393 15519 46427
rect 15519 46393 15528 46427
rect 15476 46384 15528 46393
rect 18328 46384 18380 46436
rect 23112 46384 23164 46436
rect 23296 46384 23348 46436
rect 25504 46495 25556 46504
rect 25504 46461 25513 46495
rect 25513 46461 25547 46495
rect 25547 46461 25556 46495
rect 25780 46495 25832 46504
rect 25504 46452 25556 46461
rect 25780 46461 25789 46495
rect 25789 46461 25823 46495
rect 25823 46461 25832 46495
rect 25780 46452 25832 46461
rect 26056 46452 26108 46504
rect 26516 46452 26568 46504
rect 2412 46316 2464 46368
rect 13820 46316 13872 46368
rect 14004 46316 14056 46368
rect 21456 46316 21508 46368
rect 22192 46359 22244 46368
rect 22192 46325 22201 46359
rect 22201 46325 22235 46359
rect 22235 46325 22244 46359
rect 22192 46316 22244 46325
rect 23020 46316 23072 46368
rect 25504 46316 25556 46368
rect 29092 46359 29144 46368
rect 29092 46325 29101 46359
rect 29101 46325 29135 46359
rect 29135 46325 29144 46359
rect 29092 46316 29144 46325
rect 31116 46316 31168 46368
rect 5915 46214 5967 46266
rect 5979 46214 6031 46266
rect 6043 46214 6095 46266
rect 6107 46214 6159 46266
rect 6171 46214 6223 46266
rect 15846 46214 15898 46266
rect 15910 46214 15962 46266
rect 15974 46214 16026 46266
rect 16038 46214 16090 46266
rect 16102 46214 16154 46266
rect 25776 46214 25828 46266
rect 25840 46214 25892 46266
rect 25904 46214 25956 46266
rect 25968 46214 26020 46266
rect 26032 46214 26084 46266
rect 30932 46248 30984 46300
rect 31392 46248 31444 46300
rect 12900 46112 12952 46164
rect 14648 46155 14700 46164
rect 14648 46121 14657 46155
rect 14657 46121 14691 46155
rect 14691 46121 14700 46155
rect 14648 46112 14700 46121
rect 19892 46112 19944 46164
rect 22284 46155 22336 46164
rect 22284 46121 22293 46155
rect 22293 46121 22327 46155
rect 22327 46121 22336 46155
rect 22284 46112 22336 46121
rect 1492 45908 1544 45960
rect 2228 45908 2280 45960
rect 12624 46044 12676 46096
rect 13268 46044 13320 46096
rect 14372 46044 14424 46096
rect 17960 46044 18012 46096
rect 22836 46112 22888 46164
rect 23388 46112 23440 46164
rect 26884 46112 26936 46164
rect 27252 46112 27304 46164
rect 29368 46112 29420 46164
rect 31760 46112 31812 46164
rect 25228 46044 25280 46096
rect 25412 46044 25464 46096
rect 31024 46044 31076 46096
rect 31852 46044 31904 46096
rect 12440 45976 12492 46028
rect 13820 45976 13872 46028
rect 2320 45883 2372 45892
rect 2320 45849 2329 45883
rect 2329 45849 2363 45883
rect 2363 45849 2372 45883
rect 2320 45840 2372 45849
rect 11520 45840 11572 45892
rect 12164 45883 12216 45892
rect 12164 45849 12173 45883
rect 12173 45849 12207 45883
rect 12207 45849 12216 45883
rect 12164 45840 12216 45849
rect 12716 45840 12768 45892
rect 1400 45815 1452 45824
rect 1400 45781 1409 45815
rect 1409 45781 1443 45815
rect 1443 45781 1452 45815
rect 1400 45772 1452 45781
rect 2228 45772 2280 45824
rect 2504 45772 2556 45824
rect 2688 45815 2740 45824
rect 2688 45781 2697 45815
rect 2697 45781 2731 45815
rect 2731 45781 2740 45815
rect 2688 45772 2740 45781
rect 10048 45772 10100 45824
rect 11704 45772 11756 45824
rect 11980 45772 12032 45824
rect 12900 45772 12952 45824
rect 13268 45908 13320 45960
rect 18880 45976 18932 46028
rect 20720 45976 20772 46028
rect 21916 45976 21968 46028
rect 22192 45908 22244 45960
rect 15200 45840 15252 45892
rect 15752 45883 15804 45892
rect 15752 45849 15761 45883
rect 15761 45849 15795 45883
rect 15795 45849 15804 45883
rect 15752 45840 15804 45849
rect 18236 45840 18288 45892
rect 19892 45883 19944 45892
rect 19892 45849 19901 45883
rect 19901 45849 19935 45883
rect 19935 45849 19944 45883
rect 19892 45840 19944 45849
rect 22468 45976 22520 46028
rect 22836 45976 22888 46028
rect 23020 45951 23072 45960
rect 23020 45917 23029 45951
rect 23029 45917 23063 45951
rect 23063 45917 23072 45951
rect 23020 45908 23072 45917
rect 25044 45976 25096 46028
rect 25688 45976 25740 46028
rect 13268 45772 13320 45824
rect 16948 45772 17000 45824
rect 17408 45772 17460 45824
rect 25412 45840 25464 45892
rect 29184 45908 29236 45960
rect 29368 45908 29420 45960
rect 29736 45951 29788 45960
rect 29736 45917 29745 45951
rect 29745 45917 29779 45951
rect 29779 45917 29788 45951
rect 29736 45908 29788 45917
rect 30012 45951 30064 45960
rect 30012 45917 30021 45951
rect 30021 45917 30055 45951
rect 30055 45917 30064 45951
rect 30012 45908 30064 45917
rect 28356 45840 28408 45892
rect 23020 45772 23072 45824
rect 23296 45772 23348 45824
rect 23756 45772 23808 45824
rect 24032 45772 24084 45824
rect 25320 45772 25372 45824
rect 25688 45772 25740 45824
rect 29184 45772 29236 45824
rect 10880 45670 10932 45722
rect 10944 45670 10996 45722
rect 11008 45670 11060 45722
rect 11072 45670 11124 45722
rect 11136 45670 11188 45722
rect 20811 45670 20863 45722
rect 20875 45670 20927 45722
rect 20939 45670 20991 45722
rect 21003 45670 21055 45722
rect 21067 45670 21119 45722
rect 2688 45568 2740 45620
rect 14004 45568 14056 45620
rect 15752 45568 15804 45620
rect 20352 45568 20404 45620
rect 24676 45568 24728 45620
rect 2320 45543 2372 45552
rect 2320 45509 2329 45543
rect 2329 45509 2363 45543
rect 2363 45509 2372 45543
rect 2320 45500 2372 45509
rect 2412 45500 2464 45552
rect 12532 45543 12584 45552
rect 12532 45509 12541 45543
rect 12541 45509 12575 45543
rect 12575 45509 12584 45543
rect 12532 45500 12584 45509
rect 12808 45500 12860 45552
rect 1584 45475 1636 45484
rect 1584 45441 1593 45475
rect 1593 45441 1627 45475
rect 1627 45441 1636 45475
rect 1584 45432 1636 45441
rect 13268 45500 13320 45552
rect 16948 45500 17000 45552
rect 18420 45500 18472 45552
rect 13728 45475 13780 45484
rect 12532 45364 12584 45416
rect 7472 45296 7524 45348
rect 13728 45441 13737 45475
rect 13737 45441 13771 45475
rect 13771 45441 13780 45475
rect 13728 45432 13780 45441
rect 14188 45432 14240 45484
rect 18512 45432 18564 45484
rect 13360 45296 13412 45348
rect 19984 45339 20036 45348
rect 19984 45305 19993 45339
rect 19993 45305 20027 45339
rect 20027 45305 20036 45339
rect 19984 45296 20036 45305
rect 21180 45500 21232 45552
rect 22100 45500 22152 45552
rect 22652 45500 22704 45552
rect 24768 45500 24820 45552
rect 25320 45568 25372 45620
rect 24952 45500 25004 45552
rect 25504 45500 25556 45552
rect 28908 45568 28960 45620
rect 26424 45500 26476 45552
rect 27804 45500 27856 45552
rect 20720 45432 20772 45484
rect 21916 45475 21968 45484
rect 21916 45441 21925 45475
rect 21925 45441 21959 45475
rect 21959 45441 21968 45475
rect 21916 45432 21968 45441
rect 22468 45432 22520 45484
rect 23756 45432 23808 45484
rect 20904 45364 20956 45416
rect 20996 45364 21048 45416
rect 24032 45407 24084 45416
rect 24032 45373 24041 45407
rect 24041 45373 24075 45407
rect 24075 45373 24084 45407
rect 24032 45364 24084 45373
rect 28356 45432 28408 45484
rect 29736 45500 29788 45552
rect 29552 45475 29604 45484
rect 29552 45441 29561 45475
rect 29561 45441 29595 45475
rect 29595 45441 29604 45475
rect 29552 45432 29604 45441
rect 24768 45364 24820 45416
rect 25044 45364 25096 45416
rect 25320 45364 25372 45416
rect 28540 45364 28592 45416
rect 30012 45364 30064 45416
rect 1768 45228 1820 45280
rect 12624 45228 12676 45280
rect 19524 45228 19576 45280
rect 22468 45228 22520 45280
rect 24676 45228 24728 45280
rect 24952 45271 25004 45280
rect 24952 45237 24961 45271
rect 24961 45237 24995 45271
rect 24995 45237 25004 45271
rect 24952 45228 25004 45237
rect 29276 45296 29328 45348
rect 31852 45704 31904 45756
rect 28908 45228 28960 45280
rect 29092 45228 29144 45280
rect 31760 45228 31812 45280
rect 5915 45126 5967 45178
rect 5979 45126 6031 45178
rect 6043 45126 6095 45178
rect 6107 45126 6159 45178
rect 6171 45126 6223 45178
rect 15846 45126 15898 45178
rect 15910 45126 15962 45178
rect 15974 45126 16026 45178
rect 16038 45126 16090 45178
rect 16102 45126 16154 45178
rect 25776 45126 25828 45178
rect 25840 45126 25892 45178
rect 25904 45126 25956 45178
rect 25968 45126 26020 45178
rect 26032 45126 26084 45178
rect 7472 45024 7524 45076
rect 12256 45024 12308 45076
rect 16764 45024 16816 45076
rect 16948 45024 17000 45076
rect 22284 45024 22336 45076
rect 28724 45024 28776 45076
rect 10048 44931 10100 44940
rect 10048 44897 10057 44931
rect 10057 44897 10091 44931
rect 10091 44897 10100 44931
rect 10048 44888 10100 44897
rect 1400 44820 1452 44872
rect 13084 44956 13136 45008
rect 19432 44956 19484 45008
rect 20904 44956 20956 45008
rect 12900 44888 12952 44940
rect 19800 44931 19852 44940
rect 19800 44897 19809 44931
rect 19809 44897 19843 44931
rect 19843 44897 19852 44931
rect 19800 44888 19852 44897
rect 20996 44931 21048 44940
rect 20996 44897 21005 44931
rect 21005 44897 21039 44931
rect 21039 44897 21048 44931
rect 20996 44888 21048 44897
rect 24492 44956 24544 45008
rect 26332 44956 26384 45008
rect 29092 44956 29144 45008
rect 29276 44956 29328 45008
rect 29644 44956 29696 45008
rect 31852 44956 31904 45008
rect 25044 44931 25096 44940
rect 1676 44752 1728 44804
rect 9772 44752 9824 44804
rect 12992 44820 13044 44872
rect 13360 44863 13412 44872
rect 13360 44829 13369 44863
rect 13369 44829 13403 44863
rect 13403 44829 13412 44863
rect 13360 44820 13412 44829
rect 13912 44820 13964 44872
rect 17132 44820 17184 44872
rect 19340 44820 19392 44872
rect 25044 44897 25053 44931
rect 25053 44897 25087 44931
rect 25087 44897 25096 44931
rect 25044 44888 25096 44897
rect 25320 44888 25372 44940
rect 28356 44888 28408 44940
rect 28908 44888 28960 44940
rect 12532 44752 12584 44804
rect 15292 44752 15344 44804
rect 17868 44752 17920 44804
rect 19984 44752 20036 44804
rect 20628 44752 20680 44804
rect 10416 44684 10468 44736
rect 13268 44684 13320 44736
rect 14648 44684 14700 44736
rect 15752 44727 15804 44736
rect 15752 44693 15761 44727
rect 15761 44693 15795 44727
rect 15795 44693 15804 44727
rect 15752 44684 15804 44693
rect 21180 44684 21232 44736
rect 22652 44820 22704 44872
rect 23664 44820 23716 44872
rect 23756 44820 23808 44872
rect 24492 44820 24544 44872
rect 27160 44863 27212 44872
rect 22376 44752 22428 44804
rect 24768 44752 24820 44804
rect 27160 44829 27169 44863
rect 27169 44829 27203 44863
rect 27203 44829 27212 44863
rect 27160 44820 27212 44829
rect 28264 44863 28316 44872
rect 28264 44829 28273 44863
rect 28273 44829 28307 44863
rect 28307 44829 28316 44863
rect 28264 44820 28316 44829
rect 28724 44863 28776 44872
rect 28724 44829 28733 44863
rect 28733 44829 28767 44863
rect 28767 44829 28776 44863
rect 28724 44820 28776 44829
rect 29736 44863 29788 44872
rect 29736 44829 29745 44863
rect 29745 44829 29779 44863
rect 29779 44829 29788 44863
rect 29736 44820 29788 44829
rect 30012 44863 30064 44872
rect 30012 44829 30021 44863
rect 30021 44829 30055 44863
rect 30055 44829 30064 44863
rect 30012 44820 30064 44829
rect 22652 44684 22704 44736
rect 23664 44684 23716 44736
rect 25044 44684 25096 44736
rect 25136 44684 25188 44736
rect 26884 44684 26936 44736
rect 28908 44727 28960 44736
rect 28908 44693 28917 44727
rect 28917 44693 28951 44727
rect 28951 44693 28960 44727
rect 28908 44684 28960 44693
rect 29644 44684 29696 44736
rect 10880 44582 10932 44634
rect 10944 44582 10996 44634
rect 11008 44582 11060 44634
rect 11072 44582 11124 44634
rect 11136 44582 11188 44634
rect 20811 44582 20863 44634
rect 20875 44582 20927 44634
rect 20939 44582 20991 44634
rect 21003 44582 21055 44634
rect 21067 44582 21119 44634
rect 1676 44412 1728 44464
rect 2596 44480 2648 44532
rect 2780 44344 2832 44396
rect 12348 44480 12400 44532
rect 12440 44480 12492 44532
rect 14740 44480 14792 44532
rect 17776 44480 17828 44532
rect 19892 44480 19944 44532
rect 20628 44480 20680 44532
rect 23664 44480 23716 44532
rect 24492 44523 24544 44532
rect 24492 44489 24501 44523
rect 24501 44489 24535 44523
rect 24535 44489 24544 44523
rect 24492 44480 24544 44489
rect 27160 44480 27212 44532
rect 27436 44480 27488 44532
rect 30012 44480 30064 44532
rect 11704 44412 11756 44464
rect 11612 44344 11664 44396
rect 12072 44387 12124 44396
rect 12072 44353 12081 44387
rect 12081 44353 12115 44387
rect 12115 44353 12124 44387
rect 12072 44344 12124 44353
rect 12808 44412 12860 44464
rect 13176 44412 13228 44464
rect 14188 44455 14240 44464
rect 14188 44421 14197 44455
rect 14197 44421 14231 44455
rect 14231 44421 14240 44455
rect 14188 44412 14240 44421
rect 11796 44319 11848 44328
rect 11796 44285 11805 44319
rect 11805 44285 11839 44319
rect 11839 44285 11848 44319
rect 11796 44276 11848 44285
rect 12532 44344 12584 44396
rect 15476 44412 15528 44464
rect 15660 44412 15712 44464
rect 16304 44412 16356 44464
rect 17224 44455 17276 44464
rect 17224 44421 17233 44455
rect 17233 44421 17267 44455
rect 17267 44421 17276 44455
rect 17224 44412 17276 44421
rect 17684 44412 17736 44464
rect 19524 44455 19576 44464
rect 19524 44421 19533 44455
rect 19533 44421 19567 44455
rect 19567 44421 19576 44455
rect 19524 44412 19576 44421
rect 21272 44412 21324 44464
rect 23296 44412 23348 44464
rect 12716 44276 12768 44328
rect 18052 44344 18104 44396
rect 17132 44319 17184 44328
rect 12072 44208 12124 44260
rect 13544 44208 13596 44260
rect 15384 44208 15436 44260
rect 17132 44285 17141 44319
rect 17141 44285 17175 44319
rect 17175 44285 17184 44319
rect 17132 44276 17184 44285
rect 17592 44276 17644 44328
rect 18328 44387 18380 44396
rect 18328 44353 18337 44387
rect 18337 44353 18371 44387
rect 18371 44353 18380 44387
rect 18328 44344 18380 44353
rect 18604 44344 18656 44396
rect 22744 44344 22796 44396
rect 19248 44276 19300 44328
rect 19524 44276 19576 44328
rect 16580 44208 16632 44260
rect 24676 44412 24728 44464
rect 28356 44412 28408 44464
rect 23756 44344 23808 44396
rect 25504 44344 25556 44396
rect 26884 44344 26936 44396
rect 27988 44387 28040 44396
rect 27988 44353 27997 44387
rect 27997 44353 28031 44387
rect 28031 44353 28040 44387
rect 27988 44344 28040 44353
rect 28264 44344 28316 44396
rect 28540 44344 28592 44396
rect 28816 44344 28868 44396
rect 29828 44387 29880 44396
rect 29828 44353 29837 44387
rect 29837 44353 29871 44387
rect 29871 44353 29880 44387
rect 29828 44344 29880 44353
rect 25320 44276 25372 44328
rect 24492 44208 24544 44260
rect 30012 44251 30064 44260
rect 30012 44217 30021 44251
rect 30021 44217 30055 44251
rect 30055 44217 30064 44251
rect 30012 44208 30064 44217
rect 12992 44140 13044 44192
rect 17684 44140 17736 44192
rect 18052 44140 18104 44192
rect 18788 44140 18840 44192
rect 20996 44140 21048 44192
rect 23296 44140 23348 44192
rect 5915 44038 5967 44090
rect 5979 44038 6031 44090
rect 6043 44038 6095 44090
rect 6107 44038 6159 44090
rect 6171 44038 6223 44090
rect 15846 44038 15898 44090
rect 15910 44038 15962 44090
rect 15974 44038 16026 44090
rect 16038 44038 16090 44090
rect 16102 44038 16154 44090
rect 25776 44038 25828 44090
rect 25840 44038 25892 44090
rect 25904 44038 25956 44090
rect 25968 44038 26020 44090
rect 26032 44038 26084 44090
rect 12532 43936 12584 43988
rect 13728 43936 13780 43988
rect 15200 43936 15252 43988
rect 16580 43936 16632 43988
rect 17776 43936 17828 43988
rect 19708 43936 19760 43988
rect 24308 43936 24360 43988
rect 26332 43936 26384 43988
rect 9680 43868 9732 43920
rect 12716 43868 12768 43920
rect 12992 43868 13044 43920
rect 19156 43868 19208 43920
rect 19892 43868 19944 43920
rect 23756 43868 23808 43920
rect 1768 43775 1820 43784
rect 1768 43741 1777 43775
rect 1777 43741 1811 43775
rect 1811 43741 1820 43775
rect 1768 43732 1820 43741
rect 10416 43800 10468 43852
rect 12348 43800 12400 43852
rect 1676 43664 1728 43716
rect 2596 43707 2648 43716
rect 2596 43673 2605 43707
rect 2605 43673 2639 43707
rect 2639 43673 2648 43707
rect 2596 43664 2648 43673
rect 9772 43664 9824 43716
rect 10140 43772 10192 43781
rect 10140 43738 10149 43772
rect 10149 43738 10183 43772
rect 10183 43738 10192 43772
rect 10324 43775 10376 43784
rect 10140 43729 10192 43738
rect 10324 43741 10333 43775
rect 10333 43741 10367 43775
rect 10367 43741 10376 43775
rect 10324 43732 10376 43741
rect 14372 43800 14424 43852
rect 14556 43800 14608 43852
rect 17132 43800 17184 43852
rect 19800 43843 19852 43852
rect 19800 43809 19809 43843
rect 19809 43809 19843 43843
rect 19843 43809 19852 43843
rect 20996 43843 21048 43852
rect 19800 43800 19852 43809
rect 20996 43809 21005 43843
rect 21005 43809 21039 43843
rect 21039 43809 21048 43843
rect 20996 43800 21048 43809
rect 23664 43800 23716 43852
rect 11520 43664 11572 43716
rect 12808 43732 12860 43784
rect 13084 43732 13136 43784
rect 14188 43732 14240 43784
rect 16304 43732 16356 43784
rect 16396 43732 16448 43784
rect 14096 43664 14148 43716
rect 14464 43707 14516 43716
rect 14464 43673 14473 43707
rect 14473 43673 14507 43707
rect 14507 43673 14516 43707
rect 14464 43664 14516 43673
rect 14648 43707 14700 43716
rect 14648 43673 14657 43707
rect 14657 43673 14691 43707
rect 14691 43673 14700 43707
rect 14648 43664 14700 43673
rect 15568 43664 15620 43716
rect 19248 43664 19300 43716
rect 19984 43732 20036 43784
rect 22008 43775 22060 43784
rect 22008 43741 22017 43775
rect 22017 43741 22051 43775
rect 22051 43741 22060 43775
rect 22008 43732 22060 43741
rect 22468 43775 22520 43784
rect 22468 43741 22477 43775
rect 22477 43741 22511 43775
rect 22511 43741 22520 43775
rect 22468 43732 22520 43741
rect 23756 43775 23808 43784
rect 23756 43741 23765 43775
rect 23765 43741 23799 43775
rect 23799 43741 23808 43775
rect 23756 43732 23808 43741
rect 24492 43800 24544 43852
rect 24676 43843 24728 43852
rect 24676 43809 24685 43843
rect 24685 43809 24719 43843
rect 24719 43809 24728 43843
rect 24676 43800 24728 43809
rect 28264 43843 28316 43852
rect 28264 43809 28273 43843
rect 28273 43809 28307 43843
rect 28307 43809 28316 43843
rect 28264 43800 28316 43809
rect 24032 43732 24084 43784
rect 24768 43732 24820 43784
rect 26884 43732 26936 43784
rect 28356 43732 28408 43784
rect 29828 43775 29880 43784
rect 29828 43741 29837 43775
rect 29837 43741 29871 43775
rect 29871 43741 29880 43775
rect 29828 43732 29880 43741
rect 1952 43639 2004 43648
rect 1952 43605 1961 43639
rect 1961 43605 1995 43639
rect 1995 43605 2004 43639
rect 1952 43596 2004 43605
rect 9956 43596 10008 43648
rect 12164 43596 12216 43648
rect 13084 43596 13136 43648
rect 20168 43596 20220 43648
rect 22192 43596 22244 43648
rect 23756 43596 23808 43648
rect 28264 43664 28316 43716
rect 25136 43596 25188 43648
rect 26424 43596 26476 43648
rect 30012 43639 30064 43648
rect 30012 43605 30021 43639
rect 30021 43605 30055 43639
rect 30055 43605 30064 43639
rect 30012 43596 30064 43605
rect 10880 43494 10932 43546
rect 10944 43494 10996 43546
rect 11008 43494 11060 43546
rect 11072 43494 11124 43546
rect 11136 43494 11188 43546
rect 20811 43494 20863 43546
rect 20875 43494 20927 43546
rect 20939 43494 20991 43546
rect 21003 43494 21055 43546
rect 21067 43494 21119 43546
rect 9588 43435 9640 43444
rect 9588 43401 9597 43435
rect 9597 43401 9631 43435
rect 9631 43401 9640 43435
rect 9588 43392 9640 43401
rect 9864 43392 9916 43444
rect 9956 43392 10008 43444
rect 18144 43392 18196 43444
rect 19708 43392 19760 43444
rect 20536 43392 20588 43444
rect 24584 43392 24636 43444
rect 1676 43324 1728 43376
rect 1952 43324 2004 43376
rect 9404 43324 9456 43376
rect 1768 43299 1820 43308
rect 1768 43265 1777 43299
rect 1777 43265 1811 43299
rect 1811 43265 1820 43299
rect 1768 43256 1820 43265
rect 2228 43256 2280 43308
rect 2504 43256 2556 43308
rect 10048 43299 10100 43308
rect 10048 43265 10057 43299
rect 10057 43265 10091 43299
rect 10091 43265 10100 43299
rect 10232 43299 10284 43308
rect 10048 43256 10100 43265
rect 10232 43265 10241 43299
rect 10241 43265 10275 43299
rect 10275 43265 10284 43299
rect 10232 43256 10284 43265
rect 12808 43324 12860 43376
rect 14556 43324 14608 43376
rect 19616 43324 19668 43376
rect 13084 43299 13136 43308
rect 13084 43265 13093 43299
rect 13093 43265 13127 43299
rect 13127 43265 13136 43299
rect 13084 43256 13136 43265
rect 15016 43299 15068 43308
rect 15016 43265 15025 43299
rect 15025 43265 15059 43299
rect 15059 43265 15068 43299
rect 15016 43256 15068 43265
rect 15476 43256 15528 43308
rect 16304 43256 16356 43308
rect 17040 43299 17092 43308
rect 17040 43265 17049 43299
rect 17049 43265 17083 43299
rect 17083 43265 17092 43299
rect 17040 43256 17092 43265
rect 12072 43188 12124 43240
rect 12808 43231 12860 43240
rect 12808 43197 12817 43231
rect 12817 43197 12851 43231
rect 12851 43197 12860 43231
rect 12808 43188 12860 43197
rect 13268 43188 13320 43240
rect 10324 43120 10376 43172
rect 14280 43120 14332 43172
rect 15200 43163 15252 43172
rect 15200 43129 15209 43163
rect 15209 43129 15243 43163
rect 15243 43129 15252 43163
rect 15200 43120 15252 43129
rect 20628 43188 20680 43240
rect 25136 43324 25188 43376
rect 29552 43324 29604 43376
rect 29828 43324 29880 43376
rect 30104 43367 30156 43376
rect 30104 43333 30113 43367
rect 30113 43333 30147 43367
rect 30147 43333 30156 43367
rect 30104 43324 30156 43333
rect 23664 43256 23716 43308
rect 24768 43256 24820 43308
rect 25320 43256 25372 43308
rect 24032 43188 24084 43240
rect 24492 43188 24544 43240
rect 14096 43052 14148 43104
rect 16212 43052 16264 43104
rect 21364 43052 21416 43104
rect 22376 43095 22428 43104
rect 22376 43061 22385 43095
rect 22385 43061 22419 43095
rect 22419 43061 22428 43095
rect 22376 43052 22428 43061
rect 23296 43052 23348 43104
rect 23664 43120 23716 43172
rect 24584 43120 24636 43172
rect 25136 43120 25188 43172
rect 25320 43120 25372 43172
rect 29092 43299 29144 43308
rect 29092 43265 29101 43299
rect 29101 43265 29135 43299
rect 29135 43265 29144 43299
rect 29092 43256 29144 43265
rect 29920 43299 29972 43308
rect 29920 43265 29929 43299
rect 29929 43265 29963 43299
rect 29963 43265 29972 43299
rect 29920 43256 29972 43265
rect 30104 43188 30156 43240
rect 24768 43052 24820 43104
rect 26424 43052 26476 43104
rect 27804 43095 27856 43104
rect 27804 43061 27813 43095
rect 27813 43061 27847 43095
rect 27847 43061 27856 43095
rect 27804 43052 27856 43061
rect 27988 43052 28040 43104
rect 29276 43095 29328 43104
rect 29276 43061 29285 43095
rect 29285 43061 29319 43095
rect 29319 43061 29328 43095
rect 29276 43052 29328 43061
rect 29552 43052 29604 43104
rect 5915 42950 5967 43002
rect 5979 42950 6031 43002
rect 6043 42950 6095 43002
rect 6107 42950 6159 43002
rect 6171 42950 6223 43002
rect 15846 42950 15898 43002
rect 15910 42950 15962 43002
rect 15974 42950 16026 43002
rect 16038 42950 16090 43002
rect 16102 42950 16154 43002
rect 25776 42950 25828 43002
rect 25840 42950 25892 43002
rect 25904 42950 25956 43002
rect 25968 42950 26020 43002
rect 26032 42950 26084 43002
rect 1768 42848 1820 42900
rect 2596 42848 2648 42900
rect 12808 42848 12860 42900
rect 23664 42848 23716 42900
rect 14004 42780 14056 42832
rect 24676 42848 24728 42900
rect 1584 42687 1636 42696
rect 1584 42653 1593 42687
rect 1593 42653 1627 42687
rect 1627 42653 1636 42687
rect 1584 42644 1636 42653
rect 2228 42687 2280 42696
rect 2228 42653 2237 42687
rect 2237 42653 2271 42687
rect 2271 42653 2280 42687
rect 2228 42644 2280 42653
rect 9680 42712 9732 42764
rect 11520 42712 11572 42764
rect 15016 42712 15068 42764
rect 15200 42712 15252 42764
rect 10416 42687 10468 42696
rect 10416 42653 10425 42687
rect 10425 42653 10459 42687
rect 10459 42653 10468 42687
rect 10416 42644 10468 42653
rect 14372 42687 14424 42696
rect 11980 42576 12032 42628
rect 14372 42653 14381 42687
rect 14381 42653 14415 42687
rect 14415 42653 14424 42687
rect 14372 42644 14424 42653
rect 15476 42644 15528 42696
rect 15660 42687 15712 42696
rect 15660 42653 15669 42687
rect 15669 42653 15703 42687
rect 15703 42653 15712 42687
rect 15660 42644 15712 42653
rect 17132 42712 17184 42764
rect 21916 42755 21968 42764
rect 21916 42721 21925 42755
rect 21925 42721 21959 42755
rect 21959 42721 21968 42755
rect 21916 42712 21968 42721
rect 23296 42712 23348 42764
rect 24492 42712 24544 42764
rect 24768 42780 24820 42832
rect 15108 42576 15160 42628
rect 18420 42644 18472 42696
rect 20076 42644 20128 42696
rect 22284 42644 22336 42696
rect 28264 42848 28316 42900
rect 28632 42848 28684 42900
rect 29828 42848 29880 42900
rect 25136 42780 25188 42832
rect 25780 42712 25832 42764
rect 25136 42644 25188 42696
rect 18604 42576 18656 42628
rect 25688 42576 25740 42628
rect 25872 42619 25924 42628
rect 25872 42585 25881 42619
rect 25881 42585 25915 42619
rect 25915 42585 25924 42619
rect 25872 42576 25924 42585
rect 26240 42644 26292 42696
rect 28264 42644 28316 42696
rect 28908 42712 28960 42764
rect 12992 42508 13044 42560
rect 15384 42551 15436 42560
rect 15384 42517 15393 42551
rect 15393 42517 15427 42551
rect 15427 42517 15436 42551
rect 15384 42508 15436 42517
rect 16396 42508 16448 42560
rect 18236 42551 18288 42560
rect 18236 42517 18245 42551
rect 18245 42517 18279 42551
rect 18279 42517 18288 42551
rect 18236 42508 18288 42517
rect 18972 42508 19024 42560
rect 22284 42508 22336 42560
rect 22652 42551 22704 42560
rect 22652 42517 22661 42551
rect 22661 42517 22695 42551
rect 22695 42517 22704 42551
rect 22652 42508 22704 42517
rect 24676 42508 24728 42560
rect 25320 42508 25372 42560
rect 25964 42551 26016 42560
rect 25964 42517 25973 42551
rect 25973 42517 26007 42551
rect 26007 42517 26016 42551
rect 25964 42508 26016 42517
rect 26056 42508 26108 42560
rect 28356 42576 28408 42628
rect 28816 42508 28868 42560
rect 29000 42508 29052 42560
rect 29644 42508 29696 42560
rect 29736 42508 29788 42560
rect 10880 42406 10932 42458
rect 10944 42406 10996 42458
rect 11008 42406 11060 42458
rect 11072 42406 11124 42458
rect 11136 42406 11188 42458
rect 20811 42406 20863 42458
rect 20875 42406 20927 42458
rect 20939 42406 20991 42458
rect 21003 42406 21055 42458
rect 21067 42406 21119 42458
rect 10416 42304 10468 42356
rect 11888 42304 11940 42356
rect 14648 42304 14700 42356
rect 15108 42304 15160 42356
rect 17040 42304 17092 42356
rect 19248 42304 19300 42356
rect 21364 42304 21416 42356
rect 23296 42304 23348 42356
rect 25780 42304 25832 42356
rect 14464 42236 14516 42288
rect 1584 42211 1636 42220
rect 1584 42177 1593 42211
rect 1593 42177 1627 42211
rect 1627 42177 1636 42211
rect 1584 42168 1636 42177
rect 8392 42211 8444 42220
rect 8392 42177 8401 42211
rect 8401 42177 8435 42211
rect 8435 42177 8444 42211
rect 8392 42168 8444 42177
rect 9956 42032 10008 42084
rect 10048 42032 10100 42084
rect 10232 42168 10284 42220
rect 15752 42236 15804 42288
rect 16948 42236 17000 42288
rect 14280 42100 14332 42152
rect 14556 42100 14608 42152
rect 16672 42168 16724 42220
rect 17684 42211 17736 42220
rect 17684 42177 17718 42211
rect 17718 42177 17736 42211
rect 17684 42168 17736 42177
rect 20076 42168 20128 42220
rect 22100 42236 22152 42288
rect 22192 42236 22244 42288
rect 10324 42032 10376 42084
rect 12072 42032 12124 42084
rect 16856 42100 16908 42152
rect 17408 42143 17460 42152
rect 17408 42109 17417 42143
rect 17417 42109 17451 42143
rect 17451 42109 17460 42143
rect 17408 42100 17460 42109
rect 18880 42100 18932 42152
rect 20628 42168 20680 42220
rect 26240 42236 26292 42288
rect 26424 42236 26476 42288
rect 27988 42304 28040 42356
rect 29644 42304 29696 42356
rect 29736 42304 29788 42356
rect 30104 42304 30156 42356
rect 27436 42236 27488 42288
rect 27712 42236 27764 42288
rect 25412 42168 25464 42220
rect 26516 42168 26568 42220
rect 17132 42032 17184 42084
rect 18788 42075 18840 42084
rect 18788 42041 18797 42075
rect 18797 42041 18831 42075
rect 18831 42041 18840 42075
rect 18788 42032 18840 42041
rect 11980 41964 12032 42016
rect 14096 42007 14148 42016
rect 14096 41973 14105 42007
rect 14105 41973 14139 42007
rect 14139 41973 14148 42007
rect 14096 41964 14148 41973
rect 16672 41964 16724 42016
rect 18512 41964 18564 42016
rect 19524 41964 19576 42016
rect 20260 41964 20312 42016
rect 21456 41964 21508 42016
rect 25780 42100 25832 42152
rect 24768 42032 24820 42084
rect 25964 42032 26016 42084
rect 26056 42032 26108 42084
rect 26332 42032 26384 42084
rect 26700 42032 26752 42084
rect 27804 42168 27856 42220
rect 28356 42236 28408 42288
rect 28908 42236 28960 42288
rect 28264 42168 28316 42220
rect 28540 42168 28592 42220
rect 27436 42100 27488 42152
rect 29920 42211 29972 42220
rect 29920 42177 29929 42211
rect 29929 42177 29963 42211
rect 29963 42177 29972 42211
rect 29920 42168 29972 42177
rect 31392 42304 31444 42356
rect 30656 42236 30708 42288
rect 30472 42168 30524 42220
rect 24676 41964 24728 42016
rect 25320 41964 25372 42016
rect 27436 41964 27488 42016
rect 27620 42032 27672 42084
rect 28356 42032 28408 42084
rect 29092 42032 29144 42084
rect 27988 41964 28040 42016
rect 29460 42007 29512 42016
rect 29460 41973 29469 42007
rect 29469 41973 29503 42007
rect 29503 41973 29512 42007
rect 29460 41964 29512 41973
rect 29644 42032 29696 42084
rect 29920 42032 29972 42084
rect 30012 41964 30064 42016
rect 5915 41862 5967 41914
rect 5979 41862 6031 41914
rect 6043 41862 6095 41914
rect 6107 41862 6159 41914
rect 6171 41862 6223 41914
rect 15846 41862 15898 41914
rect 15910 41862 15962 41914
rect 15974 41862 16026 41914
rect 16038 41862 16090 41914
rect 16102 41862 16154 41914
rect 25776 41862 25828 41914
rect 25840 41862 25892 41914
rect 25904 41862 25956 41914
rect 25968 41862 26020 41914
rect 26032 41862 26084 41914
rect 10324 41760 10376 41812
rect 12900 41760 12952 41812
rect 15660 41760 15712 41812
rect 17224 41760 17276 41812
rect 18512 41735 18564 41744
rect 12072 41624 12124 41676
rect 18512 41701 18521 41735
rect 18521 41701 18555 41735
rect 18555 41701 18564 41735
rect 18512 41692 18564 41701
rect 20628 41760 20680 41812
rect 21824 41803 21876 41812
rect 21824 41769 21833 41803
rect 21833 41769 21867 41803
rect 21867 41769 21876 41803
rect 21824 41760 21876 41769
rect 22008 41760 22060 41812
rect 22100 41692 22152 41744
rect 22192 41692 22244 41744
rect 17776 41624 17828 41676
rect 1584 41599 1636 41608
rect 1584 41565 1593 41599
rect 1593 41565 1627 41599
rect 1627 41565 1636 41599
rect 1584 41556 1636 41565
rect 8392 41556 8444 41608
rect 10048 41556 10100 41608
rect 14096 41599 14148 41608
rect 14096 41565 14105 41599
rect 14105 41565 14139 41599
rect 14139 41565 14148 41599
rect 14096 41556 14148 41565
rect 15384 41556 15436 41608
rect 17960 41556 18012 41608
rect 19340 41624 19392 41676
rect 20168 41624 20220 41676
rect 25320 41624 25372 41676
rect 27988 41760 28040 41812
rect 28816 41760 28868 41812
rect 29828 41760 29880 41812
rect 25964 41692 26016 41744
rect 26424 41735 26476 41744
rect 26424 41701 26433 41735
rect 26433 41701 26467 41735
rect 26467 41701 26476 41735
rect 26424 41692 26476 41701
rect 30564 41760 30616 41812
rect 25688 41667 25740 41676
rect 25688 41633 25697 41667
rect 25697 41633 25731 41667
rect 25731 41633 25740 41667
rect 25688 41624 25740 41633
rect 19892 41556 19944 41608
rect 20720 41556 20772 41608
rect 12348 41488 12400 41540
rect 18236 41488 18288 41540
rect 19708 41531 19760 41540
rect 19708 41497 19717 41531
rect 19717 41497 19751 41531
rect 19751 41497 19760 41531
rect 19708 41488 19760 41497
rect 20076 41488 20128 41540
rect 23572 41599 23624 41608
rect 23572 41565 23581 41599
rect 23581 41565 23615 41599
rect 23615 41565 23624 41599
rect 23572 41556 23624 41565
rect 24768 41556 24820 41608
rect 24032 41488 24084 41540
rect 24308 41488 24360 41540
rect 27528 41556 27580 41608
rect 28172 41556 28224 41608
rect 25136 41488 25188 41540
rect 18144 41420 18196 41472
rect 19524 41420 19576 41472
rect 20720 41420 20772 41472
rect 24860 41420 24912 41472
rect 25504 41488 25556 41540
rect 26056 41488 26108 41540
rect 27712 41488 27764 41540
rect 25780 41420 25832 41472
rect 26516 41420 26568 41472
rect 27988 41420 28040 41472
rect 28540 41556 28592 41608
rect 28724 41559 28733 41586
rect 28733 41559 28767 41586
rect 28767 41559 28776 41586
rect 28724 41534 28776 41559
rect 28816 41596 28868 41608
rect 28816 41562 28825 41596
rect 28825 41562 28859 41596
rect 28859 41562 28868 41596
rect 29184 41624 29236 41676
rect 28816 41556 28868 41562
rect 29920 41599 29972 41608
rect 29920 41565 29929 41599
rect 29929 41565 29963 41599
rect 29963 41565 29972 41599
rect 29920 41556 29972 41565
rect 30104 41556 30156 41608
rect 29092 41420 29144 41472
rect 30104 41420 30156 41472
rect 30288 41420 30340 41472
rect 31116 41488 31168 41540
rect 31392 41760 31444 41812
rect 30472 41420 30524 41472
rect 30656 41420 30708 41472
rect 30840 41420 30892 41472
rect 10880 41318 10932 41370
rect 10944 41318 10996 41370
rect 11008 41318 11060 41370
rect 11072 41318 11124 41370
rect 11136 41318 11188 41370
rect 20811 41318 20863 41370
rect 20875 41318 20927 41370
rect 20939 41318 20991 41370
rect 21003 41318 21055 41370
rect 21067 41318 21119 41370
rect 31116 41352 31168 41404
rect 15292 41216 15344 41268
rect 17592 41216 17644 41268
rect 18604 41259 18656 41268
rect 18604 41225 18613 41259
rect 18613 41225 18647 41259
rect 18647 41225 18656 41259
rect 18604 41216 18656 41225
rect 19984 41216 20036 41268
rect 1860 41148 1912 41200
rect 1584 41123 1636 41132
rect 1584 41089 1593 41123
rect 1593 41089 1627 41123
rect 1627 41089 1636 41123
rect 1584 41080 1636 41089
rect 16396 41148 16448 41200
rect 16672 41123 16724 41132
rect 15752 41012 15804 41064
rect 16672 41089 16681 41123
rect 16681 41089 16715 41123
rect 16715 41089 16724 41123
rect 16672 41080 16724 41089
rect 17500 41080 17552 41132
rect 18328 41148 18380 41200
rect 19616 41148 19668 41200
rect 19708 41148 19760 41200
rect 21916 41216 21968 41268
rect 22008 41216 22060 41268
rect 22468 41216 22520 41268
rect 22284 41148 22336 41200
rect 23112 41216 23164 41268
rect 25412 41216 25464 41268
rect 25780 41259 25832 41268
rect 25780 41225 25789 41259
rect 25789 41225 25823 41259
rect 25823 41225 25832 41259
rect 25780 41216 25832 41225
rect 26240 41216 26292 41268
rect 27712 41259 27764 41268
rect 27712 41225 27721 41259
rect 27721 41225 27755 41259
rect 27755 41225 27764 41259
rect 27712 41216 27764 41225
rect 27896 41216 27948 41268
rect 28080 41216 28132 41268
rect 19340 41080 19392 41132
rect 21364 41080 21416 41132
rect 21640 41080 21692 41132
rect 22468 41123 22520 41132
rect 22468 41089 22477 41123
rect 22477 41089 22511 41123
rect 22511 41089 22520 41123
rect 22468 41080 22520 41089
rect 22744 41080 22796 41132
rect 23204 41080 23256 41132
rect 23388 41080 23440 41132
rect 20168 41012 20220 41064
rect 20444 41055 20496 41064
rect 20444 41021 20453 41055
rect 20453 41021 20487 41055
rect 20487 41021 20496 41055
rect 20444 41012 20496 41021
rect 17500 40944 17552 40996
rect 18696 40944 18748 40996
rect 19892 40987 19944 40996
rect 8208 40876 8260 40928
rect 17040 40876 17092 40928
rect 17592 40876 17644 40928
rect 19892 40953 19901 40987
rect 19901 40953 19935 40987
rect 19935 40953 19944 40987
rect 19892 40944 19944 40953
rect 21180 40944 21232 40996
rect 21732 40944 21784 40996
rect 22008 40944 22060 40996
rect 21272 40876 21324 40928
rect 21548 40876 21600 40928
rect 23572 40944 23624 40996
rect 24768 41012 24820 41064
rect 27620 41080 27672 41132
rect 28172 41148 28224 41200
rect 28264 41148 28316 41200
rect 28724 41216 28776 41268
rect 28908 41216 28960 41268
rect 26424 41012 26476 41064
rect 24676 40944 24728 40996
rect 25136 40944 25188 40996
rect 27436 40944 27488 40996
rect 22928 40876 22980 40928
rect 23296 40876 23348 40928
rect 27528 40876 27580 40928
rect 28172 40876 28224 40928
rect 28816 40876 28868 40928
rect 31852 41216 31904 41268
rect 29920 41123 29972 41132
rect 29920 41089 29934 41123
rect 29934 41089 29968 41123
rect 29968 41089 29972 41123
rect 30104 41123 30156 41132
rect 29920 41080 29972 41089
rect 30104 41089 30113 41123
rect 30113 41089 30147 41123
rect 30147 41089 30156 41123
rect 30104 41080 30156 41089
rect 29828 40876 29880 40928
rect 5915 40774 5967 40826
rect 5979 40774 6031 40826
rect 6043 40774 6095 40826
rect 6107 40774 6159 40826
rect 6171 40774 6223 40826
rect 15846 40774 15898 40826
rect 15910 40774 15962 40826
rect 15974 40774 16026 40826
rect 16038 40774 16090 40826
rect 16102 40774 16154 40826
rect 25776 40774 25828 40826
rect 25840 40774 25892 40826
rect 25904 40774 25956 40826
rect 25968 40774 26020 40826
rect 26032 40774 26084 40826
rect 8668 40672 8720 40724
rect 10140 40672 10192 40724
rect 17408 40672 17460 40724
rect 17868 40715 17920 40724
rect 17868 40681 17877 40715
rect 17877 40681 17911 40715
rect 17911 40681 17920 40715
rect 17868 40672 17920 40681
rect 19340 40715 19392 40724
rect 19340 40681 19349 40715
rect 19349 40681 19383 40715
rect 19383 40681 19392 40715
rect 19340 40672 19392 40681
rect 23480 40672 23532 40724
rect 9864 40604 9916 40656
rect 8392 40536 8444 40588
rect 8208 40511 8260 40520
rect 8208 40477 8217 40511
rect 8217 40477 8251 40511
rect 8251 40477 8260 40511
rect 8208 40468 8260 40477
rect 16948 40604 17000 40656
rect 17316 40604 17368 40656
rect 10140 40536 10192 40588
rect 10048 40511 10100 40520
rect 10048 40477 10057 40511
rect 10057 40477 10091 40511
rect 10091 40477 10100 40511
rect 10324 40536 10376 40588
rect 11244 40536 11296 40588
rect 19892 40536 19944 40588
rect 10048 40468 10100 40477
rect 15752 40511 15804 40520
rect 15752 40477 15761 40511
rect 15761 40477 15795 40511
rect 15795 40477 15804 40511
rect 15752 40468 15804 40477
rect 16948 40468 17000 40520
rect 18052 40468 18104 40520
rect 9680 40332 9732 40384
rect 11336 40400 11388 40452
rect 10140 40332 10192 40384
rect 14004 40332 14056 40384
rect 16856 40332 16908 40384
rect 17960 40332 18012 40384
rect 22468 40604 22520 40656
rect 27804 40604 27856 40656
rect 23480 40536 23532 40588
rect 25780 40536 25832 40588
rect 22100 40468 22152 40520
rect 22284 40468 22336 40520
rect 22468 40468 22520 40520
rect 23572 40511 23624 40520
rect 23572 40477 23581 40511
rect 23581 40477 23615 40511
rect 23615 40477 23624 40511
rect 23572 40468 23624 40477
rect 24308 40468 24360 40520
rect 25872 40443 25924 40452
rect 19616 40332 19668 40384
rect 25872 40409 25881 40443
rect 25881 40409 25915 40443
rect 25915 40409 25924 40443
rect 25872 40400 25924 40409
rect 26056 40443 26108 40452
rect 26056 40409 26065 40443
rect 26065 40409 26099 40443
rect 26099 40409 26108 40443
rect 26056 40400 26108 40409
rect 26332 40332 26384 40384
rect 27528 40511 27580 40520
rect 27528 40477 27549 40511
rect 27549 40477 27580 40511
rect 27528 40468 27580 40477
rect 27436 40332 27488 40384
rect 28356 40536 28408 40588
rect 29920 40511 29972 40520
rect 29920 40477 29929 40511
rect 29929 40477 29963 40511
rect 29963 40477 29972 40511
rect 29920 40468 29972 40477
rect 28356 40400 28408 40452
rect 29000 40400 29052 40452
rect 10880 40230 10932 40282
rect 10944 40230 10996 40282
rect 11008 40230 11060 40282
rect 11072 40230 11124 40282
rect 11136 40230 11188 40282
rect 20811 40230 20863 40282
rect 20875 40230 20927 40282
rect 20939 40230 20991 40282
rect 21003 40230 21055 40282
rect 21067 40230 21119 40282
rect 8668 40171 8720 40180
rect 8668 40137 8677 40171
rect 8677 40137 8711 40171
rect 8711 40137 8720 40171
rect 8668 40128 8720 40137
rect 10324 40128 10376 40180
rect 19984 40171 20036 40180
rect 19984 40137 19993 40171
rect 19993 40137 20027 40171
rect 20027 40137 20036 40171
rect 19984 40128 20036 40137
rect 22744 40171 22796 40180
rect 1584 40035 1636 40044
rect 1584 40001 1593 40035
rect 1593 40001 1627 40035
rect 1627 40001 1636 40035
rect 1584 39992 1636 40001
rect 8392 39992 8444 40044
rect 10140 40060 10192 40112
rect 12900 40060 12952 40112
rect 15752 40060 15804 40112
rect 17040 40103 17092 40112
rect 17040 40069 17049 40103
rect 17049 40069 17083 40103
rect 17083 40069 17092 40103
rect 17040 40060 17092 40069
rect 19708 40060 19760 40112
rect 20444 40060 20496 40112
rect 21456 40060 21508 40112
rect 21180 40035 21232 40044
rect 9864 39856 9916 39908
rect 21180 40001 21189 40035
rect 21189 40001 21223 40035
rect 21223 40001 21232 40035
rect 21180 39992 21232 40001
rect 21640 40060 21692 40112
rect 22744 40137 22753 40171
rect 22753 40137 22787 40171
rect 22787 40137 22796 40171
rect 22744 40128 22796 40137
rect 23204 40171 23256 40180
rect 23204 40137 23213 40171
rect 23213 40137 23247 40171
rect 23247 40137 23256 40171
rect 23204 40128 23256 40137
rect 26056 40128 26108 40180
rect 26240 40128 26292 40180
rect 27528 40128 27580 40180
rect 27620 40171 27672 40180
rect 27620 40137 27629 40171
rect 27629 40137 27663 40171
rect 27663 40137 27672 40171
rect 27620 40128 27672 40137
rect 22652 40060 22704 40112
rect 22468 39992 22520 40044
rect 22744 39992 22796 40044
rect 23572 39992 23624 40044
rect 24308 40035 24360 40044
rect 10140 39924 10192 39976
rect 23296 39924 23348 39976
rect 23480 39924 23532 39976
rect 24308 40001 24317 40035
rect 24317 40001 24351 40035
rect 24351 40001 24360 40035
rect 24308 39992 24360 40001
rect 28172 40060 28224 40112
rect 27436 40035 27488 40044
rect 27436 40001 27445 40035
rect 27445 40001 27479 40035
rect 27479 40001 27488 40035
rect 27436 39992 27488 40001
rect 28540 40060 28592 40112
rect 28816 40060 28868 40112
rect 28356 39992 28408 40044
rect 28172 39967 28224 39976
rect 28172 39933 28181 39967
rect 28181 39933 28215 39967
rect 28215 39933 28224 39967
rect 28172 39924 28224 39933
rect 10600 39856 10652 39908
rect 18236 39856 18288 39908
rect 21456 39856 21508 39908
rect 22100 39856 22152 39908
rect 9956 39788 10008 39840
rect 11520 39788 11572 39840
rect 12164 39788 12216 39840
rect 16580 39788 16632 39840
rect 19616 39788 19668 39840
rect 21824 39788 21876 39840
rect 24768 39856 24820 39908
rect 27620 39856 27672 39908
rect 23480 39788 23532 39840
rect 24584 39788 24636 39840
rect 24676 39788 24728 39840
rect 25136 39788 25188 39840
rect 27528 39788 27580 39840
rect 29920 39856 29972 39908
rect 30196 39856 30248 39908
rect 30012 39831 30064 39840
rect 30012 39797 30021 39831
rect 30021 39797 30055 39831
rect 30055 39797 30064 39831
rect 30012 39788 30064 39797
rect 5915 39686 5967 39738
rect 5979 39686 6031 39738
rect 6043 39686 6095 39738
rect 6107 39686 6159 39738
rect 6171 39686 6223 39738
rect 15846 39686 15898 39738
rect 15910 39686 15962 39738
rect 15974 39686 16026 39738
rect 16038 39686 16090 39738
rect 16102 39686 16154 39738
rect 25776 39686 25828 39738
rect 25840 39686 25892 39738
rect 25904 39686 25956 39738
rect 25968 39686 26020 39738
rect 26032 39686 26084 39738
rect 11888 39584 11940 39636
rect 13912 39584 13964 39636
rect 14280 39627 14332 39636
rect 14280 39593 14289 39627
rect 14289 39593 14323 39627
rect 14323 39593 14332 39627
rect 14280 39584 14332 39593
rect 16948 39584 17000 39636
rect 18696 39627 18748 39636
rect 13544 39516 13596 39568
rect 18696 39593 18705 39627
rect 18705 39593 18739 39627
rect 18739 39593 18748 39627
rect 18696 39584 18748 39593
rect 10600 39491 10652 39500
rect 10600 39457 10609 39491
rect 10609 39457 10643 39491
rect 10643 39457 10652 39491
rect 10600 39448 10652 39457
rect 16580 39491 16632 39500
rect 16580 39457 16589 39491
rect 16589 39457 16623 39491
rect 16623 39457 16632 39491
rect 16580 39448 16632 39457
rect 20720 39448 20772 39500
rect 23204 39584 23256 39636
rect 26608 39584 26660 39636
rect 28264 39584 28316 39636
rect 28908 39584 28960 39636
rect 24492 39516 24544 39568
rect 1584 39423 1636 39432
rect 1584 39389 1593 39423
rect 1593 39389 1627 39423
rect 1627 39389 1636 39423
rect 1584 39380 1636 39389
rect 11428 39380 11480 39432
rect 11612 39423 11664 39432
rect 11612 39389 11621 39423
rect 11621 39389 11655 39423
rect 11655 39389 11664 39423
rect 11612 39380 11664 39389
rect 15016 39380 15068 39432
rect 11704 39312 11756 39364
rect 14188 39355 14240 39364
rect 14188 39321 14197 39355
rect 14197 39321 14231 39355
rect 14231 39321 14240 39355
rect 14188 39312 14240 39321
rect 8576 39244 8628 39296
rect 10048 39244 10100 39296
rect 12164 39244 12216 39296
rect 12716 39244 12768 39296
rect 15384 39312 15436 39364
rect 17408 39312 17460 39364
rect 15660 39244 15712 39296
rect 17224 39244 17276 39296
rect 17592 39423 17644 39432
rect 17592 39389 17626 39423
rect 17626 39389 17644 39423
rect 17592 39380 17644 39389
rect 22928 39380 22980 39432
rect 23296 39423 23348 39432
rect 23296 39389 23305 39423
rect 23305 39389 23339 39423
rect 23339 39389 23348 39423
rect 23296 39380 23348 39389
rect 24584 39423 24636 39432
rect 24584 39389 24593 39423
rect 24593 39389 24627 39423
rect 24627 39389 24636 39423
rect 24584 39380 24636 39389
rect 18696 39312 18748 39364
rect 22652 39312 22704 39364
rect 26240 39380 26292 39432
rect 27988 39423 28040 39432
rect 27988 39389 27997 39423
rect 27997 39389 28031 39423
rect 28031 39389 28040 39423
rect 27988 39380 28040 39389
rect 29460 39380 29512 39432
rect 24768 39312 24820 39364
rect 25872 39312 25924 39364
rect 17868 39244 17920 39296
rect 18420 39244 18472 39296
rect 20168 39244 20220 39296
rect 22284 39287 22336 39296
rect 22284 39253 22293 39287
rect 22293 39253 22327 39287
rect 22327 39253 22336 39287
rect 22284 39244 22336 39253
rect 24676 39244 24728 39296
rect 28172 39287 28224 39296
rect 28172 39253 28181 39287
rect 28181 39253 28215 39287
rect 28215 39253 28224 39287
rect 28172 39244 28224 39253
rect 28908 39287 28960 39296
rect 28908 39253 28917 39287
rect 28917 39253 28951 39287
rect 28951 39253 28960 39287
rect 28908 39244 28960 39253
rect 29184 39244 29236 39296
rect 29644 39244 29696 39296
rect 30104 39244 30156 39296
rect 10880 39142 10932 39194
rect 10944 39142 10996 39194
rect 11008 39142 11060 39194
rect 11072 39142 11124 39194
rect 11136 39142 11188 39194
rect 20811 39142 20863 39194
rect 20875 39142 20927 39194
rect 20939 39142 20991 39194
rect 21003 39142 21055 39194
rect 21067 39142 21119 39194
rect 11704 39040 11756 39092
rect 11888 39040 11940 39092
rect 17224 39083 17276 39092
rect 8392 39015 8444 39024
rect 8392 38981 8401 39015
rect 8401 38981 8435 39015
rect 8435 38981 8444 39015
rect 8392 38972 8444 38981
rect 8576 39015 8628 39024
rect 8576 38981 8585 39015
rect 8585 38981 8619 39015
rect 8619 38981 8628 39015
rect 8576 38972 8628 38981
rect 1584 38947 1636 38956
rect 1584 38913 1593 38947
rect 1593 38913 1627 38947
rect 1627 38913 1636 38947
rect 1584 38904 1636 38913
rect 12532 38972 12584 39024
rect 17224 39049 17233 39083
rect 17233 39049 17267 39083
rect 17267 39049 17276 39083
rect 17224 39040 17276 39049
rect 18512 39040 18564 39092
rect 12164 38947 12216 38956
rect 12164 38913 12173 38947
rect 12173 38913 12207 38947
rect 12207 38913 12216 38947
rect 12164 38904 12216 38913
rect 12992 38904 13044 38956
rect 16580 38972 16632 39024
rect 17868 38972 17920 39024
rect 19524 39015 19576 39024
rect 19524 38981 19533 39015
rect 19533 38981 19567 39015
rect 19567 38981 19576 39015
rect 19524 38972 19576 38981
rect 20812 39015 20864 39024
rect 20812 38981 20821 39015
rect 20821 38981 20855 39015
rect 20855 38981 20864 39015
rect 20812 38972 20864 38981
rect 22652 39040 22704 39092
rect 23572 39040 23624 39092
rect 24768 39040 24820 39092
rect 23020 38972 23072 39024
rect 25964 39040 26016 39092
rect 26056 39040 26108 39092
rect 28356 39040 28408 39092
rect 28632 39040 28684 39092
rect 29000 38972 29052 39024
rect 29736 38972 29788 39024
rect 9036 38768 9088 38820
rect 12164 38768 12216 38820
rect 16304 38904 16356 38956
rect 18420 38904 18472 38956
rect 14096 38879 14148 38888
rect 14096 38845 14105 38879
rect 14105 38845 14139 38879
rect 14139 38845 14148 38879
rect 14096 38836 14148 38845
rect 17408 38836 17460 38888
rect 13452 38768 13504 38820
rect 20076 38904 20128 38956
rect 20168 38904 20220 38956
rect 23572 38836 23624 38888
rect 24584 38904 24636 38956
rect 24952 38904 25004 38956
rect 25228 38904 25280 38956
rect 27528 38904 27580 38956
rect 29828 38947 29880 38956
rect 25872 38836 25924 38888
rect 29828 38913 29837 38947
rect 29837 38913 29871 38947
rect 29871 38913 29880 38947
rect 29828 38904 29880 38913
rect 21088 38768 21140 38820
rect 22928 38768 22980 38820
rect 23664 38768 23716 38820
rect 11796 38700 11848 38752
rect 12992 38700 13044 38752
rect 15568 38700 15620 38752
rect 17408 38700 17460 38752
rect 19340 38700 19392 38752
rect 22744 38700 22796 38752
rect 23848 38700 23900 38752
rect 24952 38768 25004 38820
rect 26056 38768 26108 38820
rect 28632 38700 28684 38752
rect 29368 38700 29420 38752
rect 29920 38700 29972 38752
rect 5915 38598 5967 38650
rect 5979 38598 6031 38650
rect 6043 38598 6095 38650
rect 6107 38598 6159 38650
rect 6171 38598 6223 38650
rect 15846 38598 15898 38650
rect 15910 38598 15962 38650
rect 15974 38598 16026 38650
rect 16038 38598 16090 38650
rect 16102 38598 16154 38650
rect 25776 38598 25828 38650
rect 25840 38598 25892 38650
rect 25904 38598 25956 38650
rect 25968 38598 26020 38650
rect 26032 38598 26084 38650
rect 11244 38496 11296 38548
rect 17684 38496 17736 38548
rect 18052 38539 18104 38548
rect 18052 38505 18061 38539
rect 18061 38505 18095 38539
rect 18095 38505 18104 38539
rect 18052 38496 18104 38505
rect 20812 38496 20864 38548
rect 21088 38539 21140 38548
rect 21088 38505 21097 38539
rect 21097 38505 21131 38539
rect 21131 38505 21140 38539
rect 21088 38496 21140 38505
rect 22928 38496 22980 38548
rect 16488 38428 16540 38480
rect 22192 38428 22244 38480
rect 11428 38360 11480 38412
rect 12624 38360 12676 38412
rect 16212 38360 16264 38412
rect 22928 38360 22980 38412
rect 1584 38335 1636 38344
rect 1584 38301 1593 38335
rect 1593 38301 1627 38335
rect 1627 38301 1636 38335
rect 1584 38292 1636 38301
rect 9772 38292 9824 38344
rect 9956 38335 10008 38344
rect 9956 38301 9990 38335
rect 9990 38301 10008 38335
rect 9956 38292 10008 38301
rect 12164 38292 12216 38344
rect 14096 38335 14148 38344
rect 14096 38301 14105 38335
rect 14105 38301 14139 38335
rect 14139 38301 14148 38335
rect 14096 38292 14148 38301
rect 17960 38335 18012 38344
rect 12992 38224 13044 38276
rect 16672 38224 16724 38276
rect 17960 38301 17969 38335
rect 17969 38301 18003 38335
rect 18003 38301 18012 38335
rect 17960 38292 18012 38301
rect 19340 38292 19392 38344
rect 19984 38292 20036 38344
rect 21548 38292 21600 38344
rect 23572 38428 23624 38480
rect 23664 38428 23716 38480
rect 23388 38360 23440 38412
rect 24032 38360 24084 38412
rect 25228 38496 25280 38548
rect 25504 38496 25556 38548
rect 25228 38360 25280 38412
rect 25872 38360 25924 38412
rect 9864 38156 9916 38208
rect 15476 38199 15528 38208
rect 15476 38165 15485 38199
rect 15485 38165 15519 38199
rect 15519 38165 15528 38199
rect 15476 38156 15528 38165
rect 15660 38156 15712 38208
rect 18880 38156 18932 38208
rect 23848 38156 23900 38208
rect 24124 38156 24176 38208
rect 25780 38292 25832 38344
rect 28908 38496 28960 38548
rect 30380 38496 30432 38548
rect 28172 38428 28224 38480
rect 29828 38428 29880 38480
rect 25504 38224 25556 38276
rect 26608 38292 26660 38344
rect 29184 38292 29236 38344
rect 30196 38292 30248 38344
rect 30380 38292 30432 38344
rect 26056 38224 26108 38276
rect 26240 38224 26292 38276
rect 26608 38156 26660 38208
rect 28264 38199 28316 38208
rect 28264 38165 28273 38199
rect 28273 38165 28307 38199
rect 28307 38165 28316 38199
rect 28264 38156 28316 38165
rect 30196 38156 30248 38208
rect 10880 38054 10932 38106
rect 10944 38054 10996 38106
rect 11008 38054 11060 38106
rect 11072 38054 11124 38106
rect 11136 38054 11188 38106
rect 20811 38054 20863 38106
rect 20875 38054 20927 38106
rect 20939 38054 20991 38106
rect 21003 38054 21055 38106
rect 21067 38054 21119 38106
rect 8392 37952 8444 38004
rect 10048 37952 10100 38004
rect 11612 37952 11664 38004
rect 12716 37952 12768 38004
rect 12992 37995 13044 38004
rect 12992 37961 13001 37995
rect 13001 37961 13035 37995
rect 13035 37961 13044 37995
rect 12992 37952 13044 37961
rect 14188 37952 14240 38004
rect 14556 37952 14608 38004
rect 16672 37995 16724 38004
rect 16672 37961 16681 37995
rect 16681 37961 16715 37995
rect 16715 37961 16724 37995
rect 16672 37952 16724 37961
rect 18512 37952 18564 38004
rect 22652 37952 22704 38004
rect 9036 37927 9088 37936
rect 9036 37893 9045 37927
rect 9045 37893 9079 37927
rect 9079 37893 9088 37927
rect 9036 37884 9088 37893
rect 9864 37927 9916 37936
rect 9864 37893 9873 37927
rect 9873 37893 9907 37927
rect 9907 37893 9916 37927
rect 9864 37884 9916 37893
rect 12164 37884 12216 37936
rect 14004 37927 14056 37936
rect 1400 37816 1452 37868
rect 8300 37859 8352 37868
rect 8300 37825 8309 37859
rect 8309 37825 8343 37859
rect 8343 37825 8352 37859
rect 8300 37816 8352 37825
rect 9588 37816 9640 37868
rect 11428 37816 11480 37868
rect 12440 37816 12492 37868
rect 11612 37791 11664 37800
rect 11612 37757 11621 37791
rect 11621 37757 11655 37791
rect 11655 37757 11664 37791
rect 11612 37748 11664 37757
rect 14004 37893 14013 37927
rect 14013 37893 14047 37927
rect 14047 37893 14056 37927
rect 14004 37884 14056 37893
rect 15476 37884 15528 37936
rect 17316 37859 17368 37868
rect 13728 37680 13780 37732
rect 17316 37825 17325 37859
rect 17325 37825 17359 37859
rect 17359 37825 17368 37859
rect 17316 37816 17368 37825
rect 18236 37884 18288 37936
rect 21732 37884 21784 37936
rect 24584 37884 24636 37936
rect 25228 37952 25280 38004
rect 26056 37995 26108 38004
rect 26056 37961 26065 37995
rect 26065 37961 26099 37995
rect 26099 37961 26108 37995
rect 26056 37952 26108 37961
rect 27252 37995 27304 38004
rect 27252 37961 27261 37995
rect 27261 37961 27295 37995
rect 27295 37961 27304 37995
rect 27252 37952 27304 37961
rect 27620 37952 27672 38004
rect 28816 37952 28868 38004
rect 29828 37952 29880 38004
rect 24878 37927 24930 37936
rect 24878 37893 24887 37927
rect 24887 37893 24921 37927
rect 24921 37893 24930 37927
rect 25872 37927 25924 37936
rect 24878 37884 24930 37893
rect 25872 37893 25881 37927
rect 25881 37893 25915 37927
rect 25915 37893 25924 37927
rect 25872 37884 25924 37893
rect 26608 37884 26660 37936
rect 17224 37748 17276 37800
rect 19616 37816 19668 37868
rect 23664 37859 23716 37868
rect 23664 37825 23673 37859
rect 23673 37825 23707 37859
rect 23707 37825 23716 37859
rect 23664 37816 23716 37825
rect 24124 37816 24176 37868
rect 25044 37859 25096 37868
rect 24492 37723 24544 37732
rect 24492 37689 24501 37723
rect 24501 37689 24535 37723
rect 24535 37689 24544 37723
rect 24492 37680 24544 37689
rect 25044 37825 25053 37859
rect 25053 37825 25087 37859
rect 25087 37825 25096 37859
rect 25044 37816 25096 37825
rect 26976 37816 27028 37868
rect 28172 37884 28224 37936
rect 28264 37859 28316 37868
rect 25228 37748 25280 37800
rect 26240 37748 26292 37800
rect 28264 37825 28273 37859
rect 28273 37825 28307 37859
rect 28307 37825 28316 37859
rect 28264 37816 28316 37825
rect 29460 37816 29512 37868
rect 29828 37816 29880 37868
rect 9128 37612 9180 37664
rect 12256 37612 12308 37664
rect 15660 37612 15712 37664
rect 16212 37612 16264 37664
rect 18328 37612 18380 37664
rect 20168 37655 20220 37664
rect 20168 37621 20177 37655
rect 20177 37621 20211 37655
rect 20211 37621 20220 37655
rect 20168 37612 20220 37621
rect 24768 37612 24820 37664
rect 25044 37612 25096 37664
rect 28356 37612 28408 37664
rect 28724 37612 28776 37664
rect 29000 37612 29052 37664
rect 5915 37510 5967 37562
rect 5979 37510 6031 37562
rect 6043 37510 6095 37562
rect 6107 37510 6159 37562
rect 6171 37510 6223 37562
rect 15846 37510 15898 37562
rect 15910 37510 15962 37562
rect 15974 37510 16026 37562
rect 16038 37510 16090 37562
rect 16102 37510 16154 37562
rect 25776 37510 25828 37562
rect 25840 37510 25892 37562
rect 25904 37510 25956 37562
rect 25968 37510 26020 37562
rect 26032 37510 26084 37562
rect 2504 37408 2556 37460
rect 9588 37451 9640 37460
rect 9588 37417 9597 37451
rect 9597 37417 9631 37451
rect 9631 37417 9640 37451
rect 9588 37408 9640 37417
rect 8208 37204 8260 37256
rect 12164 37408 12216 37460
rect 12440 37451 12492 37460
rect 12440 37417 12449 37451
rect 12449 37417 12483 37451
rect 12483 37417 12492 37451
rect 12440 37408 12492 37417
rect 13544 37408 13596 37460
rect 17224 37451 17276 37460
rect 11796 37340 11848 37392
rect 12532 37340 12584 37392
rect 17224 37417 17233 37451
rect 17233 37417 17267 37451
rect 17267 37417 17276 37451
rect 17224 37408 17276 37417
rect 27160 37408 27212 37460
rect 27252 37408 27304 37460
rect 27528 37408 27580 37460
rect 29184 37408 29236 37460
rect 29552 37408 29604 37460
rect 17684 37340 17736 37392
rect 8300 37136 8352 37188
rect 12532 37204 12584 37256
rect 12716 37247 12768 37256
rect 12716 37213 12725 37247
rect 12725 37213 12759 37247
rect 12759 37213 12768 37247
rect 12716 37204 12768 37213
rect 13728 37272 13780 37324
rect 18236 37315 18288 37324
rect 18236 37281 18245 37315
rect 18245 37281 18279 37315
rect 18279 37281 18288 37315
rect 18236 37272 18288 37281
rect 21916 37340 21968 37392
rect 18972 37272 19024 37324
rect 11704 37068 11756 37120
rect 12256 37136 12308 37188
rect 15200 37204 15252 37256
rect 15016 37136 15068 37188
rect 12808 37068 12860 37120
rect 13544 37068 13596 37120
rect 16672 37204 16724 37256
rect 18420 37247 18472 37256
rect 18420 37213 18429 37247
rect 18429 37213 18463 37247
rect 18463 37213 18472 37247
rect 18420 37204 18472 37213
rect 19248 37247 19300 37256
rect 15568 37136 15620 37188
rect 19248 37213 19257 37247
rect 19257 37213 19291 37247
rect 19291 37213 19300 37247
rect 19248 37204 19300 37213
rect 16488 37111 16540 37120
rect 16488 37077 16497 37111
rect 16497 37077 16531 37111
rect 16531 37077 16540 37111
rect 16488 37068 16540 37077
rect 19892 37136 19944 37188
rect 21272 37247 21324 37256
rect 21272 37213 21281 37247
rect 21281 37213 21315 37247
rect 21315 37213 21324 37247
rect 21272 37204 21324 37213
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 22284 37204 22336 37256
rect 24584 37315 24636 37324
rect 24584 37281 24593 37315
rect 24593 37281 24627 37315
rect 24627 37281 24636 37315
rect 24584 37272 24636 37281
rect 24768 37340 24820 37392
rect 25504 37272 25556 37324
rect 26976 37340 27028 37392
rect 28632 37340 28684 37392
rect 21732 37136 21784 37188
rect 27620 37247 27672 37256
rect 27620 37213 27629 37247
rect 27629 37213 27663 37247
rect 27663 37213 27672 37247
rect 27620 37204 27672 37213
rect 29552 37272 29604 37324
rect 29828 37272 29880 37324
rect 27988 37204 28040 37256
rect 28632 37247 28684 37256
rect 28632 37213 28641 37247
rect 28641 37213 28675 37247
rect 28675 37213 28684 37247
rect 28632 37204 28684 37213
rect 28172 37136 28224 37188
rect 21824 37068 21876 37120
rect 22008 37068 22060 37120
rect 24584 37068 24636 37120
rect 26056 37068 26108 37120
rect 27528 37068 27580 37120
rect 28264 37068 28316 37120
rect 29092 37204 29144 37256
rect 29460 37204 29512 37256
rect 30104 37136 30156 37188
rect 29460 37068 29512 37120
rect 10880 36966 10932 37018
rect 10944 36966 10996 37018
rect 11008 36966 11060 37018
rect 11072 36966 11124 37018
rect 11136 36966 11188 37018
rect 20811 36966 20863 37018
rect 20875 36966 20927 37018
rect 20939 36966 20991 37018
rect 21003 36966 21055 37018
rect 21067 36966 21119 37018
rect 13452 36864 13504 36916
rect 15016 36907 15068 36916
rect 15016 36873 15025 36907
rect 15025 36873 15059 36907
rect 15059 36873 15068 36907
rect 15016 36864 15068 36873
rect 9128 36839 9180 36848
rect 9128 36805 9137 36839
rect 9137 36805 9171 36839
rect 9171 36805 9180 36839
rect 9128 36796 9180 36805
rect 1584 36771 1636 36780
rect 1584 36737 1593 36771
rect 1593 36737 1627 36771
rect 1627 36737 1636 36771
rect 1584 36728 1636 36737
rect 8852 36728 8904 36780
rect 9588 36728 9640 36780
rect 13544 36728 13596 36780
rect 13728 36771 13780 36780
rect 13728 36737 13737 36771
rect 13737 36737 13771 36771
rect 13771 36737 13780 36771
rect 13728 36728 13780 36737
rect 16488 36864 16540 36916
rect 23020 36864 23072 36916
rect 26424 36864 26476 36916
rect 28264 36864 28316 36916
rect 15936 36796 15988 36848
rect 16580 36796 16632 36848
rect 22928 36796 22980 36848
rect 15476 36774 15528 36780
rect 15476 36740 15485 36774
rect 15485 36740 15519 36774
rect 15519 36740 15528 36774
rect 15476 36728 15528 36740
rect 15844 36728 15896 36780
rect 17224 36728 17276 36780
rect 18972 36771 19024 36780
rect 18972 36737 18981 36771
rect 18981 36737 19015 36771
rect 19015 36737 19024 36771
rect 18972 36728 19024 36737
rect 21180 36728 21232 36780
rect 22008 36728 22060 36780
rect 22100 36771 22152 36780
rect 22100 36737 22109 36771
rect 22109 36737 22143 36771
rect 22143 36737 22152 36771
rect 22100 36728 22152 36737
rect 16304 36660 16356 36712
rect 21732 36660 21784 36712
rect 21916 36660 21968 36712
rect 22652 36660 22704 36712
rect 17316 36592 17368 36644
rect 18420 36592 18472 36644
rect 19892 36592 19944 36644
rect 25136 36728 25188 36780
rect 26424 36728 26476 36780
rect 27620 36771 27672 36780
rect 27620 36737 27629 36771
rect 27629 36737 27663 36771
rect 27663 36737 27672 36771
rect 27620 36728 27672 36737
rect 27988 36728 28040 36780
rect 28632 36771 28684 36780
rect 28632 36737 28641 36771
rect 28641 36737 28675 36771
rect 28675 36737 28684 36771
rect 28632 36728 28684 36737
rect 29184 36796 29236 36848
rect 29000 36771 29052 36780
rect 29000 36737 29009 36771
rect 29009 36737 29043 36771
rect 29043 36737 29052 36771
rect 29000 36728 29052 36737
rect 29092 36728 29144 36780
rect 29828 36771 29880 36780
rect 29828 36737 29837 36771
rect 29837 36737 29871 36771
rect 29871 36737 29880 36771
rect 29828 36728 29880 36737
rect 30104 36771 30156 36780
rect 24768 36660 24820 36712
rect 25780 36660 25832 36712
rect 26148 36703 26200 36712
rect 26148 36669 26157 36703
rect 26157 36669 26191 36703
rect 26191 36669 26200 36703
rect 26148 36660 26200 36669
rect 28356 36660 28408 36712
rect 14924 36524 14976 36576
rect 16580 36524 16632 36576
rect 19340 36524 19392 36576
rect 19800 36524 19852 36576
rect 20076 36524 20128 36576
rect 21824 36524 21876 36576
rect 26056 36592 26108 36644
rect 26884 36592 26936 36644
rect 29000 36592 29052 36644
rect 30104 36737 30113 36771
rect 30113 36737 30147 36771
rect 30147 36737 30156 36771
rect 30104 36728 30156 36737
rect 30104 36592 30156 36644
rect 31300 36592 31352 36644
rect 22560 36524 22612 36576
rect 23388 36524 23440 36576
rect 25228 36524 25280 36576
rect 25596 36524 25648 36576
rect 27620 36524 27672 36576
rect 28724 36524 28776 36576
rect 5915 36422 5967 36474
rect 5979 36422 6031 36474
rect 6043 36422 6095 36474
rect 6107 36422 6159 36474
rect 6171 36422 6223 36474
rect 15846 36422 15898 36474
rect 15910 36422 15962 36474
rect 15974 36422 16026 36474
rect 16038 36422 16090 36474
rect 16102 36422 16154 36474
rect 25776 36422 25828 36474
rect 25840 36422 25892 36474
rect 25904 36422 25956 36474
rect 25968 36422 26020 36474
rect 26032 36422 26084 36474
rect 8208 36363 8260 36372
rect 8208 36329 8217 36363
rect 8217 36329 8251 36363
rect 8251 36329 8260 36363
rect 8208 36320 8260 36329
rect 11336 36320 11388 36372
rect 15200 36363 15252 36372
rect 9036 36252 9088 36304
rect 9680 36252 9732 36304
rect 15200 36329 15209 36363
rect 15209 36329 15243 36363
rect 15243 36329 15252 36363
rect 15200 36320 15252 36329
rect 15752 36320 15804 36372
rect 19248 36320 19300 36372
rect 26884 36320 26936 36372
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 8300 36116 8352 36168
rect 9680 36159 9732 36168
rect 9680 36125 9689 36159
rect 9689 36125 9723 36159
rect 9723 36125 9732 36159
rect 9680 36116 9732 36125
rect 20352 36184 20404 36236
rect 20628 36184 20680 36236
rect 15016 36159 15068 36168
rect 15016 36125 15025 36159
rect 15025 36125 15059 36159
rect 15059 36125 15068 36159
rect 15016 36116 15068 36125
rect 16856 36116 16908 36168
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 21456 36227 21508 36236
rect 21456 36193 21465 36227
rect 21465 36193 21499 36227
rect 21499 36193 21508 36227
rect 21456 36184 21508 36193
rect 21180 36159 21232 36168
rect 21180 36125 21189 36159
rect 21189 36125 21223 36159
rect 21223 36125 21232 36159
rect 21180 36116 21232 36125
rect 22100 36116 22152 36168
rect 23664 36252 23716 36304
rect 24768 36252 24820 36304
rect 25964 36252 26016 36304
rect 26516 36252 26568 36304
rect 29920 36252 29972 36304
rect 30564 36252 30616 36304
rect 31392 36252 31444 36304
rect 24032 36184 24084 36236
rect 28172 36184 28224 36236
rect 29368 36184 29420 36236
rect 29552 36184 29604 36236
rect 24768 36116 24820 36168
rect 24952 36159 25004 36168
rect 24952 36125 24961 36159
rect 24961 36125 24995 36159
rect 24995 36125 25004 36159
rect 24952 36116 25004 36125
rect 25136 36116 25188 36168
rect 25780 36116 25832 36168
rect 26884 36116 26936 36168
rect 27436 36116 27488 36168
rect 28356 36159 28408 36168
rect 10048 36048 10100 36100
rect 11980 36048 12032 36100
rect 21824 36048 21876 36100
rect 22284 36048 22336 36100
rect 22560 36048 22612 36100
rect 22928 36048 22980 36100
rect 25872 36091 25924 36100
rect 20352 36023 20404 36032
rect 20352 35989 20361 36023
rect 20361 35989 20395 36023
rect 20395 35989 20404 36023
rect 20352 35980 20404 35989
rect 21916 35980 21968 36032
rect 25872 36057 25881 36091
rect 25881 36057 25915 36091
rect 25915 36057 25924 36091
rect 25872 36048 25924 36057
rect 26240 36048 26292 36100
rect 28356 36125 28365 36159
rect 28365 36125 28399 36159
rect 28399 36125 28408 36159
rect 28356 36116 28408 36125
rect 29920 36159 29972 36168
rect 29920 36125 29929 36159
rect 29929 36125 29963 36159
rect 29963 36125 29972 36159
rect 29920 36116 29972 36125
rect 28264 36048 28316 36100
rect 26056 36023 26108 36032
rect 26056 35989 26065 36023
rect 26065 35989 26099 36023
rect 26099 35989 26108 36023
rect 26056 35980 26108 35989
rect 27436 35980 27488 36032
rect 28356 35980 28408 36032
rect 28632 35980 28684 36032
rect 29184 35980 29236 36032
rect 29368 35980 29420 36032
rect 29552 36023 29604 36032
rect 29552 35989 29561 36023
rect 29561 35989 29595 36023
rect 29595 35989 29604 36023
rect 29552 35980 29604 35989
rect 10880 35878 10932 35930
rect 10944 35878 10996 35930
rect 11008 35878 11060 35930
rect 11072 35878 11124 35930
rect 11136 35878 11188 35930
rect 20811 35878 20863 35930
rect 20875 35878 20927 35930
rect 20939 35878 20991 35930
rect 21003 35878 21055 35930
rect 21067 35878 21119 35930
rect 20536 35776 20588 35828
rect 23664 35776 23716 35828
rect 24032 35776 24084 35828
rect 24768 35776 24820 35828
rect 25964 35776 26016 35828
rect 27988 35776 28040 35828
rect 30288 35776 30340 35828
rect 30840 35776 30892 35828
rect 8852 35751 8904 35760
rect 8852 35717 8861 35751
rect 8861 35717 8895 35751
rect 8895 35717 8904 35751
rect 8852 35708 8904 35717
rect 9036 35751 9088 35760
rect 9036 35717 9045 35751
rect 9045 35717 9079 35751
rect 9079 35717 9088 35751
rect 9036 35708 9088 35717
rect 16672 35708 16724 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 19524 35640 19576 35692
rect 20352 35640 20404 35692
rect 21272 35640 21324 35692
rect 22376 35683 22428 35692
rect 22376 35649 22385 35683
rect 22385 35649 22419 35683
rect 22419 35649 22428 35683
rect 22376 35640 22428 35649
rect 15476 35572 15528 35624
rect 20812 35615 20864 35624
rect 19708 35504 19760 35556
rect 20812 35581 20821 35615
rect 20821 35581 20855 35615
rect 20855 35581 20864 35615
rect 20812 35572 20864 35581
rect 22100 35572 22152 35624
rect 22284 35572 22336 35624
rect 23204 35640 23256 35692
rect 24768 35683 24820 35692
rect 21364 35504 21416 35556
rect 24768 35649 24777 35683
rect 24777 35649 24811 35683
rect 24811 35649 24820 35683
rect 24768 35640 24820 35649
rect 24308 35615 24360 35624
rect 24308 35581 24317 35615
rect 24317 35581 24351 35615
rect 24351 35581 24360 35615
rect 24308 35572 24360 35581
rect 27620 35640 27672 35692
rect 28816 35708 28868 35760
rect 28264 35640 28316 35692
rect 29920 35640 29972 35692
rect 28816 35615 28868 35624
rect 28816 35581 28825 35615
rect 28825 35581 28859 35615
rect 28859 35581 28868 35615
rect 28816 35572 28868 35581
rect 29092 35615 29144 35624
rect 29092 35581 29101 35615
rect 29101 35581 29135 35615
rect 29135 35581 29144 35615
rect 29092 35572 29144 35581
rect 30288 35572 30340 35624
rect 3976 35436 4028 35488
rect 13360 35436 13412 35488
rect 19800 35436 19852 35488
rect 26332 35436 26384 35488
rect 26516 35436 26568 35488
rect 27620 35436 27672 35488
rect 5915 35334 5967 35386
rect 5979 35334 6031 35386
rect 6043 35334 6095 35386
rect 6107 35334 6159 35386
rect 6171 35334 6223 35386
rect 15846 35334 15898 35386
rect 15910 35334 15962 35386
rect 15974 35334 16026 35386
rect 16038 35334 16090 35386
rect 16102 35334 16154 35386
rect 25776 35334 25828 35386
rect 25840 35334 25892 35386
rect 25904 35334 25956 35386
rect 25968 35334 26020 35386
rect 26032 35334 26084 35386
rect 9680 35232 9732 35284
rect 11612 35232 11664 35284
rect 12348 35275 12400 35284
rect 12348 35241 12357 35275
rect 12357 35241 12391 35275
rect 12391 35241 12400 35275
rect 12348 35232 12400 35241
rect 14096 35232 14148 35284
rect 19248 35232 19300 35284
rect 16396 35164 16448 35216
rect 17316 35096 17368 35148
rect 19708 35232 19760 35284
rect 20812 35275 20864 35284
rect 20812 35241 20821 35275
rect 20821 35241 20855 35275
rect 20855 35241 20864 35275
rect 20812 35232 20864 35241
rect 23112 35232 23164 35284
rect 24124 35232 24176 35284
rect 28816 35232 28868 35284
rect 24768 35164 24820 35216
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 1584 35028 1636 35037
rect 10324 35028 10376 35080
rect 10600 34960 10652 35012
rect 12624 35028 12676 35080
rect 14556 35071 14608 35080
rect 14556 35037 14565 35071
rect 14565 35037 14599 35071
rect 14599 35037 14608 35071
rect 14556 35028 14608 35037
rect 15108 35028 15160 35080
rect 18604 35071 18656 35080
rect 18604 35037 18613 35071
rect 18613 35037 18647 35071
rect 18647 35037 18656 35071
rect 18604 35028 18656 35037
rect 18788 35028 18840 35080
rect 20444 35028 20496 35080
rect 21180 35028 21232 35080
rect 22100 35071 22152 35080
rect 22100 35037 22109 35071
rect 22109 35037 22143 35071
rect 22143 35037 22152 35071
rect 22100 35028 22152 35037
rect 14096 34960 14148 35012
rect 17408 34960 17460 35012
rect 19800 34960 19852 35012
rect 4068 34892 4120 34944
rect 16948 34892 17000 34944
rect 17960 34892 18012 34944
rect 18420 34892 18472 34944
rect 19064 34892 19116 34944
rect 21824 34892 21876 34944
rect 24032 35028 24084 35080
rect 26332 35096 26384 35148
rect 27068 35071 27120 35080
rect 27068 35037 27077 35071
rect 27077 35037 27111 35071
rect 27111 35037 27120 35071
rect 27068 35028 27120 35037
rect 28172 35071 28224 35080
rect 28172 35037 28181 35071
rect 28181 35037 28215 35071
rect 28215 35037 28224 35071
rect 28172 35028 28224 35037
rect 30012 35028 30064 35080
rect 30380 35028 30432 35080
rect 28264 34960 28316 35012
rect 27620 34892 27672 34944
rect 30012 34935 30064 34944
rect 30012 34901 30021 34935
rect 30021 34901 30055 34935
rect 30055 34901 30064 34935
rect 30012 34892 30064 34901
rect 10880 34790 10932 34842
rect 10944 34790 10996 34842
rect 11008 34790 11060 34842
rect 11072 34790 11124 34842
rect 11136 34790 11188 34842
rect 20811 34790 20863 34842
rect 20875 34790 20927 34842
rect 20939 34790 20991 34842
rect 21003 34790 21055 34842
rect 21067 34790 21119 34842
rect 9772 34688 9824 34740
rect 13912 34688 13964 34740
rect 17960 34688 18012 34740
rect 19064 34731 19116 34740
rect 19064 34697 19073 34731
rect 19073 34697 19107 34731
rect 19107 34697 19116 34731
rect 19064 34688 19116 34697
rect 20444 34731 20496 34740
rect 20444 34697 20453 34731
rect 20453 34697 20487 34731
rect 20487 34697 20496 34731
rect 20444 34688 20496 34697
rect 27620 34688 27672 34740
rect 28908 34731 28960 34740
rect 28908 34697 28917 34731
rect 28917 34697 28951 34731
rect 28951 34697 28960 34731
rect 28908 34688 28960 34697
rect 29184 34688 29236 34740
rect 29552 34688 29604 34740
rect 13176 34620 13228 34672
rect 15752 34620 15804 34672
rect 18696 34620 18748 34672
rect 20076 34620 20128 34672
rect 24952 34620 25004 34672
rect 1400 34552 1452 34604
rect 9680 34595 9732 34604
rect 9680 34561 9689 34595
rect 9689 34561 9723 34595
rect 9723 34561 9732 34595
rect 9680 34552 9732 34561
rect 9864 34552 9916 34604
rect 12992 34552 13044 34604
rect 14004 34552 14056 34604
rect 14096 34595 14148 34604
rect 14096 34561 14105 34595
rect 14105 34561 14139 34595
rect 14139 34561 14148 34595
rect 14740 34595 14792 34604
rect 14096 34552 14148 34561
rect 14740 34561 14749 34595
rect 14749 34561 14783 34595
rect 14783 34561 14792 34595
rect 14740 34552 14792 34561
rect 19616 34595 19668 34604
rect 19616 34561 19625 34595
rect 19625 34561 19659 34595
rect 19659 34561 19668 34595
rect 19616 34552 19668 34561
rect 20260 34595 20312 34604
rect 20260 34561 20269 34595
rect 20269 34561 20303 34595
rect 20303 34561 20312 34595
rect 20260 34552 20312 34561
rect 27068 34552 27120 34604
rect 10784 34416 10836 34468
rect 17316 34527 17368 34536
rect 17316 34493 17325 34527
rect 17325 34493 17359 34527
rect 17359 34493 17368 34527
rect 17316 34484 17368 34493
rect 17408 34527 17460 34536
rect 17408 34493 17417 34527
rect 17417 34493 17451 34527
rect 17451 34493 17460 34527
rect 18328 34527 18380 34536
rect 17408 34484 17460 34493
rect 18328 34493 18337 34527
rect 18337 34493 18371 34527
rect 18371 34493 18380 34527
rect 18328 34484 18380 34493
rect 19892 34484 19944 34536
rect 20444 34484 20496 34536
rect 26240 34484 26292 34536
rect 29092 34552 29144 34604
rect 30840 34688 30892 34740
rect 29000 34484 29052 34536
rect 13820 34416 13872 34468
rect 27160 34416 27212 34468
rect 27528 34416 27580 34468
rect 29552 34484 29604 34536
rect 11796 34391 11848 34400
rect 11796 34357 11805 34391
rect 11805 34357 11839 34391
rect 11839 34357 11848 34391
rect 11796 34348 11848 34357
rect 11888 34348 11940 34400
rect 14924 34391 14976 34400
rect 14924 34357 14933 34391
rect 14933 34357 14967 34391
rect 14967 34357 14976 34391
rect 14924 34348 14976 34357
rect 17224 34348 17276 34400
rect 17500 34348 17552 34400
rect 21732 34348 21784 34400
rect 24768 34348 24820 34400
rect 26884 34348 26936 34400
rect 29828 34348 29880 34400
rect 5915 34246 5967 34298
rect 5979 34246 6031 34298
rect 6043 34246 6095 34298
rect 6107 34246 6159 34298
rect 6171 34246 6223 34298
rect 15846 34246 15898 34298
rect 15910 34246 15962 34298
rect 15974 34246 16026 34298
rect 16038 34246 16090 34298
rect 16102 34246 16154 34298
rect 25776 34246 25828 34298
rect 25840 34246 25892 34298
rect 25904 34246 25956 34298
rect 25968 34246 26020 34298
rect 26032 34246 26084 34298
rect 9680 34144 9732 34196
rect 14004 34144 14056 34196
rect 12992 34076 13044 34128
rect 13728 34076 13780 34128
rect 17868 34076 17920 34128
rect 11244 34008 11296 34060
rect 11888 34008 11940 34060
rect 13084 34008 13136 34060
rect 17316 34008 17368 34060
rect 1584 33983 1636 33992
rect 1584 33949 1593 33983
rect 1593 33949 1627 33983
rect 1627 33949 1636 33983
rect 1584 33940 1636 33949
rect 10784 33983 10836 33992
rect 10784 33949 10793 33983
rect 10793 33949 10827 33983
rect 10827 33949 10836 33983
rect 10784 33940 10836 33949
rect 13820 33940 13872 33992
rect 15108 33940 15160 33992
rect 17500 33940 17552 33992
rect 12992 33872 13044 33924
rect 9956 33804 10008 33856
rect 11520 33804 11572 33856
rect 11612 33804 11664 33856
rect 12348 33804 12400 33856
rect 13544 33847 13596 33856
rect 13544 33813 13553 33847
rect 13553 33813 13587 33847
rect 13587 33813 13596 33847
rect 13544 33804 13596 33813
rect 13728 33872 13780 33924
rect 18052 33915 18104 33924
rect 18052 33881 18061 33915
rect 18061 33881 18095 33915
rect 18095 33881 18104 33915
rect 18052 33872 18104 33881
rect 19616 34144 19668 34196
rect 25044 34144 25096 34196
rect 19524 34076 19576 34128
rect 19892 34076 19944 34128
rect 25596 34076 25648 34128
rect 25964 34076 26016 34128
rect 26700 34144 26752 34196
rect 28172 34187 28224 34196
rect 28172 34153 28181 34187
rect 28181 34153 28215 34187
rect 28215 34153 28224 34187
rect 28172 34144 28224 34153
rect 24860 34008 24912 34060
rect 19984 33983 20036 33992
rect 19984 33949 19993 33983
rect 19993 33949 20027 33983
rect 20027 33949 20036 33983
rect 19984 33940 20036 33949
rect 23296 33940 23348 33992
rect 25044 33940 25096 33992
rect 26700 34008 26752 34060
rect 25780 33983 25832 33992
rect 25780 33949 25789 33983
rect 25789 33949 25823 33983
rect 25823 33949 25832 33983
rect 25780 33940 25832 33949
rect 26884 33940 26936 33992
rect 27988 33983 28040 33992
rect 27988 33949 27997 33983
rect 27997 33949 28031 33983
rect 28031 33949 28040 33983
rect 27988 33940 28040 33949
rect 28816 33940 28868 33992
rect 29828 33983 29880 33992
rect 29828 33949 29837 33983
rect 29837 33949 29871 33983
rect 29871 33949 29880 33983
rect 29828 33940 29880 33949
rect 17408 33804 17460 33856
rect 25688 33872 25740 33924
rect 27252 33872 27304 33924
rect 19432 33847 19484 33856
rect 19432 33813 19441 33847
rect 19441 33813 19475 33847
rect 19475 33813 19484 33847
rect 19432 33804 19484 33813
rect 28908 33847 28960 33856
rect 28908 33813 28917 33847
rect 28917 33813 28951 33847
rect 28951 33813 28960 33847
rect 28908 33804 28960 33813
rect 29368 33804 29420 33856
rect 29828 33804 29880 33856
rect 30012 33847 30064 33856
rect 30012 33813 30021 33847
rect 30021 33813 30055 33847
rect 30055 33813 30064 33847
rect 30012 33804 30064 33813
rect 10880 33702 10932 33754
rect 10944 33702 10996 33754
rect 11008 33702 11060 33754
rect 11072 33702 11124 33754
rect 11136 33702 11188 33754
rect 20811 33702 20863 33754
rect 20875 33702 20927 33754
rect 20939 33702 20991 33754
rect 21003 33702 21055 33754
rect 21067 33702 21119 33754
rect 12072 33600 12124 33652
rect 13728 33600 13780 33652
rect 11520 33532 11572 33584
rect 13268 33532 13320 33584
rect 17316 33600 17368 33652
rect 24768 33600 24820 33652
rect 26240 33643 26292 33652
rect 1400 33464 1452 33516
rect 11244 33464 11296 33516
rect 11612 33507 11664 33516
rect 11612 33473 11621 33507
rect 11621 33473 11655 33507
rect 11655 33473 11664 33507
rect 11612 33464 11664 33473
rect 12992 33464 13044 33516
rect 16212 33464 16264 33516
rect 16948 33532 17000 33584
rect 19524 33532 19576 33584
rect 19892 33575 19944 33584
rect 19892 33541 19901 33575
rect 19901 33541 19935 33575
rect 19935 33541 19944 33575
rect 19892 33532 19944 33541
rect 25136 33532 25188 33584
rect 17500 33507 17552 33516
rect 10784 33439 10836 33448
rect 10324 33371 10376 33380
rect 10324 33337 10333 33371
rect 10333 33337 10367 33371
rect 10367 33337 10376 33371
rect 10324 33328 10376 33337
rect 10784 33405 10793 33439
rect 10793 33405 10827 33439
rect 10827 33405 10836 33439
rect 10784 33396 10836 33405
rect 13084 33439 13136 33448
rect 13084 33405 13093 33439
rect 13093 33405 13127 33439
rect 13127 33405 13136 33439
rect 13084 33396 13136 33405
rect 15200 33396 15252 33448
rect 17500 33473 17509 33507
rect 17509 33473 17543 33507
rect 17543 33473 17552 33507
rect 17500 33464 17552 33473
rect 19432 33464 19484 33516
rect 24676 33507 24728 33516
rect 24676 33473 24685 33507
rect 24685 33473 24719 33507
rect 24719 33473 24728 33507
rect 24676 33464 24728 33473
rect 24768 33464 24820 33516
rect 25044 33507 25096 33516
rect 25044 33473 25053 33507
rect 25053 33473 25087 33507
rect 25087 33473 25096 33507
rect 26240 33609 26249 33643
rect 26249 33609 26283 33643
rect 26283 33609 26292 33643
rect 26240 33600 26292 33609
rect 25872 33575 25924 33584
rect 25872 33541 25881 33575
rect 25881 33541 25915 33575
rect 25915 33541 25924 33575
rect 25872 33532 25924 33541
rect 26148 33532 26200 33584
rect 25044 33464 25096 33473
rect 17408 33396 17460 33448
rect 18328 33396 18380 33448
rect 26884 33532 26936 33584
rect 27988 33464 28040 33516
rect 25964 33396 26016 33448
rect 27160 33396 27212 33448
rect 28264 33396 28316 33448
rect 11612 33328 11664 33380
rect 12624 33371 12676 33380
rect 12624 33337 12633 33371
rect 12633 33337 12667 33371
rect 12667 33337 12676 33371
rect 12624 33328 12676 33337
rect 14740 33328 14792 33380
rect 15016 33371 15068 33380
rect 15016 33337 15025 33371
rect 15025 33337 15059 33371
rect 15059 33337 15068 33371
rect 15016 33328 15068 33337
rect 24676 33328 24728 33380
rect 25872 33328 25924 33380
rect 9772 33260 9824 33312
rect 20628 33303 20680 33312
rect 20628 33269 20637 33303
rect 20637 33269 20671 33303
rect 20671 33269 20680 33303
rect 20628 33260 20680 33269
rect 26332 33260 26384 33312
rect 29276 33303 29328 33312
rect 29276 33269 29285 33303
rect 29285 33269 29319 33303
rect 29319 33269 29328 33303
rect 29276 33260 29328 33269
rect 30840 33260 30892 33312
rect 5915 33158 5967 33210
rect 5979 33158 6031 33210
rect 6043 33158 6095 33210
rect 6107 33158 6159 33210
rect 6171 33158 6223 33210
rect 15846 33158 15898 33210
rect 15910 33158 15962 33210
rect 15974 33158 16026 33210
rect 16038 33158 16090 33210
rect 16102 33158 16154 33210
rect 25776 33158 25828 33210
rect 25840 33158 25892 33210
rect 25904 33158 25956 33210
rect 25968 33158 26020 33210
rect 26032 33158 26084 33210
rect 10600 33056 10652 33108
rect 11336 33056 11388 33108
rect 14372 33056 14424 33108
rect 16212 33099 16264 33108
rect 11244 32988 11296 33040
rect 16212 33065 16221 33099
rect 16221 33065 16255 33099
rect 16255 33065 16264 33099
rect 16212 33056 16264 33065
rect 18972 33056 19024 33108
rect 20260 33056 20312 33108
rect 1492 32852 1544 32904
rect 9864 32852 9916 32904
rect 16580 32988 16632 33040
rect 22928 33056 22980 33108
rect 20536 32988 20588 33040
rect 25780 32988 25832 33040
rect 17408 32963 17460 32972
rect 17408 32929 17417 32963
rect 17417 32929 17451 32963
rect 17451 32929 17460 32963
rect 19708 32963 19760 32972
rect 17408 32920 17460 32929
rect 19708 32929 19717 32963
rect 19717 32929 19751 32963
rect 19751 32929 19760 32963
rect 19708 32920 19760 32929
rect 11612 32852 11664 32904
rect 13636 32852 13688 32904
rect 14924 32852 14976 32904
rect 17132 32895 17184 32904
rect 17132 32861 17141 32895
rect 17141 32861 17175 32895
rect 17175 32861 17184 32895
rect 17132 32852 17184 32861
rect 19432 32852 19484 32904
rect 20536 32895 20588 32904
rect 20536 32861 20545 32895
rect 20545 32861 20579 32895
rect 20579 32861 20588 32895
rect 20536 32852 20588 32861
rect 21272 32895 21324 32904
rect 21272 32861 21281 32895
rect 21281 32861 21315 32895
rect 21315 32861 21324 32895
rect 21272 32852 21324 32861
rect 21916 32920 21968 32972
rect 22468 32895 22520 32904
rect 22468 32861 22477 32895
rect 22477 32861 22511 32895
rect 22511 32861 22520 32895
rect 22468 32852 22520 32861
rect 29736 32920 29788 32972
rect 22928 32852 22980 32904
rect 23940 32852 23992 32904
rect 25872 32852 25924 32904
rect 26884 32852 26936 32904
rect 28724 32895 28776 32904
rect 28724 32861 28733 32895
rect 28733 32861 28767 32895
rect 28767 32861 28776 32895
rect 28724 32852 28776 32861
rect 9680 32784 9732 32836
rect 2596 32716 2648 32768
rect 11520 32716 11572 32768
rect 14280 32784 14332 32836
rect 14464 32827 14516 32836
rect 14464 32793 14498 32827
rect 14498 32793 14516 32827
rect 14464 32784 14516 32793
rect 17040 32784 17092 32836
rect 19064 32784 19116 32836
rect 24032 32784 24084 32836
rect 24952 32784 25004 32836
rect 14740 32716 14792 32768
rect 18052 32716 18104 32768
rect 20720 32716 20772 32768
rect 22008 32716 22060 32768
rect 23296 32716 23348 32768
rect 25044 32716 25096 32768
rect 29736 32784 29788 32836
rect 30564 32784 30616 32836
rect 25596 32716 25648 32768
rect 27988 32716 28040 32768
rect 28448 32716 28500 32768
rect 28632 32716 28684 32768
rect 28908 32759 28960 32768
rect 28908 32725 28917 32759
rect 28917 32725 28951 32759
rect 28951 32725 28960 32759
rect 28908 32716 28960 32725
rect 30196 32716 30248 32768
rect 10880 32614 10932 32666
rect 10944 32614 10996 32666
rect 11008 32614 11060 32666
rect 11072 32614 11124 32666
rect 11136 32614 11188 32666
rect 20811 32614 20863 32666
rect 20875 32614 20927 32666
rect 20939 32614 20991 32666
rect 21003 32614 21055 32666
rect 21067 32614 21119 32666
rect 10416 32512 10468 32564
rect 13176 32555 13228 32564
rect 13176 32521 13185 32555
rect 13185 32521 13219 32555
rect 13219 32521 13228 32555
rect 13176 32512 13228 32521
rect 14464 32512 14516 32564
rect 18052 32512 18104 32564
rect 18696 32512 18748 32564
rect 19064 32512 19116 32564
rect 20536 32512 20588 32564
rect 23664 32512 23716 32564
rect 9772 32487 9824 32496
rect 9772 32453 9781 32487
rect 9781 32453 9815 32487
rect 9815 32453 9824 32487
rect 9772 32444 9824 32453
rect 11152 32444 11204 32496
rect 11520 32444 11572 32496
rect 11796 32444 11848 32496
rect 13636 32444 13688 32496
rect 17132 32444 17184 32496
rect 17408 32444 17460 32496
rect 1584 32419 1636 32428
rect 1584 32385 1593 32419
rect 1593 32385 1627 32419
rect 1627 32385 1636 32419
rect 1584 32376 1636 32385
rect 9680 32376 9732 32428
rect 14372 32419 14424 32428
rect 14372 32385 14381 32419
rect 14381 32385 14415 32419
rect 14415 32385 14424 32419
rect 14372 32376 14424 32385
rect 14464 32385 14470 32412
rect 14470 32385 14504 32412
rect 14504 32385 14516 32412
rect 14464 32360 14516 32385
rect 14556 32419 14608 32428
rect 14556 32385 14570 32419
rect 14570 32385 14604 32419
rect 14604 32385 14608 32419
rect 14556 32376 14608 32385
rect 14740 32419 14792 32428
rect 14740 32385 14749 32419
rect 14749 32385 14783 32419
rect 14783 32385 14792 32419
rect 14740 32376 14792 32385
rect 15108 32376 15160 32428
rect 18788 32419 18840 32428
rect 18788 32385 18797 32419
rect 18797 32385 18831 32419
rect 18831 32385 18840 32419
rect 18788 32376 18840 32385
rect 20168 32444 20220 32496
rect 22192 32487 22244 32496
rect 22192 32453 22201 32487
rect 22201 32453 22235 32487
rect 22235 32453 22244 32487
rect 22192 32444 22244 32453
rect 22468 32444 22520 32496
rect 19892 32419 19944 32428
rect 19892 32385 19926 32419
rect 19926 32385 19944 32419
rect 19892 32376 19944 32385
rect 21824 32376 21876 32428
rect 22100 32419 22152 32428
rect 22100 32385 22109 32419
rect 22109 32385 22143 32419
rect 22143 32385 22152 32419
rect 22100 32376 22152 32385
rect 22744 32376 22796 32428
rect 18328 32308 18380 32360
rect 18604 32308 18656 32360
rect 11060 32240 11112 32292
rect 11244 32240 11296 32292
rect 22376 32308 22428 32360
rect 22744 32240 22796 32292
rect 23020 32240 23072 32292
rect 2320 32172 2372 32224
rect 12348 32172 12400 32224
rect 15752 32172 15804 32224
rect 16304 32172 16356 32224
rect 18420 32172 18472 32224
rect 24032 32376 24084 32428
rect 26332 32376 26384 32428
rect 25872 32351 25924 32360
rect 25872 32317 25881 32351
rect 25881 32317 25915 32351
rect 25915 32317 25924 32351
rect 25872 32308 25924 32317
rect 28080 32376 28132 32428
rect 28172 32240 28224 32292
rect 28724 32419 28776 32428
rect 28724 32385 28733 32419
rect 28733 32385 28767 32419
rect 28767 32385 28776 32419
rect 28724 32376 28776 32385
rect 29000 32376 29052 32428
rect 29828 32308 29880 32360
rect 29368 32240 29420 32292
rect 26240 32172 26292 32224
rect 27712 32172 27764 32224
rect 5915 32070 5967 32122
rect 5979 32070 6031 32122
rect 6043 32070 6095 32122
rect 6107 32070 6159 32122
rect 6171 32070 6223 32122
rect 15846 32070 15898 32122
rect 15910 32070 15962 32122
rect 15974 32070 16026 32122
rect 16038 32070 16090 32122
rect 16102 32070 16154 32122
rect 25776 32070 25828 32122
rect 25840 32070 25892 32122
rect 25904 32070 25956 32122
rect 25968 32070 26020 32122
rect 26032 32070 26084 32122
rect 9680 31900 9732 31952
rect 11244 31900 11296 31952
rect 11428 31968 11480 32020
rect 13084 31968 13136 32020
rect 14280 32011 14332 32020
rect 14280 31977 14289 32011
rect 14289 31977 14323 32011
rect 14323 31977 14332 32011
rect 14280 31968 14332 31977
rect 15568 31968 15620 32020
rect 19892 31968 19944 32020
rect 22192 31968 22244 32020
rect 11336 31832 11388 31884
rect 12072 31832 12124 31884
rect 1860 31807 1912 31816
rect 1860 31773 1869 31807
rect 1869 31773 1903 31807
rect 1903 31773 1912 31807
rect 1860 31764 1912 31773
rect 2504 31764 2556 31816
rect 2596 31807 2648 31816
rect 2596 31773 2605 31807
rect 2605 31773 2639 31807
rect 2639 31773 2648 31807
rect 2596 31764 2648 31773
rect 9772 31764 9824 31816
rect 10048 31764 10100 31816
rect 11060 31764 11112 31816
rect 13820 31832 13872 31884
rect 11152 31696 11204 31748
rect 15936 31900 15988 31952
rect 18972 31900 19024 31952
rect 21916 31900 21968 31952
rect 22100 31900 22152 31952
rect 22652 31968 22704 32020
rect 23204 31968 23256 32020
rect 23572 31968 23624 32020
rect 24032 31968 24084 32020
rect 24676 31968 24728 32020
rect 26056 31900 26108 31952
rect 28448 31968 28500 32020
rect 30380 31968 30432 32020
rect 28264 31900 28316 31952
rect 29736 31900 29788 31952
rect 18144 31832 18196 31884
rect 18788 31832 18840 31884
rect 19984 31832 20036 31884
rect 22468 31875 22520 31884
rect 22468 31841 22477 31875
rect 22477 31841 22511 31875
rect 22511 31841 22520 31875
rect 22468 31832 22520 31841
rect 24124 31832 24176 31884
rect 14096 31807 14148 31816
rect 14096 31773 14105 31807
rect 14105 31773 14139 31807
rect 14139 31773 14148 31807
rect 14096 31764 14148 31773
rect 16672 31764 16724 31816
rect 17684 31764 17736 31816
rect 18236 31764 18288 31816
rect 20720 31764 20772 31816
rect 21272 31764 21324 31816
rect 21916 31807 21968 31816
rect 15016 31696 15068 31748
rect 1676 31671 1728 31680
rect 1676 31637 1685 31671
rect 1685 31637 1719 31671
rect 1719 31637 1728 31671
rect 1676 31628 1728 31637
rect 12164 31628 12216 31680
rect 12808 31628 12860 31680
rect 15292 31628 15344 31680
rect 15568 31628 15620 31680
rect 15660 31628 15712 31680
rect 16764 31628 16816 31680
rect 18696 31696 18748 31748
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22100 31764 22152 31816
rect 25412 31832 25464 31884
rect 25596 31832 25648 31884
rect 27252 31875 27304 31884
rect 27252 31841 27261 31875
rect 27261 31841 27295 31875
rect 27295 31841 27304 31875
rect 27252 31832 27304 31841
rect 27712 31832 27764 31884
rect 28080 31832 28132 31884
rect 28724 31832 28776 31884
rect 23112 31696 23164 31748
rect 24676 31764 24728 31816
rect 23572 31696 23624 31748
rect 26240 31764 26292 31816
rect 30380 31832 30432 31884
rect 23664 31628 23716 31680
rect 27068 31696 27120 31748
rect 27344 31739 27396 31748
rect 27344 31705 27353 31739
rect 27353 31705 27387 31739
rect 27387 31705 27396 31739
rect 27344 31696 27396 31705
rect 30104 31764 30156 31816
rect 30840 31900 30892 31952
rect 26792 31628 26844 31680
rect 29368 31696 29420 31748
rect 30012 31628 30064 31680
rect 30196 31628 30248 31680
rect 30564 31628 30616 31680
rect 10880 31526 10932 31578
rect 10944 31526 10996 31578
rect 11008 31526 11060 31578
rect 11072 31526 11124 31578
rect 11136 31526 11188 31578
rect 20811 31526 20863 31578
rect 20875 31526 20927 31578
rect 20939 31526 20991 31578
rect 21003 31526 21055 31578
rect 21067 31526 21119 31578
rect 4068 31424 4120 31476
rect 2504 31356 2556 31408
rect 3976 31356 4028 31408
rect 12072 31424 12124 31476
rect 13268 31467 13320 31476
rect 13268 31433 13277 31467
rect 13277 31433 13311 31467
rect 13311 31433 13320 31467
rect 13268 31424 13320 31433
rect 14004 31424 14056 31476
rect 14556 31424 14608 31476
rect 15016 31424 15068 31476
rect 13084 31356 13136 31408
rect 15384 31356 15436 31408
rect 15568 31356 15620 31408
rect 1860 31331 1912 31340
rect 1860 31297 1869 31331
rect 1869 31297 1903 31331
rect 1903 31297 1912 31331
rect 1860 31288 1912 31297
rect 2320 31288 2372 31340
rect 9680 31331 9732 31340
rect 9680 31297 9689 31331
rect 9689 31297 9723 31331
rect 9723 31297 9732 31331
rect 9680 31288 9732 31297
rect 15108 31288 15160 31340
rect 15660 31288 15712 31340
rect 15936 31331 15988 31340
rect 15936 31297 15945 31331
rect 15945 31297 15979 31331
rect 15979 31297 15988 31331
rect 17316 31424 17368 31476
rect 21824 31424 21876 31476
rect 23112 31467 23164 31476
rect 23112 31433 23121 31467
rect 23121 31433 23155 31467
rect 23155 31433 23164 31467
rect 23112 31424 23164 31433
rect 24768 31424 24820 31476
rect 24860 31424 24912 31476
rect 19524 31356 19576 31408
rect 15936 31288 15988 31297
rect 18328 31288 18380 31340
rect 22100 31288 22152 31340
rect 22560 31356 22612 31408
rect 26976 31424 27028 31476
rect 27712 31424 27764 31476
rect 27528 31356 27580 31408
rect 30012 31356 30064 31408
rect 23020 31288 23072 31340
rect 23572 31331 23624 31340
rect 23572 31297 23581 31331
rect 23581 31297 23615 31331
rect 23615 31297 23624 31331
rect 23572 31288 23624 31297
rect 23940 31288 23992 31340
rect 24124 31288 24176 31340
rect 25504 31288 25556 31340
rect 9956 31152 10008 31204
rect 16672 31220 16724 31272
rect 1400 31084 1452 31136
rect 13452 31084 13504 31136
rect 16948 31152 17000 31204
rect 18512 31220 18564 31272
rect 22192 31220 22244 31272
rect 26332 31288 26384 31340
rect 26700 31288 26752 31340
rect 26976 31288 27028 31340
rect 27068 31288 27120 31340
rect 27252 31288 27304 31340
rect 27528 31263 27580 31272
rect 27528 31229 27537 31263
rect 27537 31229 27571 31263
rect 27571 31229 27580 31263
rect 27528 31220 27580 31229
rect 29368 31288 29420 31340
rect 29552 31263 29604 31272
rect 29552 31229 29561 31263
rect 29561 31229 29595 31263
rect 29595 31229 29604 31263
rect 29552 31220 29604 31229
rect 30012 31220 30064 31272
rect 14188 31084 14240 31136
rect 15200 31084 15252 31136
rect 15660 31084 15712 31136
rect 16764 31127 16816 31136
rect 16764 31093 16773 31127
rect 16773 31093 16807 31127
rect 16807 31093 16816 31127
rect 16764 31084 16816 31093
rect 18144 31084 18196 31136
rect 18788 31127 18840 31136
rect 18788 31093 18797 31127
rect 18797 31093 18831 31127
rect 18831 31093 18840 31127
rect 18788 31084 18840 31093
rect 19064 31084 19116 31136
rect 23204 31084 23256 31136
rect 23664 31084 23716 31136
rect 24032 31084 24084 31136
rect 26148 31152 26200 31204
rect 24676 31084 24728 31136
rect 25136 31084 25188 31136
rect 25596 31084 25648 31136
rect 29368 31152 29420 31204
rect 26332 31084 26384 31136
rect 5915 30982 5967 31034
rect 5979 30982 6031 31034
rect 6043 30982 6095 31034
rect 6107 30982 6159 31034
rect 6171 30982 6223 31034
rect 15846 30982 15898 31034
rect 15910 30982 15962 31034
rect 15974 30982 16026 31034
rect 16038 30982 16090 31034
rect 16102 30982 16154 31034
rect 25776 30982 25828 31034
rect 25840 30982 25892 31034
rect 25904 30982 25956 31034
rect 25968 30982 26020 31034
rect 26032 30982 26084 31034
rect 31484 31016 31536 31068
rect 11428 30880 11480 30932
rect 25596 30880 25648 30932
rect 26148 30880 26200 30932
rect 28356 30923 28408 30932
rect 28356 30889 28365 30923
rect 28365 30889 28399 30923
rect 28399 30889 28408 30923
rect 28356 30880 28408 30889
rect 30104 30923 30156 30932
rect 30104 30889 30113 30923
rect 30113 30889 30147 30923
rect 30147 30889 30156 30923
rect 30104 30880 30156 30889
rect 1860 30812 1912 30864
rect 9956 30744 10008 30796
rect 17960 30812 18012 30864
rect 21456 30812 21508 30864
rect 23204 30812 23256 30864
rect 25044 30812 25096 30864
rect 1768 30676 1820 30728
rect 4068 30676 4120 30728
rect 9680 30719 9732 30728
rect 9680 30685 9689 30719
rect 9689 30685 9723 30719
rect 9723 30685 9732 30719
rect 9680 30676 9732 30685
rect 9864 30719 9916 30728
rect 9864 30685 9873 30719
rect 9873 30685 9907 30719
rect 9907 30685 9916 30719
rect 9864 30676 9916 30685
rect 11244 30676 11296 30728
rect 13636 30608 13688 30660
rect 1584 30583 1636 30592
rect 1584 30549 1593 30583
rect 1593 30549 1627 30583
rect 1627 30549 1636 30583
rect 1584 30540 1636 30549
rect 2136 30583 2188 30592
rect 2136 30549 2145 30583
rect 2145 30549 2179 30583
rect 2179 30549 2188 30583
rect 2136 30540 2188 30549
rect 11244 30583 11296 30592
rect 11244 30549 11253 30583
rect 11253 30549 11287 30583
rect 11287 30549 11296 30583
rect 11244 30540 11296 30549
rect 15200 30583 15252 30592
rect 15200 30549 15209 30583
rect 15209 30549 15243 30583
rect 15243 30549 15252 30583
rect 15200 30540 15252 30549
rect 15568 30719 15620 30728
rect 15568 30685 15577 30719
rect 15577 30685 15611 30719
rect 15611 30685 15620 30719
rect 15568 30676 15620 30685
rect 18696 30719 18748 30728
rect 18696 30685 18705 30719
rect 18705 30685 18739 30719
rect 18739 30685 18748 30719
rect 18696 30676 18748 30685
rect 18972 30744 19024 30796
rect 19064 30676 19116 30728
rect 19616 30676 19668 30728
rect 22560 30744 22612 30796
rect 23940 30676 23992 30728
rect 25136 30744 25188 30796
rect 25596 30744 25648 30796
rect 28264 30744 28316 30796
rect 24952 30676 25004 30728
rect 25412 30676 25464 30728
rect 26148 30676 26200 30728
rect 27068 30676 27120 30728
rect 28632 30719 28684 30728
rect 28632 30685 28641 30719
rect 28641 30685 28675 30719
rect 28675 30685 28684 30719
rect 28632 30676 28684 30685
rect 16212 30608 16264 30660
rect 20628 30608 20680 30660
rect 20720 30608 20772 30660
rect 26332 30608 26384 30660
rect 15476 30540 15528 30592
rect 17592 30583 17644 30592
rect 17592 30549 17601 30583
rect 17601 30549 17635 30583
rect 17635 30549 17644 30583
rect 17592 30540 17644 30549
rect 18512 30583 18564 30592
rect 18512 30549 18521 30583
rect 18521 30549 18555 30583
rect 18555 30549 18564 30583
rect 18512 30540 18564 30549
rect 19524 30583 19576 30592
rect 19524 30549 19533 30583
rect 19533 30549 19567 30583
rect 19567 30549 19576 30583
rect 19524 30540 19576 30549
rect 28724 30540 28776 30592
rect 29092 30676 29144 30728
rect 29368 30676 29420 30728
rect 29092 30540 29144 30592
rect 29552 30608 29604 30660
rect 30380 30608 30432 30660
rect 31760 30608 31812 30660
rect 10880 30438 10932 30490
rect 10944 30438 10996 30490
rect 11008 30438 11060 30490
rect 11072 30438 11124 30490
rect 11136 30438 11188 30490
rect 20811 30438 20863 30490
rect 20875 30438 20927 30490
rect 20939 30438 20991 30490
rect 21003 30438 21055 30490
rect 21067 30438 21119 30490
rect 12808 30336 12860 30388
rect 13452 30336 13504 30388
rect 14740 30336 14792 30388
rect 18696 30336 18748 30388
rect 19892 30336 19944 30388
rect 11612 30268 11664 30320
rect 13728 30268 13780 30320
rect 1676 30200 1728 30252
rect 11244 30200 11296 30252
rect 14464 30268 14516 30320
rect 11428 30132 11480 30184
rect 13084 30132 13136 30184
rect 14004 30243 14056 30252
rect 14004 30209 14013 30243
rect 14013 30209 14047 30243
rect 14047 30209 14056 30243
rect 14004 30200 14056 30209
rect 14188 30243 14240 30252
rect 14188 30209 14197 30243
rect 14197 30209 14231 30243
rect 14231 30209 14240 30243
rect 17960 30268 18012 30320
rect 19432 30311 19484 30320
rect 19432 30277 19441 30311
rect 19441 30277 19475 30311
rect 19475 30277 19484 30311
rect 19432 30268 19484 30277
rect 19800 30268 19852 30320
rect 14188 30200 14240 30209
rect 18696 30200 18748 30252
rect 19064 30200 19116 30252
rect 27712 30336 27764 30388
rect 28080 30336 28132 30388
rect 28356 30336 28408 30388
rect 26148 30268 26200 30320
rect 26332 30268 26384 30320
rect 27620 30268 27672 30320
rect 30012 30336 30064 30388
rect 25412 30200 25464 30252
rect 27804 30200 27856 30252
rect 14648 30132 14700 30184
rect 25596 30175 25648 30184
rect 25596 30141 25605 30175
rect 25605 30141 25639 30175
rect 25639 30141 25648 30175
rect 25596 30132 25648 30141
rect 29368 30200 29420 30252
rect 1584 30039 1636 30048
rect 1584 30005 1593 30039
rect 1593 30005 1627 30039
rect 1627 30005 1636 30039
rect 1584 29996 1636 30005
rect 1676 29996 1728 30048
rect 14004 29996 14056 30048
rect 17776 29996 17828 30048
rect 18972 30039 19024 30048
rect 18972 30005 18981 30039
rect 18981 30005 19015 30039
rect 19015 30005 19024 30039
rect 18972 29996 19024 30005
rect 25136 30064 25188 30116
rect 28908 30132 28960 30184
rect 29552 30175 29604 30184
rect 29552 30141 29561 30175
rect 29561 30141 29595 30175
rect 29595 30141 29604 30175
rect 29552 30132 29604 30141
rect 26792 30064 26844 30116
rect 19800 30039 19852 30048
rect 19800 30005 19809 30039
rect 19809 30005 19843 30039
rect 19843 30005 19852 30039
rect 19800 29996 19852 30005
rect 25596 29996 25648 30048
rect 28080 29996 28132 30048
rect 28264 30039 28316 30048
rect 28264 30005 28273 30039
rect 28273 30005 28307 30039
rect 28307 30005 28316 30039
rect 28264 29996 28316 30005
rect 5915 29894 5967 29946
rect 5979 29894 6031 29946
rect 6043 29894 6095 29946
rect 6107 29894 6159 29946
rect 6171 29894 6223 29946
rect 15846 29894 15898 29946
rect 15910 29894 15962 29946
rect 15974 29894 16026 29946
rect 16038 29894 16090 29946
rect 16102 29894 16154 29946
rect 25776 29894 25828 29946
rect 25840 29894 25892 29946
rect 25904 29894 25956 29946
rect 25968 29894 26020 29946
rect 26032 29894 26084 29946
rect 4068 29792 4120 29844
rect 17040 29835 17092 29844
rect 17040 29801 17049 29835
rect 17049 29801 17083 29835
rect 17083 29801 17092 29835
rect 17040 29792 17092 29801
rect 18696 29835 18748 29844
rect 18696 29801 18705 29835
rect 18705 29801 18739 29835
rect 18739 29801 18748 29835
rect 18696 29792 18748 29801
rect 19892 29835 19944 29844
rect 19892 29801 19901 29835
rect 19901 29801 19935 29835
rect 19935 29801 19944 29835
rect 19892 29792 19944 29801
rect 25688 29792 25740 29844
rect 26792 29792 26844 29844
rect 27344 29792 27396 29844
rect 27804 29792 27856 29844
rect 30012 29835 30064 29844
rect 2136 29588 2188 29640
rect 25964 29724 26016 29776
rect 20720 29656 20772 29708
rect 12716 29631 12768 29640
rect 12716 29597 12725 29631
rect 12725 29597 12759 29631
rect 12759 29597 12768 29631
rect 12716 29588 12768 29597
rect 13084 29588 13136 29640
rect 14372 29631 14424 29640
rect 14372 29597 14395 29631
rect 14395 29597 14424 29631
rect 14372 29588 14424 29597
rect 14648 29588 14700 29640
rect 14740 29631 14792 29640
rect 14740 29597 14749 29631
rect 14749 29597 14783 29631
rect 14783 29597 14792 29631
rect 15752 29631 15804 29640
rect 14740 29588 14792 29597
rect 15752 29597 15761 29631
rect 15761 29597 15795 29631
rect 15795 29597 15804 29631
rect 15752 29588 15804 29597
rect 18788 29588 18840 29640
rect 19800 29588 19852 29640
rect 22100 29656 22152 29708
rect 22744 29656 22796 29708
rect 25596 29656 25648 29708
rect 1584 29495 1636 29504
rect 1584 29461 1593 29495
rect 1593 29461 1627 29495
rect 1627 29461 1636 29495
rect 1584 29452 1636 29461
rect 2136 29495 2188 29504
rect 2136 29461 2145 29495
rect 2145 29461 2179 29495
rect 2179 29461 2188 29495
rect 2136 29452 2188 29461
rect 14188 29452 14240 29504
rect 14464 29452 14516 29504
rect 19984 29452 20036 29504
rect 22836 29588 22888 29640
rect 25872 29588 25924 29640
rect 21364 29520 21416 29572
rect 22008 29520 22060 29572
rect 23112 29520 23164 29572
rect 26056 29520 26108 29572
rect 27068 29588 27120 29640
rect 28172 29724 28224 29776
rect 30012 29801 30021 29835
rect 30021 29801 30055 29835
rect 30055 29801 30064 29835
rect 30012 29792 30064 29801
rect 28080 29656 28132 29708
rect 28356 29588 28408 29640
rect 27712 29520 27764 29572
rect 21548 29452 21600 29504
rect 25872 29452 25924 29504
rect 26332 29452 26384 29504
rect 27252 29452 27304 29504
rect 27620 29495 27672 29504
rect 27620 29461 27629 29495
rect 27629 29461 27663 29495
rect 27663 29461 27672 29495
rect 28908 29495 28960 29504
rect 27620 29452 27672 29461
rect 28908 29461 28917 29495
rect 28917 29461 28951 29495
rect 28951 29461 28960 29495
rect 28908 29452 28960 29461
rect 10880 29350 10932 29402
rect 10944 29350 10996 29402
rect 11008 29350 11060 29402
rect 11072 29350 11124 29402
rect 11136 29350 11188 29402
rect 20811 29350 20863 29402
rect 20875 29350 20927 29402
rect 20939 29350 20991 29402
rect 21003 29350 21055 29402
rect 21067 29350 21119 29402
rect 15108 29248 15160 29300
rect 16856 29248 16908 29300
rect 21916 29248 21968 29300
rect 22836 29291 22888 29300
rect 22836 29257 22845 29291
rect 22845 29257 22879 29291
rect 22879 29257 22888 29291
rect 22836 29248 22888 29257
rect 23388 29248 23440 29300
rect 25136 29248 25188 29300
rect 1676 29112 1728 29164
rect 12624 29112 12676 29164
rect 13084 29180 13136 29232
rect 13912 29223 13964 29232
rect 13912 29189 13921 29223
rect 13921 29189 13955 29223
rect 13955 29189 13964 29223
rect 13912 29180 13964 29189
rect 16948 29223 17000 29232
rect 16948 29189 16982 29223
rect 16982 29189 17000 29223
rect 16948 29180 17000 29189
rect 13360 29112 13412 29164
rect 13728 29112 13780 29164
rect 15752 29112 15804 29164
rect 19616 29180 19668 29232
rect 19984 29180 20036 29232
rect 20996 29180 21048 29232
rect 21640 29180 21692 29232
rect 19524 29155 19576 29164
rect 19524 29121 19533 29155
rect 19533 29121 19567 29155
rect 19567 29121 19576 29155
rect 19524 29112 19576 29121
rect 21548 29112 21600 29164
rect 22744 29180 22796 29232
rect 22376 29112 22428 29164
rect 22652 29112 22704 29164
rect 23112 29155 23164 29164
rect 23112 29121 23121 29155
rect 23121 29121 23155 29155
rect 23155 29121 23164 29155
rect 25596 29180 25648 29232
rect 27252 29180 27304 29232
rect 23112 29112 23164 29121
rect 14648 29044 14700 29096
rect 16672 29087 16724 29096
rect 16672 29053 16681 29087
rect 16681 29053 16715 29087
rect 16715 29053 16724 29087
rect 16672 29044 16724 29053
rect 22836 29044 22888 29096
rect 26056 29112 26108 29164
rect 27712 29248 27764 29300
rect 28172 29248 28224 29300
rect 28356 29291 28408 29300
rect 28356 29257 28365 29291
rect 28365 29257 28399 29291
rect 28399 29257 28408 29291
rect 28356 29248 28408 29257
rect 30104 29248 30156 29300
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 12348 28976 12400 29028
rect 21824 28976 21876 29028
rect 27712 29112 27764 29164
rect 27252 29044 27304 29096
rect 27528 29044 27580 29096
rect 27988 29112 28040 29164
rect 28356 29112 28408 29164
rect 29460 29112 29512 29164
rect 30012 29112 30064 29164
rect 31392 29044 31444 29096
rect 10600 28908 10652 28960
rect 17316 28908 17368 28960
rect 21180 28908 21232 28960
rect 22008 28908 22060 28960
rect 28632 28976 28684 29028
rect 27620 28908 27672 28960
rect 29460 28908 29512 28960
rect 5915 28806 5967 28858
rect 5979 28806 6031 28858
rect 6043 28806 6095 28858
rect 6107 28806 6159 28858
rect 6171 28806 6223 28858
rect 15846 28806 15898 28858
rect 15910 28806 15962 28858
rect 15974 28806 16026 28858
rect 16038 28806 16090 28858
rect 16102 28806 16154 28858
rect 25776 28806 25828 28858
rect 25840 28806 25892 28858
rect 25904 28806 25956 28858
rect 25968 28806 26020 28858
rect 26032 28806 26084 28858
rect 16672 28704 16724 28756
rect 19616 28704 19668 28756
rect 20352 28704 20404 28756
rect 25136 28747 25188 28756
rect 25136 28713 25145 28747
rect 25145 28713 25179 28747
rect 25179 28713 25188 28747
rect 25136 28704 25188 28713
rect 27620 28704 27672 28756
rect 28816 28704 28868 28756
rect 14464 28636 14516 28688
rect 17316 28636 17368 28688
rect 2136 28500 2188 28552
rect 14648 28568 14700 28620
rect 2228 28432 2280 28484
rect 10784 28432 10836 28484
rect 14740 28543 14792 28552
rect 14740 28509 14749 28543
rect 14749 28509 14783 28543
rect 14783 28509 14792 28543
rect 14740 28500 14792 28509
rect 15476 28500 15528 28552
rect 17592 28568 17644 28620
rect 20076 28568 20128 28620
rect 17040 28500 17092 28552
rect 18328 28500 18380 28552
rect 16488 28432 16540 28484
rect 19708 28500 19760 28552
rect 19616 28432 19668 28484
rect 20076 28475 20128 28484
rect 20076 28441 20085 28475
rect 20085 28441 20119 28475
rect 20119 28441 20128 28475
rect 20076 28432 20128 28441
rect 20536 28636 20588 28688
rect 20996 28543 21048 28552
rect 20996 28509 21005 28543
rect 21005 28509 21039 28543
rect 21039 28509 21048 28543
rect 20996 28500 21048 28509
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 21824 28500 21876 28552
rect 22008 28543 22060 28552
rect 22008 28509 22017 28543
rect 22017 28509 22051 28543
rect 22051 28509 22060 28543
rect 22008 28500 22060 28509
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 15292 28364 15344 28416
rect 15384 28364 15436 28416
rect 16948 28407 17000 28416
rect 16948 28373 16957 28407
rect 16957 28373 16991 28407
rect 16991 28373 17000 28407
rect 16948 28364 17000 28373
rect 19524 28407 19576 28416
rect 19524 28373 19533 28407
rect 19533 28373 19567 28407
rect 19567 28373 19576 28407
rect 19524 28364 19576 28373
rect 20168 28407 20220 28416
rect 20168 28373 20177 28407
rect 20177 28373 20211 28407
rect 20211 28373 20220 28407
rect 20168 28364 20220 28373
rect 21272 28364 21324 28416
rect 21548 28364 21600 28416
rect 25136 28500 25188 28552
rect 24768 28475 24820 28484
rect 24768 28441 24777 28475
rect 24777 28441 24811 28475
rect 24811 28441 24820 28475
rect 24768 28432 24820 28441
rect 25044 28432 25096 28484
rect 29644 28636 29696 28688
rect 30104 28636 30156 28688
rect 28632 28568 28684 28620
rect 29092 28568 29144 28620
rect 27620 28500 27672 28552
rect 27988 28500 28040 28552
rect 28080 28500 28132 28552
rect 26792 28432 26844 28484
rect 27252 28407 27304 28416
rect 27252 28373 27261 28407
rect 27261 28373 27295 28407
rect 27295 28373 27304 28407
rect 27252 28364 27304 28373
rect 27988 28364 28040 28416
rect 28448 28364 28500 28416
rect 29000 28364 29052 28416
rect 29644 28500 29696 28552
rect 30012 28407 30064 28416
rect 30012 28373 30021 28407
rect 30021 28373 30055 28407
rect 30055 28373 30064 28407
rect 30012 28364 30064 28373
rect 10880 28262 10932 28314
rect 10944 28262 10996 28314
rect 11008 28262 11060 28314
rect 11072 28262 11124 28314
rect 11136 28262 11188 28314
rect 20811 28262 20863 28314
rect 20875 28262 20927 28314
rect 20939 28262 20991 28314
rect 21003 28262 21055 28314
rect 21067 28262 21119 28314
rect 13820 28160 13872 28212
rect 15844 28160 15896 28212
rect 20536 28160 20588 28212
rect 23204 28160 23256 28212
rect 23572 28160 23624 28212
rect 24032 28203 24084 28212
rect 24032 28169 24041 28203
rect 24041 28169 24075 28203
rect 24075 28169 24084 28203
rect 24032 28160 24084 28169
rect 25596 28160 25648 28212
rect 28448 28160 28500 28212
rect 28632 28160 28684 28212
rect 29368 28203 29420 28212
rect 13544 28092 13596 28144
rect 16488 28092 16540 28144
rect 15660 28024 15712 28076
rect 20168 28092 20220 28144
rect 23112 28092 23164 28144
rect 26792 28092 26844 28144
rect 27252 28092 27304 28144
rect 19524 28024 19576 28076
rect 22008 28024 22060 28076
rect 22468 28024 22520 28076
rect 23204 28024 23256 28076
rect 23848 28024 23900 28076
rect 25136 28024 25188 28076
rect 15752 27956 15804 28008
rect 28448 28024 28500 28076
rect 15476 27931 15528 27940
rect 15476 27897 15485 27931
rect 15485 27897 15519 27931
rect 15519 27897 15528 27931
rect 15476 27888 15528 27897
rect 27712 27931 27764 27940
rect 27712 27897 27721 27931
rect 27721 27897 27755 27931
rect 27755 27897 27764 27931
rect 27712 27888 27764 27897
rect 18328 27820 18380 27872
rect 19432 27820 19484 27872
rect 23572 27820 23624 27872
rect 28816 28024 28868 28076
rect 29368 28169 29377 28203
rect 29377 28169 29411 28203
rect 29411 28169 29420 28203
rect 29368 28160 29420 28169
rect 29460 28160 29512 28212
rect 29368 27956 29420 28008
rect 29552 27956 29604 28008
rect 31484 27820 31536 27872
rect 5915 27718 5967 27770
rect 5979 27718 6031 27770
rect 6043 27718 6095 27770
rect 6107 27718 6159 27770
rect 6171 27718 6223 27770
rect 15846 27718 15898 27770
rect 15910 27718 15962 27770
rect 15974 27718 16026 27770
rect 16038 27718 16090 27770
rect 16102 27718 16154 27770
rect 25776 27718 25828 27770
rect 25840 27718 25892 27770
rect 25904 27718 25956 27770
rect 25968 27718 26020 27770
rect 26032 27718 26084 27770
rect 15384 27616 15436 27668
rect 21548 27659 21600 27668
rect 21548 27625 21557 27659
rect 21557 27625 21591 27659
rect 21591 27625 21600 27659
rect 21548 27616 21600 27625
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 12072 27455 12124 27464
rect 12072 27421 12081 27455
rect 12081 27421 12115 27455
rect 12115 27421 12124 27455
rect 12072 27412 12124 27421
rect 12348 27455 12400 27464
rect 12348 27421 12382 27455
rect 12382 27421 12400 27455
rect 12348 27412 12400 27421
rect 25412 27548 25464 27600
rect 25780 27548 25832 27600
rect 26700 27616 26752 27668
rect 21824 27480 21876 27532
rect 21640 27455 21692 27464
rect 21640 27421 21649 27455
rect 21649 27421 21683 27455
rect 21683 27421 21692 27455
rect 21640 27412 21692 27421
rect 24584 27412 24636 27464
rect 25136 27455 25188 27464
rect 25136 27421 25145 27455
rect 25145 27421 25179 27455
rect 25179 27421 25188 27455
rect 25136 27412 25188 27421
rect 25412 27412 25464 27464
rect 25780 27455 25832 27464
rect 25780 27421 25789 27455
rect 25789 27421 25823 27455
rect 25823 27421 25832 27455
rect 25780 27412 25832 27421
rect 26516 27480 26568 27532
rect 26700 27480 26752 27532
rect 26148 27412 26200 27464
rect 27436 27455 27488 27464
rect 27436 27421 27445 27455
rect 27445 27421 27479 27455
rect 27479 27421 27488 27455
rect 27436 27412 27488 27421
rect 28080 27548 28132 27600
rect 29460 27548 29512 27600
rect 31484 27548 31536 27600
rect 31760 27548 31812 27600
rect 27712 27523 27764 27532
rect 27712 27489 27721 27523
rect 27721 27489 27755 27523
rect 27755 27489 27764 27523
rect 27712 27480 27764 27489
rect 28264 27480 28316 27532
rect 15292 27387 15344 27396
rect 15292 27353 15326 27387
rect 15326 27353 15344 27387
rect 15292 27344 15344 27353
rect 15752 27344 15804 27396
rect 16948 27344 17000 27396
rect 17592 27387 17644 27396
rect 17592 27353 17601 27387
rect 17601 27353 17635 27387
rect 17635 27353 17644 27387
rect 17592 27344 17644 27353
rect 21456 27344 21508 27396
rect 21916 27344 21968 27396
rect 24676 27344 24728 27396
rect 26516 27344 26568 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 12808 27276 12860 27328
rect 16488 27276 16540 27328
rect 22008 27276 22060 27328
rect 22376 27276 22428 27328
rect 22560 27276 22612 27328
rect 24216 27276 24268 27328
rect 24584 27276 24636 27328
rect 27528 27276 27580 27328
rect 28448 27412 28500 27464
rect 28908 27412 28960 27464
rect 31024 27412 31076 27464
rect 31760 27412 31812 27464
rect 29368 27344 29420 27396
rect 28080 27276 28132 27328
rect 28448 27276 28500 27328
rect 28908 27319 28960 27328
rect 28908 27285 28917 27319
rect 28917 27285 28951 27319
rect 28951 27285 28960 27319
rect 28908 27276 28960 27285
rect 10880 27174 10932 27226
rect 10944 27174 10996 27226
rect 11008 27174 11060 27226
rect 11072 27174 11124 27226
rect 11136 27174 11188 27226
rect 20811 27174 20863 27226
rect 20875 27174 20927 27226
rect 20939 27174 20991 27226
rect 21003 27174 21055 27226
rect 21067 27174 21119 27226
rect 2320 27072 2372 27124
rect 12072 27072 12124 27124
rect 15016 27004 15068 27056
rect 12532 26936 12584 26988
rect 16488 27072 16540 27124
rect 22284 27072 22336 27124
rect 22560 27072 22612 27124
rect 23204 27115 23256 27124
rect 23204 27081 23213 27115
rect 23213 27081 23247 27115
rect 23247 27081 23256 27115
rect 23204 27072 23256 27081
rect 24952 27115 25004 27124
rect 24952 27081 24961 27115
rect 24961 27081 24995 27115
rect 24995 27081 25004 27115
rect 24952 27072 25004 27081
rect 26240 27115 26292 27124
rect 26240 27081 26249 27115
rect 26249 27081 26283 27115
rect 26283 27081 26292 27115
rect 26240 27072 26292 27081
rect 27344 27072 27396 27124
rect 29184 27072 29236 27124
rect 29460 27072 29512 27124
rect 30840 27072 30892 27124
rect 15752 27004 15804 27056
rect 18880 27047 18932 27056
rect 18880 27013 18889 27047
rect 18889 27013 18923 27047
rect 18923 27013 18932 27047
rect 18880 27004 18932 27013
rect 24308 27004 24360 27056
rect 25596 27004 25648 27056
rect 25872 27004 25924 27056
rect 27252 27004 27304 27056
rect 27436 27004 27488 27056
rect 28080 27004 28132 27056
rect 22284 26979 22336 26988
rect 15752 26911 15804 26920
rect 15752 26877 15761 26911
rect 15761 26877 15795 26911
rect 15795 26877 15804 26911
rect 15752 26868 15804 26877
rect 17592 26868 17644 26920
rect 22284 26945 22293 26979
rect 22293 26945 22327 26979
rect 22327 26945 22336 26979
rect 22284 26936 22336 26945
rect 23388 26979 23440 26988
rect 23388 26945 23397 26979
rect 23397 26945 23431 26979
rect 23431 26945 23440 26979
rect 23388 26936 23440 26945
rect 24032 26936 24084 26988
rect 24400 26979 24452 26988
rect 24400 26945 24409 26979
rect 24409 26945 24443 26979
rect 24443 26945 24452 26979
rect 24400 26936 24452 26945
rect 25136 26936 25188 26988
rect 25412 26936 25464 26988
rect 27344 26936 27396 26988
rect 22468 26843 22520 26852
rect 1584 26775 1636 26784
rect 1584 26741 1593 26775
rect 1593 26741 1627 26775
rect 1627 26741 1636 26775
rect 1584 26732 1636 26741
rect 13636 26775 13688 26784
rect 13636 26741 13645 26775
rect 13645 26741 13679 26775
rect 13679 26741 13688 26775
rect 13636 26732 13688 26741
rect 15660 26732 15712 26784
rect 20168 26775 20220 26784
rect 20168 26741 20177 26775
rect 20177 26741 20211 26775
rect 20211 26741 20220 26775
rect 20168 26732 20220 26741
rect 22468 26809 22477 26843
rect 22477 26809 22511 26843
rect 22511 26809 22520 26843
rect 22468 26800 22520 26809
rect 25872 26800 25924 26852
rect 26056 26800 26108 26852
rect 26884 26868 26936 26920
rect 27160 26868 27212 26920
rect 27436 26911 27488 26920
rect 27436 26877 27445 26911
rect 27445 26877 27479 26911
rect 27479 26877 27488 26911
rect 27436 26868 27488 26877
rect 29460 26936 29512 26988
rect 30012 26911 30064 26920
rect 30012 26877 30021 26911
rect 30021 26877 30055 26911
rect 30055 26877 30064 26911
rect 30012 26868 30064 26877
rect 30564 26868 30616 26920
rect 30932 26868 30984 26920
rect 23664 26732 23716 26784
rect 24860 26732 24912 26784
rect 26240 26732 26292 26784
rect 26884 26732 26936 26784
rect 29184 26800 29236 26852
rect 30380 26800 30432 26852
rect 29460 26775 29512 26784
rect 29460 26741 29469 26775
rect 29469 26741 29503 26775
rect 29503 26741 29512 26775
rect 29460 26732 29512 26741
rect 5915 26630 5967 26682
rect 5979 26630 6031 26682
rect 6043 26630 6095 26682
rect 6107 26630 6159 26682
rect 6171 26630 6223 26682
rect 15846 26630 15898 26682
rect 15910 26630 15962 26682
rect 15974 26630 16026 26682
rect 16038 26630 16090 26682
rect 16102 26630 16154 26682
rect 25776 26630 25828 26682
rect 25840 26630 25892 26682
rect 25904 26630 25956 26682
rect 25968 26630 26020 26682
rect 26032 26630 26084 26682
rect 15568 26528 15620 26580
rect 18052 26528 18104 26580
rect 29460 26528 29512 26580
rect 29920 26528 29972 26580
rect 27436 26460 27488 26512
rect 28080 26503 28132 26512
rect 28080 26469 28089 26503
rect 28089 26469 28123 26503
rect 28123 26469 28132 26503
rect 28080 26460 28132 26469
rect 28908 26503 28960 26512
rect 28908 26469 28917 26503
rect 28917 26469 28951 26503
rect 28951 26469 28960 26503
rect 28908 26460 28960 26469
rect 15660 26435 15712 26444
rect 15660 26401 15669 26435
rect 15669 26401 15703 26435
rect 15703 26401 15712 26435
rect 15660 26392 15712 26401
rect 31392 26460 31444 26512
rect 2320 26367 2372 26376
rect 2320 26333 2329 26367
rect 2329 26333 2363 26367
rect 2363 26333 2372 26367
rect 2320 26324 2372 26333
rect 13820 26324 13872 26376
rect 15200 26324 15252 26376
rect 22928 26324 22980 26376
rect 26148 26324 26200 26376
rect 26240 26324 26292 26376
rect 27712 26324 27764 26376
rect 30380 26324 30432 26376
rect 25504 26299 25556 26308
rect 25504 26265 25513 26299
rect 25513 26265 25547 26299
rect 25547 26265 25556 26299
rect 25504 26256 25556 26265
rect 27436 26256 27488 26308
rect 28080 26256 28132 26308
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 12992 26188 13044 26240
rect 10880 26086 10932 26138
rect 10944 26086 10996 26138
rect 11008 26086 11060 26138
rect 11072 26086 11124 26138
rect 11136 26086 11188 26138
rect 20811 26086 20863 26138
rect 20875 26086 20927 26138
rect 20939 26086 20991 26138
rect 21003 26086 21055 26138
rect 21067 26086 21119 26138
rect 13268 25984 13320 26036
rect 13636 25984 13688 26036
rect 22376 25984 22428 26036
rect 22928 25984 22980 26036
rect 23848 25984 23900 26036
rect 24124 25984 24176 26036
rect 26700 25984 26752 26036
rect 28632 26027 28684 26036
rect 28632 25993 28641 26027
rect 28641 25993 28675 26027
rect 28675 25993 28684 26027
rect 28632 25984 28684 25993
rect 29092 26027 29144 26036
rect 29092 25993 29101 26027
rect 29101 25993 29135 26027
rect 29135 25993 29144 26027
rect 29092 25984 29144 25993
rect 18052 25916 18104 25968
rect 20168 25916 20220 25968
rect 13084 25891 13136 25900
rect 13084 25857 13093 25891
rect 13093 25857 13127 25891
rect 13127 25857 13136 25891
rect 13084 25848 13136 25857
rect 19340 25891 19392 25900
rect 12992 25823 13044 25832
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 19340 25857 19349 25891
rect 19349 25857 19383 25891
rect 19383 25857 19392 25891
rect 19340 25848 19392 25857
rect 22376 25848 22428 25900
rect 22652 25916 22704 25968
rect 27344 25916 27396 25968
rect 29460 25916 29512 25968
rect 30012 25959 30064 25968
rect 30012 25925 30021 25959
rect 30021 25925 30055 25959
rect 30055 25925 30064 25959
rect 30012 25916 30064 25925
rect 22744 25891 22796 25900
rect 18512 25780 18564 25832
rect 22744 25857 22753 25891
rect 22753 25857 22787 25891
rect 22787 25857 22796 25891
rect 22744 25848 22796 25857
rect 24124 25848 24176 25900
rect 27804 25891 27856 25900
rect 27804 25857 27813 25891
rect 27813 25857 27847 25891
rect 27847 25857 27856 25891
rect 27804 25848 27856 25857
rect 28080 25848 28132 25900
rect 28448 25891 28500 25900
rect 28448 25857 28457 25891
rect 28457 25857 28491 25891
rect 28491 25857 28500 25891
rect 28448 25848 28500 25857
rect 24032 25780 24084 25832
rect 29368 25780 29420 25832
rect 12532 25755 12584 25764
rect 12532 25721 12541 25755
rect 12541 25721 12575 25755
rect 12575 25721 12584 25755
rect 12532 25712 12584 25721
rect 24400 25712 24452 25764
rect 30564 25712 30616 25764
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 17868 25644 17920 25696
rect 19616 25644 19668 25696
rect 21456 25644 21508 25696
rect 5915 25542 5967 25594
rect 5979 25542 6031 25594
rect 6043 25542 6095 25594
rect 6107 25542 6159 25594
rect 6171 25542 6223 25594
rect 15846 25542 15898 25594
rect 15910 25542 15962 25594
rect 15974 25542 16026 25594
rect 16038 25542 16090 25594
rect 16102 25542 16154 25594
rect 25776 25542 25828 25594
rect 25840 25542 25892 25594
rect 25904 25542 25956 25594
rect 25968 25542 26020 25594
rect 26032 25542 26084 25594
rect 1676 25483 1728 25492
rect 1676 25449 1685 25483
rect 1685 25449 1719 25483
rect 1719 25449 1728 25483
rect 1676 25440 1728 25449
rect 2320 25440 2372 25492
rect 24400 25440 24452 25492
rect 25504 25440 25556 25492
rect 27344 25440 27396 25492
rect 28172 25440 28224 25492
rect 30012 25483 30064 25492
rect 30012 25449 30021 25483
rect 30021 25449 30055 25483
rect 30055 25449 30064 25483
rect 30012 25440 30064 25449
rect 16856 25372 16908 25424
rect 21824 25372 21876 25424
rect 27620 25372 27672 25424
rect 18328 25304 18380 25356
rect 19616 25347 19668 25356
rect 19616 25313 19625 25347
rect 19625 25313 19659 25347
rect 19659 25313 19668 25347
rect 19616 25304 19668 25313
rect 1860 25279 1912 25288
rect 1860 25245 1869 25279
rect 1869 25245 1903 25279
rect 1903 25245 1912 25279
rect 1860 25236 1912 25245
rect 16396 25279 16448 25288
rect 16396 25245 16405 25279
rect 16405 25245 16439 25279
rect 16439 25245 16448 25279
rect 16396 25236 16448 25245
rect 18512 25279 18564 25288
rect 18512 25245 18521 25279
rect 18521 25245 18555 25279
rect 18555 25245 18564 25279
rect 18512 25236 18564 25245
rect 22376 25279 22428 25288
rect 22376 25245 22385 25279
rect 22385 25245 22419 25279
rect 22419 25245 22428 25279
rect 22376 25236 22428 25245
rect 22928 25304 22980 25356
rect 24400 25304 24452 25356
rect 26332 25304 26384 25356
rect 27344 25304 27396 25356
rect 22652 25279 22704 25288
rect 17684 25211 17736 25220
rect 17684 25177 17693 25211
rect 17693 25177 17727 25211
rect 17727 25177 17736 25211
rect 17684 25168 17736 25177
rect 17868 25211 17920 25220
rect 17868 25177 17877 25211
rect 17877 25177 17911 25211
rect 17911 25177 17920 25211
rect 17868 25168 17920 25177
rect 20628 25168 20680 25220
rect 16580 25143 16632 25152
rect 16580 25109 16589 25143
rect 16589 25109 16623 25143
rect 16623 25109 16632 25143
rect 16580 25100 16632 25109
rect 18052 25100 18104 25152
rect 21272 25100 21324 25152
rect 22376 25100 22428 25152
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 22744 25279 22796 25288
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 23940 25236 23992 25288
rect 24860 25279 24912 25288
rect 24860 25245 24869 25279
rect 24869 25245 24903 25279
rect 24903 25245 24912 25279
rect 24860 25236 24912 25245
rect 26700 25236 26752 25288
rect 28080 25236 28132 25288
rect 27620 25168 27672 25220
rect 29000 25372 29052 25424
rect 29368 25372 29420 25424
rect 29000 25279 29052 25288
rect 29000 25245 29009 25279
rect 29009 25245 29043 25279
rect 29043 25245 29052 25279
rect 29000 25236 29052 25245
rect 30840 25236 30892 25288
rect 26332 25100 26384 25152
rect 27528 25100 27580 25152
rect 10880 24998 10932 25050
rect 10944 24998 10996 25050
rect 11008 24998 11060 25050
rect 11072 24998 11124 25050
rect 11136 24998 11188 25050
rect 20811 24998 20863 25050
rect 20875 24998 20927 25050
rect 20939 24998 20991 25050
rect 21003 24998 21055 25050
rect 21067 24998 21119 25050
rect 13268 24939 13320 24948
rect 13268 24905 13277 24939
rect 13277 24905 13311 24939
rect 13311 24905 13320 24939
rect 13268 24896 13320 24905
rect 20628 24939 20680 24948
rect 1860 24828 1912 24880
rect 2320 24803 2372 24812
rect 1584 24667 1636 24676
rect 1584 24633 1593 24667
rect 1593 24633 1627 24667
rect 1627 24633 1636 24667
rect 1584 24624 1636 24633
rect 2320 24769 2329 24803
rect 2329 24769 2363 24803
rect 2363 24769 2372 24803
rect 2320 24760 2372 24769
rect 12992 24828 13044 24880
rect 14004 24760 14056 24812
rect 18604 24828 18656 24880
rect 20628 24905 20637 24939
rect 20637 24905 20671 24939
rect 20671 24905 20680 24939
rect 20628 24896 20680 24905
rect 13084 24692 13136 24744
rect 13452 24692 13504 24744
rect 13912 24735 13964 24744
rect 13912 24701 13921 24735
rect 13921 24701 13955 24735
rect 13955 24701 13964 24735
rect 13912 24692 13964 24701
rect 15384 24624 15436 24676
rect 14096 24556 14148 24608
rect 16948 24556 17000 24608
rect 17500 24803 17552 24812
rect 17500 24769 17509 24803
rect 17509 24769 17543 24803
rect 17543 24769 17552 24803
rect 17500 24760 17552 24769
rect 18052 24760 18104 24812
rect 19248 24760 19300 24812
rect 21272 24803 21324 24812
rect 17868 24692 17920 24744
rect 18144 24556 18196 24608
rect 19524 24556 19576 24608
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 22100 24760 22152 24812
rect 22928 24760 22980 24812
rect 23296 24803 23348 24812
rect 23296 24769 23305 24803
rect 23305 24769 23339 24803
rect 23339 24769 23348 24803
rect 23296 24760 23348 24769
rect 21824 24735 21876 24744
rect 21824 24701 21833 24735
rect 21833 24701 21867 24735
rect 21867 24701 21876 24735
rect 21824 24692 21876 24701
rect 22008 24692 22060 24744
rect 22652 24692 22704 24744
rect 21364 24624 21416 24676
rect 23940 24896 23992 24948
rect 26700 24896 26752 24948
rect 24308 24803 24360 24812
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 27804 24828 27856 24880
rect 24400 24692 24452 24744
rect 26240 24760 26292 24812
rect 28908 24896 28960 24948
rect 29092 24896 29144 24948
rect 24584 24692 24636 24744
rect 25320 24735 25372 24744
rect 25320 24701 25329 24735
rect 25329 24701 25363 24735
rect 25363 24701 25372 24735
rect 25320 24692 25372 24701
rect 29460 24760 29512 24812
rect 27620 24692 27672 24744
rect 29092 24692 29144 24744
rect 30380 24692 30432 24744
rect 21272 24556 21324 24608
rect 22744 24556 22796 24608
rect 24860 24556 24912 24608
rect 27344 24556 27396 24608
rect 27988 24556 28040 24608
rect 28264 24556 28316 24608
rect 28724 24556 28776 24608
rect 29460 24599 29512 24608
rect 29460 24565 29469 24599
rect 29469 24565 29503 24599
rect 29503 24565 29512 24599
rect 29460 24556 29512 24565
rect 5915 24454 5967 24506
rect 5979 24454 6031 24506
rect 6043 24454 6095 24506
rect 6107 24454 6159 24506
rect 6171 24454 6223 24506
rect 15846 24454 15898 24506
rect 15910 24454 15962 24506
rect 15974 24454 16026 24506
rect 16038 24454 16090 24506
rect 16102 24454 16154 24506
rect 25776 24454 25828 24506
rect 25840 24454 25892 24506
rect 25904 24454 25956 24506
rect 25968 24454 26020 24506
rect 26032 24454 26084 24506
rect 13912 24352 13964 24404
rect 13176 24284 13228 24336
rect 17684 24352 17736 24404
rect 19248 24395 19300 24404
rect 19248 24361 19257 24395
rect 19257 24361 19291 24395
rect 19291 24361 19300 24395
rect 19248 24352 19300 24361
rect 22284 24352 22336 24404
rect 24124 24352 24176 24404
rect 27344 24352 27396 24404
rect 27528 24352 27580 24404
rect 27804 24352 27856 24404
rect 28632 24352 28684 24404
rect 29000 24352 29052 24404
rect 29184 24352 29236 24404
rect 29460 24284 29512 24336
rect 18972 24216 19024 24268
rect 12992 24148 13044 24200
rect 13452 24191 13504 24200
rect 13452 24157 13461 24191
rect 13461 24157 13495 24191
rect 13495 24157 13504 24191
rect 13452 24148 13504 24157
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 16580 24148 16632 24200
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 13268 24080 13320 24132
rect 16948 24080 17000 24132
rect 19616 24080 19668 24132
rect 19800 24191 19852 24200
rect 19800 24157 19809 24191
rect 19809 24157 19843 24191
rect 19843 24157 19852 24191
rect 21088 24191 21140 24200
rect 19800 24148 19852 24157
rect 21088 24157 21097 24191
rect 21097 24157 21131 24191
rect 21131 24157 21140 24191
rect 21088 24148 21140 24157
rect 22100 24216 22152 24268
rect 23848 24216 23900 24268
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 22928 24148 22980 24200
rect 21364 24080 21416 24132
rect 22008 24123 22060 24132
rect 22008 24089 22017 24123
rect 22017 24089 22051 24123
rect 22051 24089 22060 24123
rect 22008 24080 22060 24089
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 20720 24012 20772 24064
rect 22192 24012 22244 24064
rect 22744 24012 22796 24064
rect 23940 24148 23992 24200
rect 23572 24080 23624 24132
rect 25412 24148 25464 24200
rect 26700 24148 26752 24200
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 28908 24148 28960 24200
rect 29920 24123 29972 24132
rect 29920 24089 29929 24123
rect 29929 24089 29963 24123
rect 29963 24089 29972 24123
rect 29920 24080 29972 24089
rect 24952 24012 25004 24064
rect 26700 24012 26752 24064
rect 27804 24012 27856 24064
rect 10880 23910 10932 23962
rect 10944 23910 10996 23962
rect 11008 23910 11060 23962
rect 11072 23910 11124 23962
rect 11136 23910 11188 23962
rect 20811 23910 20863 23962
rect 20875 23910 20927 23962
rect 20939 23910 20991 23962
rect 21003 23910 21055 23962
rect 21067 23910 21119 23962
rect 10784 23808 10836 23860
rect 14280 23808 14332 23860
rect 17500 23808 17552 23860
rect 18144 23808 18196 23860
rect 22652 23808 22704 23860
rect 22836 23808 22888 23860
rect 23112 23808 23164 23860
rect 24676 23808 24728 23860
rect 25412 23851 25464 23860
rect 25412 23817 25421 23851
rect 25421 23817 25455 23851
rect 25455 23817 25464 23851
rect 25412 23808 25464 23817
rect 12992 23672 13044 23724
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 17684 23672 17736 23724
rect 18512 23672 18564 23724
rect 19156 23672 19208 23724
rect 21180 23672 21232 23724
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 21916 23672 21968 23724
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22744 23672 22796 23724
rect 24584 23715 24636 23724
rect 24584 23681 24593 23715
rect 24593 23681 24627 23715
rect 24627 23681 24636 23715
rect 24584 23672 24636 23681
rect 24952 23672 25004 23724
rect 27620 23740 27672 23792
rect 28448 23740 28500 23792
rect 28632 23715 28684 23724
rect 28632 23681 28641 23715
rect 28641 23681 28675 23715
rect 28675 23681 28684 23715
rect 28632 23672 28684 23681
rect 29184 23715 29236 23724
rect 29184 23681 29193 23715
rect 29193 23681 29227 23715
rect 29227 23681 29236 23715
rect 29184 23672 29236 23681
rect 22100 23604 22152 23656
rect 17868 23536 17920 23588
rect 21916 23536 21968 23588
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 14096 23468 14148 23520
rect 19708 23511 19760 23520
rect 19708 23477 19717 23511
rect 19717 23477 19751 23511
rect 19751 23477 19760 23511
rect 19708 23468 19760 23477
rect 24124 23604 24176 23656
rect 23112 23536 23164 23588
rect 25412 23604 25464 23656
rect 27804 23604 27856 23656
rect 27988 23579 28040 23588
rect 27988 23545 27997 23579
rect 27997 23545 28031 23579
rect 28031 23545 28040 23579
rect 27988 23536 28040 23545
rect 29000 23536 29052 23588
rect 23572 23468 23624 23520
rect 24676 23468 24728 23520
rect 24860 23468 24912 23520
rect 28724 23468 28776 23520
rect 5915 23366 5967 23418
rect 5979 23366 6031 23418
rect 6043 23366 6095 23418
rect 6107 23366 6159 23418
rect 6171 23366 6223 23418
rect 15846 23366 15898 23418
rect 15910 23366 15962 23418
rect 15974 23366 16026 23418
rect 16038 23366 16090 23418
rect 16102 23366 16154 23418
rect 25776 23366 25828 23418
rect 25840 23366 25892 23418
rect 25904 23366 25956 23418
rect 25968 23366 26020 23418
rect 26032 23366 26084 23418
rect 12992 23264 13044 23316
rect 22652 23264 22704 23316
rect 23296 23307 23348 23316
rect 23296 23273 23305 23307
rect 23305 23273 23339 23307
rect 23339 23273 23348 23307
rect 23296 23264 23348 23273
rect 24768 23264 24820 23316
rect 24860 23264 24912 23316
rect 25320 23264 25372 23316
rect 15476 23239 15528 23248
rect 15476 23205 15485 23239
rect 15485 23205 15519 23239
rect 15519 23205 15528 23239
rect 15476 23196 15528 23205
rect 14096 23171 14148 23180
rect 14096 23137 14105 23171
rect 14105 23137 14139 23171
rect 14139 23137 14148 23171
rect 14096 23128 14148 23137
rect 19708 23128 19760 23180
rect 2320 23103 2372 23112
rect 2320 23069 2329 23103
rect 2329 23069 2363 23103
rect 2363 23069 2372 23103
rect 2320 23060 2372 23069
rect 14188 23060 14240 23112
rect 17132 23060 17184 23112
rect 21180 23128 21232 23180
rect 21548 23060 21600 23112
rect 22836 23128 22888 23180
rect 29368 23264 29420 23316
rect 20720 22992 20772 23044
rect 22376 23060 22428 23112
rect 22928 23103 22980 23112
rect 22928 23069 22937 23103
rect 22937 23069 22971 23103
rect 22971 23069 22980 23103
rect 22928 23060 22980 23069
rect 23848 23060 23900 23112
rect 24584 23103 24636 23112
rect 24584 23069 24593 23103
rect 24593 23069 24627 23103
rect 24627 23069 24636 23103
rect 24584 23060 24636 23069
rect 24676 23060 24728 23112
rect 25412 23060 25464 23112
rect 27620 23128 27672 23180
rect 29368 23128 29420 23180
rect 26148 23060 26200 23112
rect 28908 23060 28960 23112
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 24952 22992 25004 23044
rect 25136 22992 25188 23044
rect 27620 22992 27672 23044
rect 29000 22992 29052 23044
rect 23020 22924 23072 22976
rect 23572 22924 23624 22976
rect 24768 22924 24820 22976
rect 25320 22924 25372 22976
rect 26700 22924 26752 22976
rect 29092 22924 29144 22976
rect 29276 22924 29328 22976
rect 10880 22822 10932 22874
rect 10944 22822 10996 22874
rect 11008 22822 11060 22874
rect 11072 22822 11124 22874
rect 11136 22822 11188 22874
rect 20811 22822 20863 22874
rect 20875 22822 20927 22874
rect 20939 22822 20991 22874
rect 21003 22822 21055 22874
rect 21067 22822 21119 22874
rect 2320 22720 2372 22772
rect 17132 22720 17184 22772
rect 18144 22720 18196 22772
rect 22192 22720 22244 22772
rect 22652 22720 22704 22772
rect 29828 22763 29880 22772
rect 29828 22729 29837 22763
rect 29837 22729 29871 22763
rect 29871 22729 29880 22763
rect 29828 22720 29880 22729
rect 22100 22652 22152 22704
rect 17868 22627 17920 22636
rect 17868 22593 17877 22627
rect 17877 22593 17911 22627
rect 17911 22593 17920 22627
rect 17868 22584 17920 22593
rect 21180 22584 21232 22636
rect 21640 22584 21692 22636
rect 22376 22652 22428 22704
rect 26700 22652 26752 22704
rect 21364 22516 21416 22568
rect 22928 22584 22980 22636
rect 23204 22584 23256 22636
rect 23480 22584 23532 22636
rect 23940 22584 23992 22636
rect 24308 22584 24360 22636
rect 25412 22627 25464 22636
rect 25136 22516 25188 22568
rect 25412 22593 25421 22627
rect 25421 22593 25455 22627
rect 25455 22593 25464 22627
rect 25412 22584 25464 22593
rect 26240 22584 26292 22636
rect 27620 22695 27672 22704
rect 27620 22661 27629 22695
rect 27629 22661 27663 22695
rect 27663 22661 27672 22695
rect 27620 22652 27672 22661
rect 29000 22584 29052 22636
rect 28632 22516 28684 22568
rect 29368 22652 29420 22704
rect 29460 22627 29512 22636
rect 29460 22593 29469 22627
rect 29469 22593 29503 22627
rect 29503 22593 29512 22627
rect 29460 22584 29512 22593
rect 31484 22516 31536 22568
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 21272 22380 21324 22432
rect 22376 22448 22428 22500
rect 25320 22380 25372 22432
rect 25596 22423 25648 22432
rect 25596 22389 25605 22423
rect 25605 22389 25639 22423
rect 25639 22389 25648 22423
rect 25596 22380 25648 22389
rect 26700 22380 26752 22432
rect 28724 22380 28776 22432
rect 5915 22278 5967 22330
rect 5979 22278 6031 22330
rect 6043 22278 6095 22330
rect 6107 22278 6159 22330
rect 6171 22278 6223 22330
rect 15846 22278 15898 22330
rect 15910 22278 15962 22330
rect 15974 22278 16026 22330
rect 16038 22278 16090 22330
rect 16102 22278 16154 22330
rect 25776 22278 25828 22330
rect 25840 22278 25892 22330
rect 25904 22278 25956 22330
rect 25968 22278 26020 22330
rect 26032 22278 26084 22330
rect 22100 22176 22152 22228
rect 22560 22176 22612 22228
rect 26240 22176 26292 22228
rect 26792 22176 26844 22228
rect 27528 22176 27580 22228
rect 28448 22176 28500 22228
rect 28908 22176 28960 22228
rect 27436 22108 27488 22160
rect 18512 21972 18564 22024
rect 22284 21972 22336 22024
rect 22744 21904 22796 21956
rect 23112 21904 23164 21956
rect 26240 22040 26292 22092
rect 27712 22040 27764 22092
rect 28632 22040 28684 22092
rect 25320 22015 25372 22024
rect 25320 21981 25354 22015
rect 25354 21981 25372 22015
rect 25320 21972 25372 21981
rect 28264 21972 28316 22024
rect 30288 22040 30340 22092
rect 29368 21972 29420 22024
rect 29920 21972 29972 22024
rect 25596 21904 25648 21956
rect 26148 21904 26200 21956
rect 27252 21947 27304 21956
rect 27252 21913 27261 21947
rect 27261 21913 27295 21947
rect 27295 21913 27304 21947
rect 27252 21904 27304 21913
rect 27804 21947 27856 21956
rect 27804 21913 27813 21947
rect 27813 21913 27847 21947
rect 27847 21913 27856 21947
rect 27804 21904 27856 21913
rect 28448 21947 28500 21956
rect 28448 21913 28457 21947
rect 28457 21913 28491 21947
rect 28491 21913 28500 21947
rect 28448 21904 28500 21913
rect 28816 21904 28868 21956
rect 29644 21947 29696 21956
rect 29644 21913 29653 21947
rect 29653 21913 29687 21947
rect 29687 21913 29696 21947
rect 29644 21904 29696 21913
rect 30012 21904 30064 21956
rect 1400 21836 1452 21888
rect 19248 21836 19300 21888
rect 22560 21879 22612 21888
rect 22560 21845 22569 21879
rect 22569 21845 22603 21879
rect 22603 21845 22612 21879
rect 22560 21836 22612 21845
rect 24400 21836 24452 21888
rect 29184 21836 29236 21888
rect 30564 21836 30616 21888
rect 10880 21734 10932 21786
rect 10944 21734 10996 21786
rect 11008 21734 11060 21786
rect 11072 21734 11124 21786
rect 11136 21734 11188 21786
rect 20811 21734 20863 21786
rect 20875 21734 20927 21786
rect 20939 21734 20991 21786
rect 21003 21734 21055 21786
rect 21067 21734 21119 21786
rect 17868 21632 17920 21684
rect 23296 21632 23348 21684
rect 24768 21632 24820 21684
rect 25412 21632 25464 21684
rect 26056 21632 26108 21684
rect 26240 21632 26292 21684
rect 27712 21632 27764 21684
rect 29000 21632 29052 21684
rect 30196 21632 30248 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 16672 21539 16724 21548
rect 1584 21403 1636 21412
rect 1584 21369 1593 21403
rect 1593 21369 1627 21403
rect 1627 21369 1636 21403
rect 1584 21360 1636 21369
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 18420 21496 18472 21548
rect 18604 21496 18656 21548
rect 19248 21539 19300 21548
rect 18144 21428 18196 21480
rect 19248 21505 19257 21539
rect 19257 21505 19291 21539
rect 19291 21505 19300 21539
rect 19248 21496 19300 21505
rect 19616 21496 19668 21548
rect 22376 21496 22428 21548
rect 24584 21564 24636 21616
rect 25596 21564 25648 21616
rect 25964 21564 26016 21616
rect 27344 21564 27396 21616
rect 28632 21564 28684 21616
rect 29920 21607 29972 21616
rect 29920 21573 29929 21607
rect 29929 21573 29963 21607
rect 29963 21573 29972 21607
rect 29920 21564 29972 21573
rect 25136 21496 25188 21548
rect 25412 21539 25464 21548
rect 25412 21505 25421 21539
rect 25421 21505 25455 21539
rect 25455 21505 25464 21539
rect 25412 21496 25464 21505
rect 24860 21428 24912 21480
rect 26792 21496 26844 21548
rect 28172 21539 28224 21548
rect 28172 21505 28181 21539
rect 28181 21505 28215 21539
rect 28215 21505 28224 21539
rect 28172 21496 28224 21505
rect 29276 21539 29328 21548
rect 29276 21505 29285 21539
rect 29285 21505 29319 21539
rect 29319 21505 29328 21539
rect 29276 21496 29328 21505
rect 29368 21428 29420 21480
rect 30196 21428 30248 21480
rect 24400 21360 24452 21412
rect 1400 21292 1452 21344
rect 16672 21292 16724 21344
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 18512 21335 18564 21344
rect 18512 21301 18521 21335
rect 18521 21301 18555 21335
rect 18555 21301 18564 21335
rect 18512 21292 18564 21301
rect 19340 21292 19392 21344
rect 5915 21190 5967 21242
rect 5979 21190 6031 21242
rect 6043 21190 6095 21242
rect 6107 21190 6159 21242
rect 6171 21190 6223 21242
rect 15846 21190 15898 21242
rect 15910 21190 15962 21242
rect 15974 21190 16026 21242
rect 16038 21190 16090 21242
rect 16102 21190 16154 21242
rect 25776 21190 25828 21242
rect 25840 21190 25892 21242
rect 25904 21190 25956 21242
rect 25968 21190 26020 21242
rect 26032 21190 26084 21242
rect 12716 21088 12768 21140
rect 23572 21088 23624 21140
rect 27436 21131 27488 21140
rect 27436 21097 27445 21131
rect 27445 21097 27479 21131
rect 27479 21097 27488 21131
rect 27436 21088 27488 21097
rect 29184 21088 29236 21140
rect 30104 21131 30156 21140
rect 30104 21097 30113 21131
rect 30113 21097 30147 21131
rect 30147 21097 30156 21131
rect 30104 21088 30156 21097
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 18052 20952 18104 21004
rect 17776 20884 17828 20936
rect 19340 20884 19392 20936
rect 24584 20927 24636 20936
rect 24584 20893 24593 20927
rect 24593 20893 24627 20927
rect 24627 20893 24636 20927
rect 24584 20884 24636 20893
rect 24860 20927 24912 20936
rect 24860 20893 24869 20927
rect 24869 20893 24903 20927
rect 24903 20893 24912 20927
rect 24860 20884 24912 20893
rect 25596 20884 25648 20936
rect 27620 20927 27672 20936
rect 27620 20893 27629 20927
rect 27629 20893 27663 20927
rect 27663 20893 27672 20927
rect 27620 20884 27672 20893
rect 28264 20927 28316 20936
rect 28264 20893 28273 20927
rect 28273 20893 28307 20927
rect 28307 20893 28316 20927
rect 28264 20884 28316 20893
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 18052 20816 18104 20868
rect 26424 20816 26476 20868
rect 26884 20816 26936 20868
rect 28816 20859 28868 20868
rect 28816 20825 28825 20859
rect 28825 20825 28859 20859
rect 28859 20825 28868 20859
rect 28816 20816 28868 20825
rect 29184 20816 29236 20868
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 20628 20791 20680 20800
rect 20628 20757 20637 20791
rect 20637 20757 20671 20791
rect 20671 20757 20680 20791
rect 20628 20748 20680 20757
rect 10880 20646 10932 20698
rect 10944 20646 10996 20698
rect 11008 20646 11060 20698
rect 11072 20646 11124 20698
rect 11136 20646 11188 20698
rect 20811 20646 20863 20698
rect 20875 20646 20927 20698
rect 20939 20646 20991 20698
rect 21003 20646 21055 20698
rect 21067 20646 21119 20698
rect 2320 20544 2372 20596
rect 31576 20544 31628 20596
rect 20628 20476 20680 20528
rect 28172 20476 28224 20528
rect 2136 20408 2188 20460
rect 16488 20408 16540 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 18052 20408 18104 20460
rect 19248 20408 19300 20460
rect 29184 20408 29236 20460
rect 17868 20340 17920 20392
rect 30012 20383 30064 20392
rect 30012 20349 30021 20383
rect 30021 20349 30055 20383
rect 30055 20349 30064 20383
rect 30012 20340 30064 20349
rect 18052 20315 18104 20324
rect 18052 20281 18061 20315
rect 18061 20281 18095 20315
rect 18095 20281 18104 20315
rect 18052 20272 18104 20281
rect 25780 20272 25832 20324
rect 27436 20272 27488 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 18236 20204 18288 20256
rect 28172 20204 28224 20256
rect 5915 20102 5967 20154
rect 5979 20102 6031 20154
rect 6043 20102 6095 20154
rect 6107 20102 6159 20154
rect 6171 20102 6223 20154
rect 15846 20102 15898 20154
rect 15910 20102 15962 20154
rect 15974 20102 16026 20154
rect 16038 20102 16090 20154
rect 16102 20102 16154 20154
rect 25776 20102 25828 20154
rect 25840 20102 25892 20154
rect 25904 20102 25956 20154
rect 25968 20102 26020 20154
rect 26032 20102 26084 20154
rect 2136 20043 2188 20052
rect 2136 20009 2145 20043
rect 2145 20009 2179 20043
rect 2179 20009 2188 20043
rect 2136 20000 2188 20009
rect 16488 20000 16540 20052
rect 19340 20000 19392 20052
rect 9680 19932 9732 19984
rect 23204 20000 23256 20052
rect 24032 20000 24084 20052
rect 28724 20000 28776 20052
rect 29000 20000 29052 20052
rect 30288 20000 30340 20052
rect 29460 19932 29512 19984
rect 29828 19932 29880 19984
rect 30196 19932 30248 19984
rect 23480 19864 23532 19916
rect 24124 19864 24176 19916
rect 2136 19796 2188 19848
rect 2320 19839 2372 19848
rect 2320 19805 2329 19839
rect 2329 19805 2363 19839
rect 2363 19805 2372 19839
rect 2320 19796 2372 19805
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 16672 19839 16724 19848
rect 16672 19805 16681 19839
rect 16681 19805 16715 19839
rect 16715 19805 16724 19839
rect 16672 19796 16724 19805
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 19248 19796 19300 19848
rect 20628 19796 20680 19848
rect 22468 19796 22520 19848
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 24860 19839 24912 19848
rect 24860 19805 24869 19839
rect 24869 19805 24903 19839
rect 24903 19805 24912 19839
rect 24860 19796 24912 19805
rect 25964 19864 26016 19916
rect 26056 19864 26108 19916
rect 27068 19864 27120 19916
rect 28264 19864 28316 19916
rect 31760 19864 31812 19916
rect 25136 19796 25188 19848
rect 27252 19796 27304 19848
rect 27988 19796 28040 19848
rect 29828 19839 29880 19848
rect 29828 19805 29837 19839
rect 29837 19805 29871 19839
rect 29871 19805 29880 19839
rect 29828 19796 29880 19805
rect 21456 19728 21508 19780
rect 22928 19728 22980 19780
rect 25504 19728 25556 19780
rect 26792 19728 26844 19780
rect 27804 19728 27856 19780
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 20720 19660 20772 19712
rect 24216 19660 24268 19712
rect 24400 19703 24452 19712
rect 24400 19669 24409 19703
rect 24409 19669 24443 19703
rect 24443 19669 24452 19703
rect 24400 19660 24452 19669
rect 30380 19728 30432 19780
rect 29184 19660 29236 19712
rect 10880 19558 10932 19610
rect 10944 19558 10996 19610
rect 11008 19558 11060 19610
rect 11072 19558 11124 19610
rect 11136 19558 11188 19610
rect 20811 19558 20863 19610
rect 20875 19558 20927 19610
rect 20939 19558 20991 19610
rect 21003 19558 21055 19610
rect 21067 19558 21119 19610
rect 2136 19499 2188 19508
rect 2136 19465 2145 19499
rect 2145 19465 2179 19499
rect 2179 19465 2188 19499
rect 2136 19456 2188 19465
rect 16672 19456 16724 19508
rect 22928 19499 22980 19508
rect 22928 19465 22937 19499
rect 22937 19465 22971 19499
rect 22971 19465 22980 19499
rect 22928 19456 22980 19465
rect 24216 19456 24268 19508
rect 28264 19456 28316 19508
rect 29184 19456 29236 19508
rect 31208 19456 31260 19508
rect 17868 19388 17920 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 18236 19320 18288 19372
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 18052 19252 18104 19304
rect 18604 19320 18656 19372
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 19248 19388 19300 19440
rect 19616 19320 19668 19372
rect 25412 19388 25464 19440
rect 27436 19388 27488 19440
rect 28172 19431 28224 19440
rect 28172 19397 28181 19431
rect 28181 19397 28215 19431
rect 28215 19397 28224 19431
rect 28172 19388 28224 19397
rect 29000 19388 29052 19440
rect 30012 19431 30064 19440
rect 30012 19397 30021 19431
rect 30021 19397 30055 19431
rect 30055 19397 30064 19431
rect 30012 19388 30064 19397
rect 21272 19320 21324 19372
rect 24400 19320 24452 19372
rect 25596 19320 25648 19372
rect 25780 19320 25832 19372
rect 23204 19252 23256 19304
rect 25136 19252 25188 19304
rect 26700 19320 26752 19372
rect 28908 19363 28960 19372
rect 28908 19329 28917 19363
rect 28917 19329 28951 19363
rect 28951 19329 28960 19363
rect 28908 19320 28960 19329
rect 29184 19320 29236 19372
rect 29644 19320 29696 19372
rect 23664 19184 23716 19236
rect 24032 19184 24084 19236
rect 25872 19184 25924 19236
rect 28908 19184 28960 19236
rect 29460 19227 29512 19236
rect 29460 19193 29469 19227
rect 29469 19193 29503 19227
rect 29503 19193 29512 19227
rect 29460 19184 29512 19193
rect 23204 19116 23256 19168
rect 5915 19014 5967 19066
rect 5979 19014 6031 19066
rect 6043 19014 6095 19066
rect 6107 19014 6159 19066
rect 6171 19014 6223 19066
rect 15846 19014 15898 19066
rect 15910 19014 15962 19066
rect 15974 19014 16026 19066
rect 16038 19014 16090 19066
rect 16102 19014 16154 19066
rect 25776 19014 25828 19066
rect 25840 19014 25892 19066
rect 25904 19014 25956 19066
rect 25968 19014 26020 19066
rect 26032 19014 26084 19066
rect 31576 19048 31628 19100
rect 31760 19048 31812 19100
rect 1400 18912 1452 18964
rect 23204 18912 23256 18964
rect 29552 18912 29604 18964
rect 25412 18844 25464 18896
rect 26608 18844 26660 18896
rect 27528 18844 27580 18896
rect 28172 18844 28224 18896
rect 28448 18844 28500 18896
rect 19340 18776 19392 18828
rect 22468 18776 22520 18828
rect 27988 18776 28040 18828
rect 24584 18751 24636 18760
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 24860 18751 24912 18760
rect 24860 18717 24869 18751
rect 24869 18717 24903 18751
rect 24903 18717 24912 18751
rect 24860 18708 24912 18717
rect 28632 18751 28684 18760
rect 28632 18717 28641 18751
rect 28641 18717 28675 18751
rect 28675 18717 28684 18751
rect 28632 18708 28684 18717
rect 29000 18776 29052 18828
rect 1492 18640 1544 18692
rect 1400 18572 1452 18624
rect 25688 18640 25740 18692
rect 25964 18640 26016 18692
rect 28448 18640 28500 18692
rect 21732 18572 21784 18624
rect 23848 18572 23900 18624
rect 31760 18572 31812 18624
rect 10880 18470 10932 18522
rect 10944 18470 10996 18522
rect 11008 18470 11060 18522
rect 11072 18470 11124 18522
rect 11136 18470 11188 18522
rect 20811 18470 20863 18522
rect 20875 18470 20927 18522
rect 20939 18470 20991 18522
rect 21003 18470 21055 18522
rect 21067 18470 21119 18522
rect 22836 18368 22888 18420
rect 28356 18368 28408 18420
rect 31668 18368 31720 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 20720 18232 20772 18284
rect 22468 18300 22520 18352
rect 24124 18300 24176 18352
rect 27988 18300 28040 18352
rect 29368 18300 29420 18352
rect 22376 18232 22428 18284
rect 23848 18275 23900 18284
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 24032 18275 24084 18284
rect 24032 18241 24041 18275
rect 24041 18241 24075 18275
rect 24075 18241 24084 18275
rect 24032 18232 24084 18241
rect 24768 18275 24820 18284
rect 24768 18241 24777 18275
rect 24777 18241 24811 18275
rect 24811 18241 24820 18275
rect 24768 18232 24820 18241
rect 24860 18232 24912 18284
rect 28264 18275 28316 18284
rect 28264 18241 28273 18275
rect 28273 18241 28307 18275
rect 28307 18241 28316 18275
rect 28264 18232 28316 18241
rect 29000 18232 29052 18284
rect 23112 18164 23164 18216
rect 25136 18164 25188 18216
rect 1584 18139 1636 18148
rect 1584 18105 1593 18139
rect 1593 18105 1627 18139
rect 1627 18105 1636 18139
rect 1584 18096 1636 18105
rect 23848 18096 23900 18148
rect 25964 18164 26016 18216
rect 27344 18164 27396 18216
rect 31024 18164 31076 18216
rect 25412 18096 25464 18148
rect 29920 18096 29972 18148
rect 30288 18096 30340 18148
rect 1400 18028 1452 18080
rect 18788 18028 18840 18080
rect 19524 18028 19576 18080
rect 23664 18071 23716 18080
rect 23664 18037 23673 18071
rect 23673 18037 23707 18071
rect 23707 18037 23716 18071
rect 23664 18028 23716 18037
rect 24216 18028 24268 18080
rect 24584 18071 24636 18080
rect 24584 18037 24593 18071
rect 24593 18037 24627 18071
rect 24627 18037 24636 18071
rect 24584 18028 24636 18037
rect 25228 18028 25280 18080
rect 29368 18028 29420 18080
rect 29828 18028 29880 18080
rect 5915 17926 5967 17978
rect 5979 17926 6031 17978
rect 6043 17926 6095 17978
rect 6107 17926 6159 17978
rect 6171 17926 6223 17978
rect 15846 17926 15898 17978
rect 15910 17926 15962 17978
rect 15974 17926 16026 17978
rect 16038 17926 16090 17978
rect 16102 17926 16154 17978
rect 25776 17926 25828 17978
rect 25840 17926 25892 17978
rect 25904 17926 25956 17978
rect 25968 17926 26020 17978
rect 26032 17926 26084 17978
rect 22008 17824 22060 17876
rect 22744 17824 22796 17876
rect 23848 17867 23900 17876
rect 23848 17833 23857 17867
rect 23857 17833 23891 17867
rect 23891 17833 23900 17867
rect 23848 17824 23900 17833
rect 24032 17824 24084 17876
rect 25688 17867 25740 17876
rect 25688 17833 25697 17867
rect 25697 17833 25731 17867
rect 25731 17833 25740 17867
rect 25688 17824 25740 17833
rect 28632 17824 28684 17876
rect 29276 17756 29328 17808
rect 19432 17688 19484 17740
rect 26608 17688 26660 17740
rect 28632 17688 28684 17740
rect 30932 17688 30984 17740
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 20352 17620 20404 17672
rect 21456 17620 21508 17672
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 23664 17620 23716 17672
rect 25596 17620 25648 17672
rect 26056 17663 26108 17672
rect 26056 17629 26065 17663
rect 26065 17629 26099 17663
rect 26099 17629 26108 17663
rect 26056 17620 26108 17629
rect 26240 17620 26292 17672
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 28816 17620 28868 17672
rect 29920 17663 29972 17672
rect 29920 17629 29929 17663
rect 29929 17629 29963 17663
rect 29963 17629 29972 17663
rect 29920 17620 29972 17629
rect 18604 17552 18656 17604
rect 18972 17552 19024 17604
rect 22836 17552 22888 17604
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 19708 17484 19760 17536
rect 28908 17484 28960 17536
rect 10880 17382 10932 17434
rect 10944 17382 10996 17434
rect 11008 17382 11060 17434
rect 11072 17382 11124 17434
rect 11136 17382 11188 17434
rect 20811 17382 20863 17434
rect 20875 17382 20927 17434
rect 20939 17382 20991 17434
rect 21003 17382 21055 17434
rect 21067 17382 21119 17434
rect 18052 17280 18104 17332
rect 21548 17280 21600 17332
rect 22376 17280 22428 17332
rect 27528 17323 27580 17332
rect 27528 17289 27537 17323
rect 27537 17289 27571 17323
rect 27571 17289 27580 17323
rect 27528 17280 27580 17289
rect 27988 17280 28040 17332
rect 28724 17280 28776 17332
rect 29184 17323 29236 17332
rect 29184 17289 29193 17323
rect 29193 17289 29227 17323
rect 29227 17289 29236 17323
rect 29184 17280 29236 17289
rect 2688 17144 2740 17196
rect 17224 17144 17276 17196
rect 18604 17187 18656 17196
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 19524 17144 19576 17196
rect 23388 17212 23440 17264
rect 19892 17187 19944 17196
rect 19340 17076 19392 17128
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 20720 17144 20772 17196
rect 21272 17144 21324 17196
rect 24216 17144 24268 17196
rect 27436 17212 27488 17264
rect 28172 17212 28224 17264
rect 30012 17212 30064 17264
rect 20352 17076 20404 17128
rect 22836 17076 22888 17128
rect 24124 17076 24176 17128
rect 27068 17144 27120 17196
rect 28908 17144 28960 17196
rect 27712 17076 27764 17128
rect 29184 17076 29236 17128
rect 30104 17076 30156 17128
rect 18696 17008 18748 17060
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 17960 16940 18012 16992
rect 18512 16940 18564 16992
rect 19524 16940 19576 16992
rect 24032 16940 24084 16992
rect 25228 16940 25280 16992
rect 5915 16838 5967 16890
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 15846 16838 15898 16890
rect 15910 16838 15962 16890
rect 15974 16838 16026 16890
rect 16038 16838 16090 16890
rect 16102 16838 16154 16890
rect 25776 16838 25828 16890
rect 25840 16838 25892 16890
rect 25904 16838 25956 16890
rect 25968 16838 26020 16890
rect 26032 16838 26084 16890
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 18972 16736 19024 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 19892 16736 19944 16788
rect 27620 16779 27672 16788
rect 27620 16745 27629 16779
rect 27629 16745 27663 16779
rect 27663 16745 27672 16779
rect 27620 16736 27672 16745
rect 18696 16668 18748 16720
rect 18880 16668 18932 16720
rect 16488 16600 16540 16652
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 16212 16575 16264 16584
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 16856 16643 16908 16652
rect 16856 16609 16865 16643
rect 16865 16609 16899 16643
rect 16899 16609 16908 16643
rect 16856 16600 16908 16609
rect 18604 16532 18656 16584
rect 19432 16668 19484 16720
rect 19892 16643 19944 16652
rect 19892 16609 19901 16643
rect 19901 16609 19935 16643
rect 19935 16609 19944 16643
rect 19892 16600 19944 16609
rect 20444 16600 20496 16652
rect 26608 16600 26660 16652
rect 27528 16600 27580 16652
rect 28816 16600 28868 16652
rect 31300 16600 31352 16652
rect 19708 16575 19760 16584
rect 19708 16541 19743 16575
rect 19743 16541 19760 16575
rect 19708 16532 19760 16541
rect 2688 16464 2740 16516
rect 18696 16464 18748 16516
rect 18880 16464 18932 16516
rect 20076 16532 20128 16584
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 21180 16532 21232 16584
rect 28264 16532 28316 16584
rect 30104 16575 30156 16584
rect 30104 16541 30113 16575
rect 30113 16541 30147 16575
rect 30147 16541 30156 16575
rect 30104 16532 30156 16541
rect 16856 16396 16908 16448
rect 19340 16396 19392 16448
rect 25044 16464 25096 16516
rect 25504 16464 25556 16516
rect 27712 16464 27764 16516
rect 28724 16464 28776 16516
rect 19892 16396 19944 16448
rect 27344 16396 27396 16448
rect 27620 16396 27672 16448
rect 29828 16396 29880 16448
rect 10880 16294 10932 16346
rect 10944 16294 10996 16346
rect 11008 16294 11060 16346
rect 11072 16294 11124 16346
rect 11136 16294 11188 16346
rect 20811 16294 20863 16346
rect 20875 16294 20927 16346
rect 20939 16294 20991 16346
rect 21003 16294 21055 16346
rect 21067 16294 21119 16346
rect 18236 16192 18288 16244
rect 18420 16192 18472 16244
rect 28356 16192 28408 16244
rect 31116 16192 31168 16244
rect 16948 16124 17000 16176
rect 17684 16124 17736 16176
rect 17776 16124 17828 16176
rect 17914 16124 17966 16176
rect 26240 16124 26292 16176
rect 27068 16124 27120 16176
rect 27344 16124 27396 16176
rect 27620 16124 27672 16176
rect 28724 16167 28776 16176
rect 28724 16133 28733 16167
rect 28733 16133 28767 16167
rect 28767 16133 28776 16167
rect 28724 16124 28776 16133
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 19340 16056 19392 16108
rect 18328 15988 18380 16040
rect 21824 16099 21876 16108
rect 21824 16065 21833 16099
rect 21833 16065 21867 16099
rect 21867 16065 21876 16099
rect 21824 16056 21876 16065
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 25228 16099 25280 16108
rect 25228 16065 25237 16099
rect 25237 16065 25271 16099
rect 25271 16065 25280 16099
rect 25228 16056 25280 16065
rect 25596 16056 25648 16108
rect 28448 16099 28500 16108
rect 28448 16065 28457 16099
rect 28457 16065 28491 16099
rect 28491 16065 28500 16099
rect 28448 16056 28500 16065
rect 29920 16099 29972 16108
rect 29920 16065 29929 16099
rect 29929 16065 29963 16099
rect 29963 16065 29972 16099
rect 29920 16056 29972 16065
rect 20352 15988 20404 16040
rect 27436 15988 27488 16040
rect 18604 15920 18656 15972
rect 21916 15920 21968 15972
rect 26148 15920 26200 15972
rect 1400 15852 1452 15904
rect 1768 15852 1820 15904
rect 16672 15852 16724 15904
rect 18052 15852 18104 15904
rect 19708 15852 19760 15904
rect 27988 15852 28040 15904
rect 28448 15852 28500 15904
rect 5915 15750 5967 15802
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 15846 15750 15898 15802
rect 15910 15750 15962 15802
rect 15974 15750 16026 15802
rect 16038 15750 16090 15802
rect 16102 15750 16154 15802
rect 25776 15750 25828 15802
rect 25840 15750 25892 15802
rect 25904 15750 25956 15802
rect 25968 15750 26020 15802
rect 26032 15750 26084 15802
rect 1768 15444 1820 15496
rect 16672 15648 16724 15700
rect 16948 15648 17000 15700
rect 28264 15648 28316 15700
rect 19340 15580 19392 15632
rect 20352 15580 20404 15632
rect 29000 15580 29052 15632
rect 20536 15512 20588 15564
rect 21640 15512 21692 15564
rect 21916 15512 21968 15564
rect 26608 15512 26660 15564
rect 26884 15512 26936 15564
rect 27712 15555 27764 15564
rect 27712 15521 27721 15555
rect 27721 15521 27755 15555
rect 27755 15521 27764 15555
rect 27712 15512 27764 15521
rect 16580 15444 16632 15496
rect 19248 15444 19300 15496
rect 19708 15487 19760 15496
rect 18420 15376 18472 15428
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 20168 15487 20220 15496
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 20444 15487 20496 15496
rect 20444 15453 20453 15487
rect 20453 15453 20487 15487
rect 20487 15453 20496 15487
rect 20444 15444 20496 15453
rect 21548 15487 21600 15496
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 24492 15444 24544 15496
rect 25596 15487 25648 15496
rect 25596 15453 25605 15487
rect 25605 15453 25639 15487
rect 25639 15453 25648 15487
rect 25596 15444 25648 15453
rect 26148 15444 26200 15496
rect 26240 15444 26292 15496
rect 27436 15487 27488 15496
rect 27436 15453 27445 15487
rect 27445 15453 27479 15487
rect 27479 15453 27488 15487
rect 27436 15444 27488 15453
rect 29000 15487 29052 15496
rect 29000 15453 29009 15487
rect 29009 15453 29043 15487
rect 29043 15453 29052 15487
rect 29000 15444 29052 15453
rect 20628 15376 20680 15428
rect 24216 15376 24268 15428
rect 24676 15376 24728 15428
rect 25412 15419 25464 15428
rect 25412 15385 25421 15419
rect 25421 15385 25455 15419
rect 25455 15385 25464 15419
rect 25412 15376 25464 15385
rect 26884 15376 26936 15428
rect 27620 15419 27672 15428
rect 27620 15385 27629 15419
rect 27629 15385 27663 15419
rect 27663 15385 27672 15419
rect 27620 15376 27672 15385
rect 29920 15419 29972 15428
rect 29920 15385 29929 15419
rect 29929 15385 29963 15419
rect 29963 15385 29972 15419
rect 29920 15376 29972 15385
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 2136 15351 2188 15360
rect 2136 15317 2145 15351
rect 2145 15317 2179 15351
rect 2179 15317 2188 15351
rect 2136 15308 2188 15317
rect 27528 15308 27580 15360
rect 10880 15206 10932 15258
rect 10944 15206 10996 15258
rect 11008 15206 11060 15258
rect 11072 15206 11124 15258
rect 11136 15206 11188 15258
rect 20811 15206 20863 15258
rect 20875 15206 20927 15258
rect 20939 15206 20991 15258
rect 21003 15206 21055 15258
rect 21067 15206 21119 15258
rect 19800 15036 19852 15088
rect 20352 15036 20404 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 20720 14968 20772 15020
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 21180 15011 21232 15020
rect 21180 14977 21189 15011
rect 21189 14977 21223 15011
rect 21223 14977 21232 15011
rect 21180 14968 21232 14977
rect 19432 14900 19484 14952
rect 20076 14900 20128 14952
rect 21548 14900 21600 14952
rect 22468 15104 22520 15156
rect 23480 15104 23532 15156
rect 25412 15104 25464 15156
rect 25228 15036 25280 15088
rect 22468 14968 22520 15020
rect 23756 14968 23808 15020
rect 24032 14968 24084 15020
rect 23204 14900 23256 14952
rect 25412 14968 25464 15020
rect 27436 15104 27488 15156
rect 28264 15147 28316 15156
rect 27620 15036 27672 15088
rect 28264 15113 28273 15147
rect 28273 15113 28307 15147
rect 28307 15113 28316 15147
rect 28264 15104 28316 15113
rect 27068 14968 27120 15020
rect 27988 14968 28040 15020
rect 28080 14968 28132 15020
rect 27528 14900 27580 14952
rect 28908 14900 28960 14952
rect 17224 14832 17276 14884
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 19984 14764 20036 14816
rect 23388 14764 23440 14816
rect 24032 14764 24084 14816
rect 25044 14807 25096 14816
rect 25044 14773 25053 14807
rect 25053 14773 25087 14807
rect 25087 14773 25096 14807
rect 25044 14764 25096 14773
rect 25412 14764 25464 14816
rect 26332 14764 26384 14816
rect 27436 14764 27488 14816
rect 5915 14662 5967 14714
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 15846 14662 15898 14714
rect 15910 14662 15962 14714
rect 15974 14662 16026 14714
rect 16038 14662 16090 14714
rect 16102 14662 16154 14714
rect 25776 14662 25828 14714
rect 25840 14662 25892 14714
rect 25904 14662 25956 14714
rect 25968 14662 26020 14714
rect 26032 14662 26084 14714
rect 1400 14560 1452 14612
rect 17224 14560 17276 14612
rect 18420 14560 18472 14612
rect 20076 14560 20128 14612
rect 21824 14560 21876 14612
rect 22468 14603 22520 14612
rect 22468 14569 22477 14603
rect 22477 14569 22511 14603
rect 22511 14569 22520 14603
rect 22468 14560 22520 14569
rect 24860 14560 24912 14612
rect 25412 14560 25464 14612
rect 6276 14492 6328 14544
rect 19524 14492 19576 14544
rect 2136 14356 2188 14408
rect 19432 14356 19484 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 20260 14424 20312 14476
rect 19984 14356 20036 14408
rect 20168 14356 20220 14408
rect 20904 14424 20956 14476
rect 23480 14424 23532 14476
rect 20628 14399 20680 14408
rect 20628 14365 20637 14399
rect 20637 14365 20671 14399
rect 20671 14365 20680 14399
rect 20628 14356 20680 14365
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 19524 14220 19576 14272
rect 20444 14288 20496 14340
rect 23112 14356 23164 14408
rect 25320 14356 25372 14408
rect 26148 14399 26200 14408
rect 26148 14365 26157 14399
rect 26157 14365 26191 14399
rect 26191 14365 26200 14399
rect 26148 14356 26200 14365
rect 27068 14535 27120 14544
rect 27068 14501 27077 14535
rect 27077 14501 27111 14535
rect 27111 14501 27120 14535
rect 27068 14492 27120 14501
rect 30840 14560 30892 14612
rect 27344 14492 27396 14544
rect 27528 14424 27580 14476
rect 27988 14492 28040 14544
rect 28264 14424 28316 14476
rect 30104 14424 30156 14476
rect 27804 14356 27856 14408
rect 29828 14399 29880 14408
rect 29828 14365 29837 14399
rect 29837 14365 29871 14399
rect 29871 14365 29880 14399
rect 29828 14356 29880 14365
rect 24400 14288 24452 14340
rect 24860 14288 24912 14340
rect 25780 14220 25832 14272
rect 28724 14288 28776 14340
rect 26792 14220 26844 14272
rect 28816 14263 28868 14272
rect 28816 14229 28825 14263
rect 28825 14229 28859 14263
rect 28859 14229 28868 14263
rect 28816 14220 28868 14229
rect 10880 14118 10932 14170
rect 10944 14118 10996 14170
rect 11008 14118 11060 14170
rect 11072 14118 11124 14170
rect 11136 14118 11188 14170
rect 20811 14118 20863 14170
rect 20875 14118 20927 14170
rect 20939 14118 20991 14170
rect 21003 14118 21055 14170
rect 21067 14118 21119 14170
rect 20536 14016 20588 14068
rect 28080 14016 28132 14068
rect 21824 13991 21876 14000
rect 21824 13957 21833 13991
rect 21833 13957 21867 13991
rect 21867 13957 21876 13991
rect 21824 13948 21876 13957
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 23388 13880 23440 13932
rect 24124 13880 24176 13932
rect 26240 13948 26292 14000
rect 27436 13991 27488 14000
rect 27436 13957 27445 13991
rect 27445 13957 27479 13991
rect 27479 13957 27488 13991
rect 27436 13948 27488 13957
rect 28540 13948 28592 14000
rect 28632 13991 28684 14000
rect 28632 13957 28641 13991
rect 28641 13957 28675 13991
rect 28675 13957 28684 13991
rect 28632 13948 28684 13957
rect 25228 13880 25280 13932
rect 25504 13880 25556 13932
rect 24584 13812 24636 13864
rect 26148 13812 26200 13864
rect 28724 13855 28776 13864
rect 28724 13821 28733 13855
rect 28733 13821 28767 13855
rect 28767 13821 28776 13855
rect 28724 13812 28776 13821
rect 28908 13812 28960 13864
rect 22376 13744 22428 13796
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 22192 13719 22244 13728
rect 22192 13685 22201 13719
rect 22201 13685 22235 13719
rect 22235 13685 22244 13719
rect 22192 13676 22244 13685
rect 23756 13719 23808 13728
rect 23756 13685 23765 13719
rect 23765 13685 23799 13719
rect 23799 13685 23808 13719
rect 23756 13676 23808 13685
rect 26240 13744 26292 13796
rect 27712 13744 27764 13796
rect 5915 13574 5967 13626
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 15846 13574 15898 13626
rect 15910 13574 15962 13626
rect 15974 13574 16026 13626
rect 16038 13574 16090 13626
rect 16102 13574 16154 13626
rect 25776 13574 25828 13626
rect 25840 13574 25892 13626
rect 25904 13574 25956 13626
rect 25968 13574 26020 13626
rect 26032 13574 26084 13626
rect 20352 13336 20404 13388
rect 20536 13268 20588 13320
rect 22192 13472 22244 13524
rect 23204 13515 23256 13524
rect 23204 13481 23213 13515
rect 23213 13481 23247 13515
rect 23247 13481 23256 13515
rect 23204 13472 23256 13481
rect 24400 13515 24452 13524
rect 24400 13481 24409 13515
rect 24409 13481 24443 13515
rect 24443 13481 24452 13515
rect 24400 13472 24452 13481
rect 26608 13472 26660 13524
rect 27436 13472 27488 13524
rect 22928 13404 22980 13456
rect 24124 13336 24176 13388
rect 20628 13200 20680 13252
rect 21272 13268 21324 13320
rect 21548 13268 21600 13320
rect 23204 13268 23256 13320
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 25136 13336 25188 13388
rect 26240 13336 26292 13388
rect 26700 13336 26752 13388
rect 28724 13472 28776 13524
rect 25412 13268 25464 13320
rect 26148 13268 26200 13320
rect 26792 13268 26844 13320
rect 31392 13404 31444 13456
rect 28724 13336 28776 13388
rect 22652 13200 22704 13252
rect 26240 13243 26292 13252
rect 26240 13209 26249 13243
rect 26249 13209 26283 13243
rect 26283 13209 26292 13243
rect 26240 13200 26292 13209
rect 26700 13200 26752 13252
rect 30012 13268 30064 13320
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 19340 13132 19392 13184
rect 19524 13132 19576 13184
rect 21364 13175 21416 13184
rect 21364 13141 21373 13175
rect 21373 13141 21407 13175
rect 21407 13141 21416 13175
rect 21364 13132 21416 13141
rect 24216 13132 24268 13184
rect 25504 13132 25556 13184
rect 28172 13200 28224 13252
rect 27068 13175 27120 13184
rect 27068 13141 27077 13175
rect 27077 13141 27111 13175
rect 27111 13141 27120 13175
rect 27068 13132 27120 13141
rect 27436 13132 27488 13184
rect 10880 13030 10932 13082
rect 10944 13030 10996 13082
rect 11008 13030 11060 13082
rect 11072 13030 11124 13082
rect 11136 13030 11188 13082
rect 20811 13030 20863 13082
rect 20875 13030 20927 13082
rect 20939 13030 20991 13082
rect 21003 13030 21055 13082
rect 21067 13030 21119 13082
rect 20628 12971 20680 12980
rect 20628 12937 20637 12971
rect 20637 12937 20671 12971
rect 20671 12937 20680 12971
rect 20628 12928 20680 12937
rect 22100 12928 22152 12980
rect 22284 12928 22336 12980
rect 22652 12928 22704 12980
rect 24860 12928 24912 12980
rect 25412 12928 25464 12980
rect 26332 12928 26384 12980
rect 27252 12928 27304 12980
rect 28264 12928 28316 12980
rect 28356 12928 28408 12980
rect 2044 12860 2096 12912
rect 28448 12903 28500 12912
rect 28448 12869 28457 12903
rect 28457 12869 28491 12903
rect 28491 12869 28500 12903
rect 28448 12860 28500 12869
rect 28724 12903 28776 12912
rect 28724 12869 28733 12903
rect 28733 12869 28767 12903
rect 28767 12869 28776 12903
rect 28724 12860 28776 12869
rect 20628 12792 20680 12844
rect 23756 12792 23808 12844
rect 24860 12835 24912 12844
rect 24860 12801 24869 12835
rect 24869 12801 24903 12835
rect 24903 12801 24912 12835
rect 24860 12792 24912 12801
rect 25412 12792 25464 12844
rect 25504 12792 25556 12844
rect 26332 12792 26384 12844
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 20812 12724 20864 12776
rect 21272 12724 21324 12776
rect 23112 12767 23164 12776
rect 23112 12733 23121 12767
rect 23121 12733 23155 12767
rect 23155 12733 23164 12767
rect 23112 12724 23164 12733
rect 23204 12767 23256 12776
rect 23204 12733 23213 12767
rect 23213 12733 23247 12767
rect 23247 12733 23256 12767
rect 23204 12724 23256 12733
rect 23388 12724 23440 12776
rect 29368 12724 29420 12776
rect 29552 12767 29604 12776
rect 29552 12733 29561 12767
rect 29561 12733 29595 12767
rect 29595 12733 29604 12767
rect 29552 12724 29604 12733
rect 2320 12656 2372 12708
rect 25044 12631 25096 12640
rect 25044 12597 25053 12631
rect 25053 12597 25087 12631
rect 25087 12597 25096 12631
rect 25044 12588 25096 12597
rect 5915 12486 5967 12538
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 15846 12486 15898 12538
rect 15910 12486 15962 12538
rect 15974 12486 16026 12538
rect 16038 12486 16090 12538
rect 16102 12486 16154 12538
rect 25776 12486 25828 12538
rect 25840 12486 25892 12538
rect 25904 12486 25956 12538
rect 25968 12486 26020 12538
rect 26032 12486 26084 12538
rect 2044 12427 2096 12436
rect 2044 12393 2053 12427
rect 2053 12393 2087 12427
rect 2087 12393 2096 12427
rect 2044 12384 2096 12393
rect 26424 12384 26476 12436
rect 27436 12384 27488 12436
rect 26792 12316 26844 12368
rect 20352 12248 20404 12300
rect 27528 12291 27580 12300
rect 2044 12180 2096 12232
rect 2688 12180 2740 12232
rect 6276 12180 6328 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 18512 12180 18564 12232
rect 20720 12223 20772 12232
rect 20720 12189 20729 12223
rect 20729 12189 20763 12223
rect 20763 12189 20772 12223
rect 20720 12180 20772 12189
rect 27528 12257 27537 12291
rect 27537 12257 27571 12291
rect 27571 12257 27580 12291
rect 27528 12248 27580 12257
rect 21916 12180 21968 12232
rect 23572 12180 23624 12232
rect 26148 12180 26200 12232
rect 28172 12223 28224 12232
rect 28172 12189 28181 12223
rect 28181 12189 28215 12223
rect 28215 12189 28224 12223
rect 28172 12180 28224 12189
rect 22836 12112 22888 12164
rect 24676 12112 24728 12164
rect 25964 12112 26016 12164
rect 29644 12112 29696 12164
rect 29920 12155 29972 12164
rect 29920 12121 29929 12155
rect 29929 12121 29963 12155
rect 29963 12121 29972 12155
rect 29920 12112 29972 12121
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 17500 12087 17552 12096
rect 17500 12053 17509 12087
rect 17509 12053 17543 12087
rect 17543 12053 17552 12087
rect 17500 12044 17552 12053
rect 17868 12044 17920 12096
rect 20352 12044 20404 12096
rect 25044 12044 25096 12096
rect 25872 12044 25924 12096
rect 26884 12044 26936 12096
rect 10880 11942 10932 11994
rect 10944 11942 10996 11994
rect 11008 11942 11060 11994
rect 11072 11942 11124 11994
rect 11136 11942 11188 11994
rect 20811 11942 20863 11994
rect 20875 11942 20927 11994
rect 20939 11942 20991 11994
rect 21003 11942 21055 11994
rect 21067 11942 21119 11994
rect 19340 11840 19392 11892
rect 19984 11840 20036 11892
rect 20628 11840 20680 11892
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 26240 11840 26292 11892
rect 27620 11840 27672 11892
rect 27804 11840 27856 11892
rect 4804 11772 4856 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 17868 11747 17920 11756
rect 17868 11713 17877 11747
rect 17877 11713 17911 11747
rect 17911 11713 17920 11747
rect 17868 11704 17920 11713
rect 19248 11704 19300 11756
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 19616 11636 19668 11688
rect 19800 11636 19852 11688
rect 20260 11704 20312 11756
rect 21364 11704 21416 11756
rect 29736 11772 29788 11824
rect 24860 11747 24912 11756
rect 24860 11713 24869 11747
rect 24869 11713 24903 11747
rect 24903 11713 24912 11747
rect 24860 11704 24912 11713
rect 25964 11704 26016 11756
rect 28816 11747 28868 11756
rect 25044 11679 25096 11688
rect 25044 11645 25053 11679
rect 25053 11645 25087 11679
rect 25087 11645 25096 11679
rect 25044 11636 25096 11645
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 19708 11543 19760 11552
rect 19708 11509 19717 11543
rect 19717 11509 19751 11543
rect 19751 11509 19760 11543
rect 19708 11500 19760 11509
rect 23204 11500 23256 11552
rect 25412 11636 25464 11688
rect 28816 11713 28825 11747
rect 28825 11713 28859 11747
rect 28859 11713 28868 11747
rect 28816 11704 28868 11713
rect 29460 11704 29512 11756
rect 29276 11679 29328 11688
rect 25872 11568 25924 11620
rect 25504 11500 25556 11552
rect 26700 11568 26752 11620
rect 26608 11500 26660 11552
rect 27528 11568 27580 11620
rect 29276 11645 29285 11679
rect 29285 11645 29319 11679
rect 29319 11645 29328 11679
rect 29276 11636 29328 11645
rect 5915 11398 5967 11450
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 15846 11398 15898 11450
rect 15910 11398 15962 11450
rect 15974 11398 16026 11450
rect 16038 11398 16090 11450
rect 16102 11398 16154 11450
rect 25776 11398 25828 11450
rect 25840 11398 25892 11450
rect 25904 11398 25956 11450
rect 25968 11398 26020 11450
rect 26032 11398 26084 11450
rect 1400 11296 1452 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 21180 11296 21232 11348
rect 21364 11296 21416 11348
rect 27528 11296 27580 11348
rect 28448 11296 28500 11348
rect 30104 11296 30156 11348
rect 19616 11228 19668 11280
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 19432 11092 19484 11144
rect 20168 11160 20220 11212
rect 20260 11160 20312 11212
rect 21640 11160 21692 11212
rect 20352 11092 20404 11144
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 19800 11024 19852 11076
rect 20628 11092 20680 11144
rect 23204 11092 23256 11144
rect 24032 11092 24084 11144
rect 24400 11092 24452 11144
rect 25136 11160 25188 11212
rect 27160 11160 27212 11212
rect 27436 11160 27488 11212
rect 21180 11024 21232 11076
rect 21456 11024 21508 11076
rect 22836 11024 22888 11076
rect 23020 11024 23072 11076
rect 25320 11092 25372 11144
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 28264 11092 28316 11144
rect 28724 11135 28776 11144
rect 28724 11101 28733 11135
rect 28733 11101 28767 11135
rect 28767 11101 28776 11135
rect 28724 11092 28776 11101
rect 28908 11092 28960 11144
rect 25412 11024 25464 11076
rect 25688 11024 25740 11076
rect 26240 11024 26292 11076
rect 24216 10956 24268 11008
rect 24400 10999 24452 11008
rect 24400 10965 24409 10999
rect 24409 10965 24443 10999
rect 24443 10965 24452 10999
rect 24400 10956 24452 10965
rect 10880 10854 10932 10906
rect 10944 10854 10996 10906
rect 11008 10854 11060 10906
rect 11072 10854 11124 10906
rect 11136 10854 11188 10906
rect 20811 10854 20863 10906
rect 20875 10854 20927 10906
rect 20939 10854 20991 10906
rect 21003 10854 21055 10906
rect 21067 10854 21119 10906
rect 20352 10752 20404 10804
rect 23204 10795 23256 10804
rect 23204 10761 23213 10795
rect 23213 10761 23247 10795
rect 23247 10761 23256 10795
rect 23204 10752 23256 10761
rect 17960 10684 18012 10736
rect 19708 10684 19760 10736
rect 17500 10616 17552 10668
rect 19432 10616 19484 10668
rect 20444 10684 20496 10736
rect 20536 10616 20588 10668
rect 22652 10616 22704 10668
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 25136 10752 25188 10804
rect 24216 10684 24268 10736
rect 28080 10795 28132 10804
rect 28080 10761 28089 10795
rect 28089 10761 28123 10795
rect 28123 10761 28132 10795
rect 28080 10752 28132 10761
rect 29368 10795 29420 10804
rect 29368 10761 29377 10795
rect 29377 10761 29411 10795
rect 29411 10761 29420 10795
rect 29368 10752 29420 10761
rect 30656 10752 30708 10804
rect 27620 10684 27672 10736
rect 19340 10548 19392 10600
rect 21548 10548 21600 10600
rect 26792 10616 26844 10668
rect 27528 10548 27580 10600
rect 26884 10480 26936 10532
rect 27252 10480 27304 10532
rect 29184 10548 29236 10600
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 21456 10412 21508 10464
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 5915 10310 5967 10362
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 15846 10310 15898 10362
rect 15910 10310 15962 10362
rect 15974 10310 16026 10362
rect 16038 10310 16090 10362
rect 16102 10310 16154 10362
rect 25776 10310 25828 10362
rect 25840 10310 25892 10362
rect 25904 10310 25956 10362
rect 25968 10310 26020 10362
rect 26032 10310 26084 10362
rect 21916 10251 21968 10260
rect 21916 10217 21925 10251
rect 21925 10217 21959 10251
rect 21959 10217 21968 10251
rect 21916 10208 21968 10217
rect 22652 10208 22704 10260
rect 23112 10251 23164 10260
rect 23112 10217 23121 10251
rect 23121 10217 23155 10251
rect 23155 10217 23164 10251
rect 23112 10208 23164 10217
rect 26332 10251 26384 10260
rect 26332 10217 26341 10251
rect 26341 10217 26375 10251
rect 26375 10217 26384 10251
rect 26332 10208 26384 10217
rect 17960 10140 18012 10192
rect 20536 10072 20588 10124
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 21640 10072 21692 10124
rect 2136 10004 2188 10056
rect 2688 10004 2740 10056
rect 20352 10004 20404 10056
rect 21180 10047 21232 10056
rect 21180 10013 21189 10047
rect 21189 10013 21223 10047
rect 21223 10013 21232 10047
rect 21180 10004 21232 10013
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 24400 10072 24452 10124
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 27068 10004 27120 10056
rect 28264 10004 28316 10056
rect 25504 9936 25556 9988
rect 26240 9979 26292 9988
rect 26240 9945 26249 9979
rect 26249 9945 26283 9979
rect 26283 9945 26292 9979
rect 29736 9979 29788 9988
rect 26240 9936 26292 9945
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2136 9911 2188 9920
rect 2136 9877 2145 9911
rect 2145 9877 2179 9911
rect 2179 9877 2188 9911
rect 2136 9868 2188 9877
rect 28816 9911 28868 9920
rect 28816 9877 28825 9911
rect 28825 9877 28859 9911
rect 28859 9877 28868 9911
rect 28816 9868 28868 9877
rect 29736 9945 29745 9979
rect 29745 9945 29779 9979
rect 29779 9945 29788 9979
rect 29736 9936 29788 9945
rect 10880 9766 10932 9818
rect 10944 9766 10996 9818
rect 11008 9766 11060 9818
rect 11072 9766 11124 9818
rect 11136 9766 11188 9818
rect 20811 9766 20863 9818
rect 20875 9766 20927 9818
rect 20939 9766 20991 9818
rect 21003 9766 21055 9818
rect 21067 9766 21119 9818
rect 20352 9664 20404 9716
rect 7564 9596 7616 9648
rect 2320 9392 2372 9444
rect 20628 9596 20680 9648
rect 21364 9664 21416 9716
rect 24032 9664 24084 9716
rect 20168 9571 20220 9580
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 20444 9571 20496 9580
rect 20444 9537 20453 9571
rect 20453 9537 20487 9571
rect 20487 9537 20496 9571
rect 30380 9596 30432 9648
rect 31852 9596 31904 9648
rect 20444 9528 20496 9537
rect 23848 9528 23900 9580
rect 25596 9528 25648 9580
rect 27068 9571 27120 9580
rect 27068 9537 27077 9571
rect 27077 9537 27111 9571
rect 27111 9537 27120 9571
rect 27068 9528 27120 9537
rect 20536 9460 20588 9512
rect 23296 9460 23348 9512
rect 26700 9460 26752 9512
rect 27436 9528 27488 9580
rect 28632 9528 28684 9580
rect 29184 9460 29236 9512
rect 22376 9324 22428 9376
rect 22652 9367 22704 9376
rect 22652 9333 22661 9367
rect 22661 9333 22695 9367
rect 22695 9333 22704 9367
rect 22652 9324 22704 9333
rect 23112 9324 23164 9376
rect 25320 9324 25372 9376
rect 5915 9222 5967 9274
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 15846 9222 15898 9274
rect 15910 9222 15962 9274
rect 15974 9222 16026 9274
rect 16038 9222 16090 9274
rect 16102 9222 16154 9274
rect 25776 9222 25828 9274
rect 25840 9222 25892 9274
rect 25904 9222 25956 9274
rect 25968 9222 26020 9274
rect 26032 9222 26084 9274
rect 2688 9120 2740 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 20444 9052 20496 9104
rect 22836 9120 22888 9172
rect 23296 9120 23348 9172
rect 30012 9163 30064 9172
rect 30012 9129 30021 9163
rect 30021 9129 30055 9163
rect 30055 9129 30064 9163
rect 30012 9120 30064 9129
rect 28724 9052 28776 9104
rect 24584 8984 24636 9036
rect 28816 9027 28868 9036
rect 28816 8993 28825 9027
rect 28825 8993 28859 9027
rect 28859 8993 28868 9027
rect 28816 8984 28868 8993
rect 2136 8916 2188 8968
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 20536 8916 20588 8968
rect 21548 8959 21600 8968
rect 21548 8925 21557 8959
rect 21557 8925 21591 8959
rect 21591 8925 21600 8959
rect 21548 8916 21600 8925
rect 22652 8916 22704 8968
rect 25320 8916 25372 8968
rect 27436 8916 27488 8968
rect 28632 8959 28684 8968
rect 28632 8925 28641 8959
rect 28641 8925 28675 8959
rect 28675 8925 28684 8959
rect 28632 8916 28684 8925
rect 29828 8959 29880 8968
rect 29828 8925 29837 8959
rect 29837 8925 29871 8959
rect 29871 8925 29880 8959
rect 29828 8916 29880 8925
rect 20168 8848 20220 8900
rect 26148 8848 26200 8900
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2136 8823 2188 8832
rect 2136 8789 2145 8823
rect 2145 8789 2179 8823
rect 2179 8789 2188 8823
rect 2136 8780 2188 8789
rect 23112 8780 23164 8832
rect 27252 8780 27304 8832
rect 28264 8823 28316 8832
rect 28264 8789 28273 8823
rect 28273 8789 28307 8823
rect 28307 8789 28316 8823
rect 28264 8780 28316 8789
rect 30380 8848 30432 8900
rect 29368 8780 29420 8832
rect 10880 8678 10932 8730
rect 10944 8678 10996 8730
rect 11008 8678 11060 8730
rect 11072 8678 11124 8730
rect 11136 8678 11188 8730
rect 20811 8678 20863 8730
rect 20875 8678 20927 8730
rect 20939 8678 20991 8730
rect 21003 8678 21055 8730
rect 21067 8678 21119 8730
rect 2136 8440 2188 8492
rect 24032 8440 24084 8492
rect 24584 8440 24636 8492
rect 25596 8508 25648 8560
rect 26148 8576 26200 8628
rect 27068 8576 27120 8628
rect 29368 8576 29420 8628
rect 30748 8576 30800 8628
rect 26516 8508 26568 8560
rect 26608 8508 26660 8560
rect 24768 8440 24820 8492
rect 25044 8440 25096 8492
rect 27068 8440 27120 8492
rect 27528 8440 27580 8492
rect 29276 8440 29328 8492
rect 25596 8372 25648 8424
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 1584 8304 1636 8313
rect 14280 8304 14332 8356
rect 29184 8372 29236 8424
rect 26424 8304 26476 8356
rect 24032 8279 24084 8288
rect 24032 8245 24041 8279
rect 24041 8245 24075 8279
rect 24075 8245 24084 8279
rect 24032 8236 24084 8245
rect 27344 8279 27396 8288
rect 27344 8245 27353 8279
rect 27353 8245 27387 8279
rect 27387 8245 27396 8279
rect 27344 8236 27396 8245
rect 27896 8236 27948 8288
rect 5915 8134 5967 8186
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 15846 8134 15898 8186
rect 15910 8134 15962 8186
rect 15974 8134 16026 8186
rect 16038 8134 16090 8186
rect 16102 8134 16154 8186
rect 25776 8134 25828 8186
rect 25840 8134 25892 8186
rect 25904 8134 25956 8186
rect 25968 8134 26020 8186
rect 26032 8134 26084 8186
rect 23112 8032 23164 8084
rect 27068 7964 27120 8016
rect 2688 7828 2740 7880
rect 24032 7896 24084 7948
rect 25504 7939 25556 7948
rect 25504 7905 25513 7939
rect 25513 7905 25547 7939
rect 25547 7905 25556 7939
rect 25504 7896 25556 7905
rect 23388 7828 23440 7880
rect 25688 7828 25740 7880
rect 26056 7828 26108 7880
rect 28264 7871 28316 7880
rect 28264 7837 28273 7871
rect 28273 7837 28307 7871
rect 28307 7837 28316 7871
rect 28264 7828 28316 7837
rect 28724 7828 28776 7880
rect 25964 7760 26016 7812
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 22652 7735 22704 7744
rect 22652 7701 22661 7735
rect 22661 7701 22695 7735
rect 22695 7701 22704 7735
rect 22652 7692 22704 7701
rect 25228 7692 25280 7744
rect 26148 7692 26200 7744
rect 28356 7735 28408 7744
rect 28356 7701 28365 7735
rect 28365 7701 28399 7735
rect 28399 7701 28408 7735
rect 28356 7692 28408 7701
rect 10880 7590 10932 7642
rect 10944 7590 10996 7642
rect 11008 7590 11060 7642
rect 11072 7590 11124 7642
rect 11136 7590 11188 7642
rect 20811 7590 20863 7642
rect 20875 7590 20927 7642
rect 20939 7590 20991 7642
rect 21003 7590 21055 7642
rect 21067 7590 21119 7642
rect 2044 7488 2096 7540
rect 28356 7488 28408 7540
rect 29092 7531 29144 7540
rect 29092 7497 29101 7531
rect 29101 7497 29135 7531
rect 29135 7497 29144 7531
rect 29092 7488 29144 7497
rect 30472 7488 30524 7540
rect 6368 7420 6420 7472
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 25688 7352 25740 7404
rect 26976 7395 27028 7404
rect 26976 7361 26985 7395
rect 26985 7361 27019 7395
rect 27019 7361 27028 7395
rect 26976 7352 27028 7361
rect 29000 7352 29052 7404
rect 25412 7284 25464 7336
rect 25504 7284 25556 7336
rect 26056 7327 26108 7336
rect 26056 7293 26065 7327
rect 26065 7293 26099 7327
rect 26099 7293 26108 7327
rect 26056 7284 26108 7293
rect 25964 7216 26016 7268
rect 26792 7284 26844 7336
rect 29184 7284 29236 7336
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 25228 7148 25280 7200
rect 26148 7148 26200 7200
rect 5915 7046 5967 7098
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 15846 7046 15898 7098
rect 15910 7046 15962 7098
rect 15974 7046 16026 7098
rect 16038 7046 16090 7098
rect 16102 7046 16154 7098
rect 25776 7046 25828 7098
rect 25840 7046 25892 7098
rect 25904 7046 25956 7098
rect 25968 7046 26020 7098
rect 26032 7046 26084 7098
rect 23388 6944 23440 6996
rect 28540 6944 28592 6996
rect 25596 6876 25648 6928
rect 26148 6876 26200 6928
rect 26976 6876 27028 6928
rect 25412 6851 25464 6860
rect 25412 6817 25421 6851
rect 25421 6817 25455 6851
rect 25455 6817 25464 6851
rect 25412 6808 25464 6817
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 25504 6740 25556 6792
rect 22008 6672 22060 6724
rect 27712 6808 27764 6860
rect 28724 6851 28776 6860
rect 28724 6817 28733 6851
rect 28733 6817 28767 6851
rect 28767 6817 28776 6851
rect 28724 6808 28776 6817
rect 27620 6783 27672 6792
rect 27620 6749 27629 6783
rect 27629 6749 27663 6783
rect 27663 6749 27672 6783
rect 27620 6740 27672 6749
rect 30196 6808 30248 6860
rect 28908 6740 28960 6792
rect 29000 6672 29052 6724
rect 22652 6604 22704 6656
rect 25688 6604 25740 6656
rect 27252 6604 27304 6656
rect 27436 6647 27488 6656
rect 27436 6613 27445 6647
rect 27445 6613 27479 6647
rect 27479 6613 27488 6647
rect 27436 6604 27488 6613
rect 28080 6647 28132 6656
rect 28080 6613 28089 6647
rect 28089 6613 28123 6647
rect 28123 6613 28132 6647
rect 28080 6604 28132 6613
rect 29092 6604 29144 6656
rect 10880 6502 10932 6554
rect 10944 6502 10996 6554
rect 11008 6502 11060 6554
rect 11072 6502 11124 6554
rect 11136 6502 11188 6554
rect 20811 6502 20863 6554
rect 20875 6502 20927 6554
rect 20939 6502 20991 6554
rect 21003 6502 21055 6554
rect 21067 6502 21119 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 24492 6400 24544 6452
rect 29276 6400 29328 6452
rect 29828 6443 29880 6452
rect 29828 6409 29837 6443
rect 29837 6409 29871 6443
rect 29871 6409 29880 6443
rect 29828 6400 29880 6409
rect 24124 6332 24176 6384
rect 28080 6332 28132 6384
rect 29368 6332 29420 6384
rect 29092 6264 29144 6316
rect 22008 6196 22060 6248
rect 28724 6196 28776 6248
rect 1584 6171 1636 6180
rect 1584 6137 1593 6171
rect 1593 6137 1627 6171
rect 1627 6137 1636 6171
rect 1584 6128 1636 6137
rect 24768 6060 24820 6112
rect 27988 6060 28040 6112
rect 29368 6103 29420 6112
rect 29368 6069 29377 6103
rect 29377 6069 29411 6103
rect 29411 6069 29420 6103
rect 29368 6060 29420 6069
rect 5915 5958 5967 6010
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 15846 5958 15898 6010
rect 15910 5958 15962 6010
rect 15974 5958 16026 6010
rect 16038 5958 16090 6010
rect 16102 5958 16154 6010
rect 25776 5958 25828 6010
rect 25840 5958 25892 6010
rect 25904 5958 25956 6010
rect 25968 5958 26020 6010
rect 26032 5958 26084 6010
rect 2688 5720 2740 5772
rect 29000 5856 29052 5908
rect 29276 5856 29328 5908
rect 25596 5763 25648 5772
rect 25596 5729 25605 5763
rect 25605 5729 25639 5763
rect 25639 5729 25648 5763
rect 25596 5720 25648 5729
rect 26148 5720 26200 5772
rect 25504 5695 25556 5704
rect 25504 5661 25513 5695
rect 25513 5661 25547 5695
rect 25547 5661 25556 5695
rect 25504 5652 25556 5661
rect 24768 5584 24820 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 25320 5559 25372 5568
rect 25320 5525 25329 5559
rect 25329 5525 25363 5559
rect 25363 5525 25372 5559
rect 25320 5516 25372 5525
rect 25780 5695 25832 5704
rect 25780 5661 25789 5695
rect 25789 5661 25823 5695
rect 25823 5661 25832 5695
rect 26608 5695 26660 5704
rect 25780 5652 25832 5661
rect 26608 5661 26617 5695
rect 26617 5661 26651 5695
rect 26651 5661 26660 5695
rect 26608 5652 26660 5661
rect 27988 5695 28040 5704
rect 27988 5661 27997 5695
rect 27997 5661 28031 5695
rect 28031 5661 28040 5695
rect 27988 5652 28040 5661
rect 28816 5652 28868 5704
rect 30104 5695 30156 5704
rect 30104 5661 30113 5695
rect 30113 5661 30147 5695
rect 30147 5661 30156 5695
rect 30104 5652 30156 5661
rect 27160 5516 27212 5568
rect 10880 5414 10932 5466
rect 10944 5414 10996 5466
rect 11008 5414 11060 5466
rect 11072 5414 11124 5466
rect 11136 5414 11188 5466
rect 20811 5414 20863 5466
rect 20875 5414 20927 5466
rect 20939 5414 20991 5466
rect 21003 5414 21055 5466
rect 21067 5414 21119 5466
rect 22284 5312 22336 5364
rect 23940 5312 23992 5364
rect 22192 5244 22244 5296
rect 24676 5244 24728 5296
rect 25504 5244 25556 5296
rect 29092 5312 29144 5364
rect 29828 5355 29880 5364
rect 29828 5321 29837 5355
rect 29837 5321 29871 5355
rect 29871 5321 29880 5355
rect 29828 5312 29880 5321
rect 2688 5176 2740 5228
rect 23204 5219 23256 5228
rect 23204 5185 23213 5219
rect 23213 5185 23247 5219
rect 23247 5185 23256 5219
rect 23204 5176 23256 5185
rect 24584 5176 24636 5228
rect 25596 5219 25648 5228
rect 25596 5185 25605 5219
rect 25605 5185 25639 5219
rect 25639 5185 25648 5219
rect 25596 5176 25648 5185
rect 27068 5176 27120 5228
rect 28172 5219 28224 5228
rect 28172 5185 28181 5219
rect 28181 5185 28215 5219
rect 28215 5185 28224 5219
rect 28172 5176 28224 5185
rect 29368 5244 29420 5296
rect 29000 5176 29052 5228
rect 29092 5176 29144 5228
rect 25504 5151 25556 5160
rect 25504 5117 25513 5151
rect 25513 5117 25547 5151
rect 25547 5117 25556 5151
rect 25504 5108 25556 5117
rect 24952 5040 25004 5092
rect 25780 5151 25832 5160
rect 25780 5117 25789 5151
rect 25789 5117 25823 5151
rect 25823 5117 25832 5151
rect 25780 5108 25832 5117
rect 26148 5108 26200 5160
rect 29920 5151 29972 5160
rect 29920 5117 29929 5151
rect 29929 5117 29963 5151
rect 29963 5117 29972 5151
rect 29920 5108 29972 5117
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 24032 5015 24084 5024
rect 24032 4981 24041 5015
rect 24041 4981 24075 5015
rect 24075 4981 24084 5015
rect 24032 4972 24084 4981
rect 27436 4972 27488 5024
rect 27712 4972 27764 5024
rect 29368 5015 29420 5024
rect 29368 4981 29377 5015
rect 29377 4981 29411 5015
rect 29411 4981 29420 5015
rect 29368 4972 29420 4981
rect 5915 4870 5967 4922
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 15846 4870 15898 4922
rect 15910 4870 15962 4922
rect 15974 4870 16026 4922
rect 16038 4870 16090 4922
rect 16102 4870 16154 4922
rect 25776 4870 25828 4922
rect 25840 4870 25892 4922
rect 25904 4870 25956 4922
rect 25968 4870 26020 4922
rect 26032 4870 26084 4922
rect 23204 4768 23256 4820
rect 24584 4700 24636 4752
rect 26884 4743 26936 4752
rect 23020 4564 23072 4616
rect 23480 4564 23532 4616
rect 25320 4632 25372 4684
rect 24584 4564 24636 4616
rect 25228 4607 25280 4616
rect 25228 4573 25237 4607
rect 25237 4573 25271 4607
rect 25271 4573 25280 4607
rect 25228 4564 25280 4573
rect 25412 4607 25464 4616
rect 25412 4573 25421 4607
rect 25421 4573 25455 4607
rect 25455 4573 25464 4607
rect 25412 4564 25464 4573
rect 26884 4709 26893 4743
rect 26893 4709 26927 4743
rect 26927 4709 26936 4743
rect 26884 4700 26936 4709
rect 26148 4632 26200 4684
rect 27712 4632 27764 4684
rect 27804 4607 27856 4616
rect 27804 4573 27813 4607
rect 27813 4573 27847 4607
rect 27847 4573 27856 4607
rect 27804 4564 27856 4573
rect 28724 4675 28776 4684
rect 28724 4641 28733 4675
rect 28733 4641 28767 4675
rect 28767 4641 28776 4675
rect 28724 4632 28776 4641
rect 29000 4632 29052 4684
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 23388 4471 23440 4480
rect 23388 4437 23397 4471
rect 23397 4437 23431 4471
rect 23431 4437 23440 4471
rect 23388 4428 23440 4437
rect 23480 4428 23532 4480
rect 25136 4428 25188 4480
rect 27712 4428 27764 4480
rect 10880 4326 10932 4378
rect 10944 4326 10996 4378
rect 11008 4326 11060 4378
rect 11072 4326 11124 4378
rect 11136 4326 11188 4378
rect 20811 4326 20863 4378
rect 20875 4326 20927 4378
rect 20939 4326 20991 4378
rect 21003 4326 21055 4378
rect 21067 4326 21119 4378
rect 27712 4224 27764 4276
rect 23388 4156 23440 4208
rect 24032 4156 24084 4208
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 27436 4131 27488 4140
rect 27436 4097 27445 4131
rect 27445 4097 27479 4131
rect 27479 4097 27488 4131
rect 27436 4088 27488 4097
rect 28172 4131 28224 4140
rect 28172 4097 28181 4131
rect 28181 4097 28215 4131
rect 28215 4097 28224 4131
rect 28172 4088 28224 4097
rect 29736 4131 29788 4140
rect 29736 4097 29745 4131
rect 29745 4097 29779 4131
rect 29779 4097 29788 4131
rect 29736 4088 29788 4097
rect 22008 4063 22060 4072
rect 22008 4029 22017 4063
rect 22017 4029 22051 4063
rect 22051 4029 22060 4063
rect 22008 4020 22060 4029
rect 23940 4063 23992 4072
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 23940 4029 23949 4063
rect 23949 4029 23983 4063
rect 23983 4029 23992 4063
rect 23940 4020 23992 4029
rect 29828 4063 29880 4072
rect 29828 4029 29837 4063
rect 29837 4029 29871 4063
rect 29871 4029 29880 4063
rect 29828 4020 29880 4029
rect 29920 4063 29972 4072
rect 29920 4029 29929 4063
rect 29929 4029 29963 4063
rect 29963 4029 29972 4063
rect 29920 4020 29972 4029
rect 23388 3995 23440 4004
rect 23388 3961 23397 3995
rect 23397 3961 23431 3995
rect 23431 3961 23440 3995
rect 23388 3952 23440 3961
rect 29092 3952 29144 4004
rect 24676 3884 24728 3936
rect 27252 3927 27304 3936
rect 27252 3893 27261 3927
rect 27261 3893 27295 3927
rect 27295 3893 27304 3927
rect 27252 3884 27304 3893
rect 28632 3927 28684 3936
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 5915 3782 5967 3834
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 15846 3782 15898 3834
rect 15910 3782 15962 3834
rect 15974 3782 16026 3834
rect 16038 3782 16090 3834
rect 16102 3782 16154 3834
rect 25776 3782 25828 3834
rect 25840 3782 25892 3834
rect 25904 3782 25956 3834
rect 25968 3782 26020 3834
rect 26032 3782 26084 3834
rect 2136 3680 2188 3732
rect 28632 3680 28684 3732
rect 29736 3612 29788 3664
rect 23940 3544 23992 3596
rect 27252 3544 27304 3596
rect 25136 3519 25188 3528
rect 25136 3485 25170 3519
rect 25170 3485 25188 3519
rect 25136 3476 25188 3485
rect 28264 3519 28316 3528
rect 28264 3485 28273 3519
rect 28273 3485 28307 3519
rect 28307 3485 28316 3519
rect 28264 3476 28316 3485
rect 29368 3476 29420 3528
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 25412 3340 25464 3392
rect 28908 3383 28960 3392
rect 28908 3349 28917 3383
rect 28917 3349 28951 3383
rect 28951 3349 28960 3383
rect 28908 3340 28960 3349
rect 10880 3238 10932 3290
rect 10944 3238 10996 3290
rect 11008 3238 11060 3290
rect 11072 3238 11124 3290
rect 11136 3238 11188 3290
rect 20811 3238 20863 3290
rect 20875 3238 20927 3290
rect 20939 3238 20991 3290
rect 21003 3238 21055 3290
rect 21067 3238 21119 3290
rect 27528 3136 27580 3188
rect 26608 3068 26660 3120
rect 1492 3000 1544 3052
rect 28816 3000 28868 3052
rect 29736 3043 29788 3052
rect 29736 3009 29745 3043
rect 29745 3009 29779 3043
rect 29779 3009 29788 3043
rect 29736 3000 29788 3009
rect 1400 2796 1452 2848
rect 5915 2694 5967 2746
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 15846 2694 15898 2746
rect 15910 2694 15962 2746
rect 15974 2694 16026 2746
rect 16038 2694 16090 2746
rect 16102 2694 16154 2746
rect 25776 2694 25828 2746
rect 25840 2694 25892 2746
rect 25904 2694 25956 2746
rect 25968 2694 26020 2746
rect 26032 2694 26084 2746
rect 26884 2592 26936 2644
rect 27896 2524 27948 2576
rect 18696 2456 18748 2508
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 16856 2388 16908 2440
rect 28264 2431 28316 2440
rect 28264 2397 28273 2431
rect 28273 2397 28307 2431
rect 28307 2397 28316 2431
rect 28264 2388 28316 2397
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 29644 2431 29696 2440
rect 29644 2397 29653 2431
rect 29653 2397 29687 2431
rect 29687 2397 29696 2431
rect 29644 2388 29696 2397
rect 25044 2320 25096 2372
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2320 2295 2372 2304
rect 2320 2261 2329 2295
rect 2329 2261 2363 2295
rect 2363 2261 2372 2295
rect 2320 2252 2372 2261
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 10880 2150 10932 2202
rect 10944 2150 10996 2202
rect 11008 2150 11060 2202
rect 11072 2150 11124 2202
rect 11136 2150 11188 2202
rect 20811 2150 20863 2202
rect 20875 2150 20927 2202
rect 20939 2150 20991 2202
rect 21003 2150 21055 2202
rect 21067 2150 21119 2202
rect 22744 1300 22796 1352
rect 28724 1300 28776 1352
<< metal2 >>
rect 3790 79656 3846 79665
rect 3790 79591 3846 79600
rect 27894 79656 27950 79665
rect 27894 79591 27950 79600
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 1306 78296 1362 78305
rect 1306 78231 1362 78240
rect 1320 76498 1348 78231
rect 1398 77616 1454 77625
rect 1398 77551 1400 77560
rect 1452 77551 1454 77560
rect 1400 77522 1452 77528
rect 2792 77042 2820 78911
rect 3804 77586 3832 79591
rect 5915 77820 6223 77840
rect 5915 77818 5921 77820
rect 5977 77818 6001 77820
rect 6057 77818 6081 77820
rect 6137 77818 6161 77820
rect 6217 77818 6223 77820
rect 5977 77766 5979 77818
rect 6159 77766 6161 77818
rect 5915 77764 5921 77766
rect 5977 77764 6001 77766
rect 6057 77764 6081 77766
rect 6137 77764 6161 77766
rect 6217 77764 6223 77766
rect 5915 77744 6223 77764
rect 15846 77820 16154 77840
rect 15846 77818 15852 77820
rect 15908 77818 15932 77820
rect 15988 77818 16012 77820
rect 16068 77818 16092 77820
rect 16148 77818 16154 77820
rect 15908 77766 15910 77818
rect 16090 77766 16092 77818
rect 15846 77764 15852 77766
rect 15908 77764 15932 77766
rect 15988 77764 16012 77766
rect 16068 77764 16092 77766
rect 16148 77764 16154 77766
rect 15846 77744 16154 77764
rect 25776 77820 26084 77840
rect 25776 77818 25782 77820
rect 25838 77818 25862 77820
rect 25918 77818 25942 77820
rect 25998 77818 26022 77820
rect 26078 77818 26084 77820
rect 25838 77766 25840 77818
rect 26020 77766 26022 77818
rect 25776 77764 25782 77766
rect 25838 77764 25862 77766
rect 25918 77764 25942 77766
rect 25998 77764 26022 77766
rect 26078 77764 26084 77766
rect 25776 77744 26084 77764
rect 27908 77722 27936 79591
rect 28814 79248 28870 79257
rect 28814 79183 28870 79192
rect 28538 78704 28594 78713
rect 28538 78639 28594 78648
rect 28170 78296 28226 78305
rect 28170 78231 28226 78240
rect 28184 77722 28212 78231
rect 27896 77716 27948 77722
rect 27896 77658 27948 77664
rect 28172 77716 28224 77722
rect 28172 77658 28224 77664
rect 3792 77580 3844 77586
rect 3792 77522 3844 77528
rect 11704 77512 11756 77518
rect 11704 77454 11756 77460
rect 27252 77512 27304 77518
rect 27252 77454 27304 77460
rect 27712 77512 27764 77518
rect 27712 77454 27764 77460
rect 10880 77276 11188 77296
rect 10880 77274 10886 77276
rect 10942 77274 10966 77276
rect 11022 77274 11046 77276
rect 11102 77274 11126 77276
rect 11182 77274 11188 77276
rect 10942 77222 10944 77274
rect 11124 77222 11126 77274
rect 10880 77220 10886 77222
rect 10942 77220 10966 77222
rect 11022 77220 11046 77222
rect 11102 77220 11126 77222
rect 11182 77220 11188 77222
rect 10880 77200 11188 77220
rect 2780 77036 2832 77042
rect 2780 76978 2832 76984
rect 1400 76968 1452 76974
rect 1398 76936 1400 76945
rect 1452 76936 1454 76945
rect 1398 76871 1454 76880
rect 8300 76900 8352 76906
rect 8300 76842 8352 76848
rect 5915 76732 6223 76752
rect 5915 76730 5921 76732
rect 5977 76730 6001 76732
rect 6057 76730 6081 76732
rect 6137 76730 6161 76732
rect 6217 76730 6223 76732
rect 5977 76678 5979 76730
rect 6159 76678 6161 76730
rect 5915 76676 5921 76678
rect 5977 76676 6001 76678
rect 6057 76676 6081 76678
rect 6137 76676 6161 76678
rect 6217 76676 6223 76678
rect 5915 76656 6223 76676
rect 1308 76492 1360 76498
rect 1308 76434 1360 76440
rect 2872 76424 2924 76430
rect 2872 76366 2924 76372
rect 2884 76265 2912 76366
rect 2870 76256 2926 76265
rect 2870 76191 2926 76200
rect 1584 75948 1636 75954
rect 1584 75890 1636 75896
rect 1596 75585 1624 75890
rect 5915 75644 6223 75664
rect 5915 75642 5921 75644
rect 5977 75642 6001 75644
rect 6057 75642 6081 75644
rect 6137 75642 6161 75644
rect 6217 75642 6223 75644
rect 5977 75590 5979 75642
rect 6159 75590 6161 75642
rect 5915 75588 5921 75590
rect 5977 75588 6001 75590
rect 6057 75588 6081 75590
rect 6137 75588 6161 75590
rect 6217 75588 6223 75590
rect 1582 75576 1638 75585
rect 5915 75568 6223 75588
rect 1582 75511 1638 75520
rect 1584 75336 1636 75342
rect 1584 75278 1636 75284
rect 1596 75041 1624 75278
rect 1582 75032 1638 75041
rect 1582 74967 1638 74976
rect 1584 74860 1636 74866
rect 1584 74802 1636 74808
rect 1596 74361 1624 74802
rect 5915 74556 6223 74576
rect 5915 74554 5921 74556
rect 5977 74554 6001 74556
rect 6057 74554 6081 74556
rect 6137 74554 6161 74556
rect 6217 74554 6223 74556
rect 5977 74502 5979 74554
rect 6159 74502 6161 74554
rect 5915 74500 5921 74502
rect 5977 74500 6001 74502
rect 6057 74500 6081 74502
rect 6137 74500 6161 74502
rect 6217 74500 6223 74502
rect 5915 74480 6223 74500
rect 1582 74352 1638 74361
rect 1582 74287 1638 74296
rect 1584 73772 1636 73778
rect 1584 73714 1636 73720
rect 1596 73681 1624 73714
rect 1582 73672 1638 73681
rect 1582 73607 1638 73616
rect 5915 73468 6223 73488
rect 5915 73466 5921 73468
rect 5977 73466 6001 73468
rect 6057 73466 6081 73468
rect 6137 73466 6161 73468
rect 6217 73466 6223 73468
rect 5977 73414 5979 73466
rect 6159 73414 6161 73466
rect 5915 73412 5921 73414
rect 5977 73412 6001 73414
rect 6057 73412 6081 73414
rect 6137 73412 6161 73414
rect 6217 73412 6223 73414
rect 5915 73392 6223 73412
rect 1584 73160 1636 73166
rect 1584 73102 1636 73108
rect 1596 73001 1624 73102
rect 1582 72992 1638 73001
rect 1582 72927 1638 72936
rect 1584 72684 1636 72690
rect 1584 72626 1636 72632
rect 1596 72321 1624 72626
rect 5915 72380 6223 72400
rect 5915 72378 5921 72380
rect 5977 72378 6001 72380
rect 6057 72378 6081 72380
rect 6137 72378 6161 72380
rect 6217 72378 6223 72380
rect 5977 72326 5979 72378
rect 6159 72326 6161 72378
rect 5915 72324 5921 72326
rect 5977 72324 6001 72326
rect 6057 72324 6081 72326
rect 6137 72324 6161 72326
rect 6217 72324 6223 72326
rect 1582 72312 1638 72321
rect 5915 72304 6223 72324
rect 1582 72247 1638 72256
rect 1584 72072 1636 72078
rect 1584 72014 1636 72020
rect 1596 71641 1624 72014
rect 8312 71670 8340 76842
rect 10784 76356 10836 76362
rect 10784 76298 10836 76304
rect 9588 73092 9640 73098
rect 9588 73034 9640 73040
rect 8300 71664 8352 71670
rect 1582 71632 1638 71641
rect 8300 71606 8352 71612
rect 1582 71567 1638 71576
rect 5915 71292 6223 71312
rect 5915 71290 5921 71292
rect 5977 71290 6001 71292
rect 6057 71290 6081 71292
rect 6137 71290 6161 71292
rect 6217 71290 6223 71292
rect 5977 71238 5979 71290
rect 6159 71238 6161 71290
rect 5915 71236 5921 71238
rect 5977 71236 6001 71238
rect 6057 71236 6081 71238
rect 6137 71236 6161 71238
rect 6217 71236 6223 71238
rect 5915 71216 6223 71236
rect 1492 71052 1544 71058
rect 1492 70994 1544 71000
rect 1400 70984 1452 70990
rect 1398 70952 1400 70961
rect 1452 70952 1454 70961
rect 1398 70887 1454 70896
rect 1504 70650 1532 70994
rect 9600 70990 9628 73034
rect 10232 73024 10284 73030
rect 10232 72966 10284 72972
rect 10244 72758 10272 72966
rect 10232 72752 10284 72758
rect 10232 72694 10284 72700
rect 9588 70984 9640 70990
rect 9588 70926 9640 70932
rect 1492 70644 1544 70650
rect 1492 70586 1544 70592
rect 1584 70508 1636 70514
rect 1584 70450 1636 70456
rect 1596 70417 1624 70450
rect 1582 70408 1638 70417
rect 1582 70343 1638 70352
rect 5915 70204 6223 70224
rect 5915 70202 5921 70204
rect 5977 70202 6001 70204
rect 6057 70202 6081 70204
rect 6137 70202 6161 70204
rect 6217 70202 6223 70204
rect 5977 70150 5979 70202
rect 6159 70150 6161 70202
rect 5915 70148 5921 70150
rect 5977 70148 6001 70150
rect 6057 70148 6081 70150
rect 6137 70148 6161 70150
rect 6217 70148 6223 70150
rect 5915 70128 6223 70148
rect 10796 69902 10824 76298
rect 10880 76188 11188 76208
rect 10880 76186 10886 76188
rect 10942 76186 10966 76188
rect 11022 76186 11046 76188
rect 11102 76186 11126 76188
rect 11182 76186 11188 76188
rect 10942 76134 10944 76186
rect 11124 76134 11126 76186
rect 10880 76132 10886 76134
rect 10942 76132 10966 76134
rect 11022 76132 11046 76134
rect 11102 76132 11126 76134
rect 11182 76132 11188 76134
rect 10880 76112 11188 76132
rect 10880 75100 11188 75120
rect 10880 75098 10886 75100
rect 10942 75098 10966 75100
rect 11022 75098 11046 75100
rect 11102 75098 11126 75100
rect 11182 75098 11188 75100
rect 10942 75046 10944 75098
rect 11124 75046 11126 75098
rect 10880 75044 10886 75046
rect 10942 75044 10966 75046
rect 11022 75044 11046 75046
rect 11102 75044 11126 75046
rect 11182 75044 11188 75046
rect 10880 75024 11188 75044
rect 10880 74012 11188 74032
rect 10880 74010 10886 74012
rect 10942 74010 10966 74012
rect 11022 74010 11046 74012
rect 11102 74010 11126 74012
rect 11182 74010 11188 74012
rect 10942 73958 10944 74010
rect 11124 73958 11126 74010
rect 10880 73956 10886 73958
rect 10942 73956 10966 73958
rect 11022 73956 11046 73958
rect 11102 73956 11126 73958
rect 11182 73956 11188 73958
rect 10880 73936 11188 73956
rect 10880 72924 11188 72944
rect 10880 72922 10886 72924
rect 10942 72922 10966 72924
rect 11022 72922 11046 72924
rect 11102 72922 11126 72924
rect 11182 72922 11188 72924
rect 10942 72870 10944 72922
rect 11124 72870 11126 72922
rect 10880 72868 10886 72870
rect 10942 72868 10966 72870
rect 11022 72868 11046 72870
rect 11102 72868 11126 72870
rect 11182 72868 11188 72870
rect 10880 72848 11188 72868
rect 10880 71836 11188 71856
rect 10880 71834 10886 71836
rect 10942 71834 10966 71836
rect 11022 71834 11046 71836
rect 11102 71834 11126 71836
rect 11182 71834 11188 71836
rect 10942 71782 10944 71834
rect 11124 71782 11126 71834
rect 10880 71780 10886 71782
rect 10942 71780 10966 71782
rect 11022 71780 11046 71782
rect 11102 71780 11126 71782
rect 11182 71780 11188 71782
rect 10880 71760 11188 71780
rect 10880 70748 11188 70768
rect 10880 70746 10886 70748
rect 10942 70746 10966 70748
rect 11022 70746 11046 70748
rect 11102 70746 11126 70748
rect 11182 70746 11188 70748
rect 10942 70694 10944 70746
rect 11124 70694 11126 70746
rect 10880 70692 10886 70694
rect 10942 70692 10966 70694
rect 11022 70692 11046 70694
rect 11102 70692 11126 70694
rect 11182 70692 11188 70694
rect 10880 70672 11188 70692
rect 11716 70582 11744 77454
rect 27160 77444 27212 77450
rect 27160 77386 27212 77392
rect 11796 77376 11848 77382
rect 11796 77318 11848 77324
rect 11808 70990 11836 77318
rect 20811 77276 21119 77296
rect 20811 77274 20817 77276
rect 20873 77274 20897 77276
rect 20953 77274 20977 77276
rect 21033 77274 21057 77276
rect 21113 77274 21119 77276
rect 20873 77222 20875 77274
rect 21055 77222 21057 77274
rect 20811 77220 20817 77222
rect 20873 77220 20897 77222
rect 20953 77220 20977 77222
rect 21033 77220 21057 77222
rect 21113 77220 21119 77222
rect 20811 77200 21119 77220
rect 13728 76968 13780 76974
rect 13728 76910 13780 76916
rect 13544 73772 13596 73778
rect 13544 73714 13596 73720
rect 13556 72078 13584 73714
rect 13544 72072 13596 72078
rect 13544 72014 13596 72020
rect 12808 71596 12860 71602
rect 12808 71538 12860 71544
rect 11796 70984 11848 70990
rect 11796 70926 11848 70932
rect 12820 70922 12848 71538
rect 12808 70916 12860 70922
rect 12808 70858 12860 70864
rect 12820 70650 12848 70858
rect 12808 70644 12860 70650
rect 12808 70586 12860 70592
rect 11704 70576 11756 70582
rect 11704 70518 11756 70524
rect 12820 70514 12848 70586
rect 12808 70508 12860 70514
rect 12808 70450 12860 70456
rect 12820 69902 12848 70450
rect 13556 70446 13584 72014
rect 13740 70514 13768 76910
rect 15846 76732 16154 76752
rect 15846 76730 15852 76732
rect 15908 76730 15932 76732
rect 15988 76730 16012 76732
rect 16068 76730 16092 76732
rect 16148 76730 16154 76732
rect 15908 76678 15910 76730
rect 16090 76678 16092 76730
rect 15846 76676 15852 76678
rect 15908 76676 15932 76678
rect 15988 76676 16012 76678
rect 16068 76676 16092 76678
rect 16148 76676 16154 76678
rect 15846 76656 16154 76676
rect 25776 76732 26084 76752
rect 25776 76730 25782 76732
rect 25838 76730 25862 76732
rect 25918 76730 25942 76732
rect 25998 76730 26022 76732
rect 26078 76730 26084 76732
rect 25838 76678 25840 76730
rect 26020 76678 26022 76730
rect 25776 76676 25782 76678
rect 25838 76676 25862 76678
rect 25918 76676 25942 76678
rect 25998 76676 26022 76678
rect 26078 76676 26084 76678
rect 25776 76656 26084 76676
rect 26332 76424 26384 76430
rect 26332 76366 26384 76372
rect 14648 76288 14700 76294
rect 14648 76230 14700 76236
rect 19984 76288 20036 76294
rect 19984 76230 20036 76236
rect 21180 76288 21232 76294
rect 21180 76230 21232 76236
rect 14556 76084 14608 76090
rect 14556 76026 14608 76032
rect 14464 75948 14516 75954
rect 14464 75890 14516 75896
rect 14476 75274 14504 75890
rect 14568 75342 14596 76026
rect 14660 76022 14688 76230
rect 14648 76016 14700 76022
rect 14648 75958 14700 75964
rect 15292 76016 15344 76022
rect 15292 75958 15344 75964
rect 15200 75744 15252 75750
rect 15200 75686 15252 75692
rect 15212 75410 15240 75686
rect 15200 75404 15252 75410
rect 15200 75346 15252 75352
rect 14556 75336 14608 75342
rect 14556 75278 14608 75284
rect 14464 75268 14516 75274
rect 14464 75210 14516 75216
rect 14476 75154 14504 75210
rect 14648 75200 14700 75206
rect 14476 75126 14596 75154
rect 14648 75142 14700 75148
rect 14568 74866 14596 75126
rect 14660 74934 14688 75142
rect 15304 75002 15332 75958
rect 19996 75954 20024 76230
rect 20811 76188 21119 76208
rect 20811 76186 20817 76188
rect 20873 76186 20897 76188
rect 20953 76186 20977 76188
rect 21033 76186 21057 76188
rect 21113 76186 21119 76188
rect 20873 76134 20875 76186
rect 21055 76134 21057 76186
rect 20811 76132 20817 76134
rect 20873 76132 20897 76134
rect 20953 76132 20977 76134
rect 21033 76132 21057 76134
rect 21113 76132 21119 76134
rect 20811 76112 21119 76132
rect 15752 75948 15804 75954
rect 15752 75890 15804 75896
rect 16764 75948 16816 75954
rect 16764 75890 16816 75896
rect 19064 75948 19116 75954
rect 19064 75890 19116 75896
rect 19984 75948 20036 75954
rect 19984 75890 20036 75896
rect 20168 75948 20220 75954
rect 20168 75890 20220 75896
rect 15292 74996 15344 75002
rect 15292 74938 15344 74944
rect 14648 74928 14700 74934
rect 14648 74870 14700 74876
rect 14556 74860 14608 74866
rect 14556 74802 14608 74808
rect 14568 74186 14596 74802
rect 15764 74458 15792 75890
rect 15846 75644 16154 75664
rect 15846 75642 15852 75644
rect 15908 75642 15932 75644
rect 15988 75642 16012 75644
rect 16068 75642 16092 75644
rect 16148 75642 16154 75644
rect 15908 75590 15910 75642
rect 16090 75590 16092 75642
rect 15846 75588 15852 75590
rect 15908 75588 15932 75590
rect 15988 75588 16012 75590
rect 16068 75588 16092 75590
rect 16148 75588 16154 75590
rect 15846 75568 16154 75588
rect 16672 75268 16724 75274
rect 16672 75210 16724 75216
rect 16488 74860 16540 74866
rect 16488 74802 16540 74808
rect 15846 74556 16154 74576
rect 15846 74554 15852 74556
rect 15908 74554 15932 74556
rect 15988 74554 16012 74556
rect 16068 74554 16092 74556
rect 16148 74554 16154 74556
rect 15908 74502 15910 74554
rect 16090 74502 16092 74554
rect 15846 74500 15852 74502
rect 15908 74500 15932 74502
rect 15988 74500 16012 74502
rect 16068 74500 16092 74502
rect 16148 74500 16154 74502
rect 15846 74480 16154 74500
rect 15752 74452 15804 74458
rect 15752 74394 15804 74400
rect 16500 74322 16528 74802
rect 16580 74792 16632 74798
rect 16580 74734 16632 74740
rect 16488 74316 16540 74322
rect 16488 74258 16540 74264
rect 14556 74180 14608 74186
rect 14556 74122 14608 74128
rect 14740 74180 14792 74186
rect 14740 74122 14792 74128
rect 14568 73914 14596 74122
rect 14556 73908 14608 73914
rect 14556 73850 14608 73856
rect 14752 73642 14780 74122
rect 14740 73636 14792 73642
rect 14740 73578 14792 73584
rect 15846 73468 16154 73488
rect 15846 73466 15852 73468
rect 15908 73466 15932 73468
rect 15988 73466 16012 73468
rect 16068 73466 16092 73468
rect 16148 73466 16154 73468
rect 15908 73414 15910 73466
rect 16090 73414 16092 73466
rect 15846 73412 15852 73414
rect 15908 73412 15932 73414
rect 15988 73412 16012 73414
rect 16068 73412 16092 73414
rect 16148 73412 16154 73414
rect 15846 73392 16154 73412
rect 15844 73160 15896 73166
rect 15842 73128 15844 73137
rect 15896 73128 15898 73137
rect 14648 73092 14700 73098
rect 14648 73034 14700 73040
rect 14740 73092 14792 73098
rect 14740 73034 14792 73040
rect 14924 73092 14976 73098
rect 15842 73063 15898 73072
rect 14924 73034 14976 73040
rect 14660 72690 14688 73034
rect 14648 72684 14700 72690
rect 14648 72626 14700 72632
rect 14660 72282 14688 72626
rect 14648 72276 14700 72282
rect 14648 72218 14700 72224
rect 14660 72078 14688 72218
rect 14752 72214 14780 73034
rect 14936 72690 14964 73034
rect 16500 72758 16528 74258
rect 16592 74186 16620 74734
rect 16580 74180 16632 74186
rect 16580 74122 16632 74128
rect 16488 72752 16540 72758
rect 16488 72694 16540 72700
rect 14924 72684 14976 72690
rect 14924 72626 14976 72632
rect 14832 72480 14884 72486
rect 14832 72422 14884 72428
rect 14740 72208 14792 72214
rect 14740 72150 14792 72156
rect 14844 72078 14872 72422
rect 15846 72380 16154 72400
rect 15846 72378 15852 72380
rect 15908 72378 15932 72380
rect 15988 72378 16012 72380
rect 16068 72378 16092 72380
rect 16148 72378 16154 72380
rect 15908 72326 15910 72378
rect 16090 72326 16092 72378
rect 15846 72324 15852 72326
rect 15908 72324 15932 72326
rect 15988 72324 16012 72326
rect 16068 72324 16092 72326
rect 16148 72324 16154 72326
rect 15846 72304 16154 72324
rect 14648 72072 14700 72078
rect 14648 72014 14700 72020
rect 14832 72072 14884 72078
rect 14832 72014 14884 72020
rect 14660 70922 14688 72014
rect 15846 71292 16154 71312
rect 15846 71290 15852 71292
rect 15908 71290 15932 71292
rect 15988 71290 16012 71292
rect 16068 71290 16092 71292
rect 16148 71290 16154 71292
rect 15908 71238 15910 71290
rect 16090 71238 16092 71290
rect 15846 71236 15852 71238
rect 15908 71236 15932 71238
rect 15988 71236 16012 71238
rect 16068 71236 16092 71238
rect 16148 71236 16154 71238
rect 15846 71216 16154 71236
rect 16396 71188 16448 71194
rect 16396 71130 16448 71136
rect 14648 70916 14700 70922
rect 14648 70858 14700 70864
rect 15568 70848 15620 70854
rect 15568 70790 15620 70796
rect 15476 70576 15528 70582
rect 15476 70518 15528 70524
rect 13728 70508 13780 70514
rect 13728 70450 13780 70456
rect 13544 70440 13596 70446
rect 13544 70382 13596 70388
rect 14832 70440 14884 70446
rect 14884 70388 14964 70394
rect 14832 70382 14964 70388
rect 1584 69896 1636 69902
rect 1584 69838 1636 69844
rect 10784 69896 10836 69902
rect 10784 69838 10836 69844
rect 12808 69896 12860 69902
rect 12808 69838 12860 69844
rect 1596 69737 1624 69838
rect 9956 69760 10008 69766
rect 1582 69728 1638 69737
rect 9956 69702 10008 69708
rect 1582 69663 1638 69672
rect 9968 69494 9996 69702
rect 10880 69660 11188 69680
rect 10880 69658 10886 69660
rect 10942 69658 10966 69660
rect 11022 69658 11046 69660
rect 11102 69658 11126 69660
rect 11182 69658 11188 69660
rect 10942 69606 10944 69658
rect 11124 69606 11126 69658
rect 10880 69604 10886 69606
rect 10942 69604 10966 69606
rect 11022 69604 11046 69606
rect 11102 69604 11126 69606
rect 11182 69604 11188 69606
rect 10880 69584 11188 69604
rect 9956 69488 10008 69494
rect 9956 69430 10008 69436
rect 1584 69420 1636 69426
rect 1584 69362 1636 69368
rect 12624 69420 12676 69426
rect 12624 69362 12676 69368
rect 1596 69057 1624 69362
rect 11336 69216 11388 69222
rect 11336 69158 11388 69164
rect 5915 69116 6223 69136
rect 5915 69114 5921 69116
rect 5977 69114 6001 69116
rect 6057 69114 6081 69116
rect 6137 69114 6161 69116
rect 6217 69114 6223 69116
rect 5977 69062 5979 69114
rect 6159 69062 6161 69114
rect 5915 69060 5921 69062
rect 5977 69060 6001 69062
rect 6057 69060 6081 69062
rect 6137 69060 6161 69062
rect 6217 69060 6223 69062
rect 1582 69048 1638 69057
rect 5915 69040 6223 69060
rect 1582 68983 1638 68992
rect 1584 68808 1636 68814
rect 1584 68750 1636 68756
rect 1400 68672 1452 68678
rect 1400 68614 1452 68620
rect 1412 68474 1440 68614
rect 1400 68468 1452 68474
rect 1400 68410 1452 68416
rect 1596 68377 1624 68750
rect 10880 68572 11188 68592
rect 10880 68570 10886 68572
rect 10942 68570 10966 68572
rect 11022 68570 11046 68572
rect 11102 68570 11126 68572
rect 11182 68570 11188 68572
rect 10942 68518 10944 68570
rect 11124 68518 11126 68570
rect 10880 68516 10886 68518
rect 10942 68516 10966 68518
rect 11022 68516 11046 68518
rect 11102 68516 11126 68518
rect 11182 68516 11188 68518
rect 10880 68496 11188 68516
rect 1582 68368 1638 68377
rect 1582 68303 1638 68312
rect 5915 68028 6223 68048
rect 5915 68026 5921 68028
rect 5977 68026 6001 68028
rect 6057 68026 6081 68028
rect 6137 68026 6161 68028
rect 6217 68026 6223 68028
rect 5977 67974 5979 68026
rect 6159 67974 6161 68026
rect 5915 67972 5921 67974
rect 5977 67972 6001 67974
rect 6057 67972 6081 67974
rect 6137 67972 6161 67974
rect 6217 67972 6223 67974
rect 5915 67952 6223 67972
rect 11244 67856 11296 67862
rect 11244 67798 11296 67804
rect 1584 67720 1636 67726
rect 1582 67688 1584 67697
rect 1636 67688 1638 67697
rect 1582 67623 1638 67632
rect 10880 67484 11188 67504
rect 10880 67482 10886 67484
rect 10942 67482 10966 67484
rect 11022 67482 11046 67484
rect 11102 67482 11126 67484
rect 11182 67482 11188 67484
rect 10942 67430 10944 67482
rect 11124 67430 11126 67482
rect 10880 67428 10886 67430
rect 10942 67428 10966 67430
rect 11022 67428 11046 67430
rect 11102 67428 11126 67430
rect 11182 67428 11188 67430
rect 10880 67408 11188 67428
rect 11256 67318 11284 67798
rect 11348 67726 11376 69158
rect 12636 68814 12664 69362
rect 12624 68808 12676 68814
rect 12624 68750 12676 68756
rect 11336 67720 11388 67726
rect 11336 67662 11388 67668
rect 12636 67658 12664 68750
rect 12808 68740 12860 68746
rect 12808 68682 12860 68688
rect 12820 68474 12848 68682
rect 12808 68468 12860 68474
rect 12808 68410 12860 68416
rect 12624 67652 12676 67658
rect 12624 67594 12676 67600
rect 11244 67312 11296 67318
rect 11244 67254 11296 67260
rect 12636 67250 12664 67594
rect 13084 67584 13136 67590
rect 13084 67526 13136 67532
rect 13096 67318 13124 67526
rect 13084 67312 13136 67318
rect 13084 67254 13136 67260
rect 1584 67244 1636 67250
rect 1584 67186 1636 67192
rect 12624 67244 12676 67250
rect 12624 67186 12676 67192
rect 1596 67017 1624 67186
rect 11244 67040 11296 67046
rect 1582 67008 1638 67017
rect 11244 66982 11296 66988
rect 1582 66943 1638 66952
rect 5915 66940 6223 66960
rect 5915 66938 5921 66940
rect 5977 66938 6001 66940
rect 6057 66938 6081 66940
rect 6137 66938 6161 66940
rect 6217 66938 6223 66940
rect 5977 66886 5979 66938
rect 6159 66886 6161 66938
rect 5915 66884 5921 66886
rect 5977 66884 6001 66886
rect 6057 66884 6081 66886
rect 6137 66884 6161 66886
rect 6217 66884 6223 66886
rect 5915 66864 6223 66884
rect 1584 66632 1636 66638
rect 1584 66574 1636 66580
rect 1596 66337 1624 66574
rect 10880 66396 11188 66416
rect 10880 66394 10886 66396
rect 10942 66394 10966 66396
rect 11022 66394 11046 66396
rect 11102 66394 11126 66396
rect 11182 66394 11188 66396
rect 10942 66342 10944 66394
rect 11124 66342 11126 66394
rect 10880 66340 10886 66342
rect 10942 66340 10966 66342
rect 11022 66340 11046 66342
rect 11102 66340 11126 66342
rect 11182 66340 11188 66342
rect 1582 66328 1638 66337
rect 10880 66320 11188 66340
rect 1582 66263 1638 66272
rect 11256 66230 11284 66982
rect 11336 66496 11388 66502
rect 11336 66438 11388 66444
rect 11244 66224 11296 66230
rect 11244 66166 11296 66172
rect 1584 66156 1636 66162
rect 1584 66098 1636 66104
rect 1596 65793 1624 66098
rect 5915 65852 6223 65872
rect 5915 65850 5921 65852
rect 5977 65850 6001 65852
rect 6057 65850 6081 65852
rect 6137 65850 6161 65852
rect 6217 65850 6223 65852
rect 5977 65798 5979 65850
rect 6159 65798 6161 65850
rect 5915 65796 5921 65798
rect 5977 65796 6001 65798
rect 6057 65796 6081 65798
rect 6137 65796 6161 65798
rect 6217 65796 6223 65798
rect 1582 65784 1638 65793
rect 5915 65776 6223 65796
rect 1582 65719 1638 65728
rect 1584 65544 1636 65550
rect 1584 65486 1636 65492
rect 1596 65113 1624 65486
rect 11244 65408 11296 65414
rect 11244 65350 11296 65356
rect 10880 65308 11188 65328
rect 10880 65306 10886 65308
rect 10942 65306 10966 65308
rect 11022 65306 11046 65308
rect 11102 65306 11126 65308
rect 11182 65306 11188 65308
rect 10942 65254 10944 65306
rect 11124 65254 11126 65306
rect 10880 65252 10886 65254
rect 10942 65252 10966 65254
rect 11022 65252 11046 65254
rect 11102 65252 11126 65254
rect 11182 65252 11188 65254
rect 10880 65232 11188 65252
rect 1582 65104 1638 65113
rect 1582 65039 1638 65048
rect 5915 64764 6223 64784
rect 5915 64762 5921 64764
rect 5977 64762 6001 64764
rect 6057 64762 6081 64764
rect 6137 64762 6161 64764
rect 6217 64762 6223 64764
rect 5977 64710 5979 64762
rect 6159 64710 6161 64762
rect 5915 64708 5921 64710
rect 5977 64708 6001 64710
rect 6057 64708 6081 64710
rect 6137 64708 6161 64710
rect 6217 64708 6223 64710
rect 5915 64688 6223 64708
rect 11256 64462 11284 65350
rect 1584 64456 1636 64462
rect 1582 64424 1584 64433
rect 11244 64456 11296 64462
rect 1636 64424 1638 64433
rect 11244 64398 11296 64404
rect 1582 64359 1638 64368
rect 10880 64220 11188 64240
rect 10880 64218 10886 64220
rect 10942 64218 10966 64220
rect 11022 64218 11046 64220
rect 11102 64218 11126 64220
rect 11182 64218 11188 64220
rect 10942 64166 10944 64218
rect 11124 64166 11126 64218
rect 10880 64164 10886 64166
rect 10942 64164 10966 64166
rect 11022 64164 11046 64166
rect 11102 64164 11126 64166
rect 11182 64164 11188 64166
rect 10880 64144 11188 64164
rect 11348 64122 11376 66438
rect 12636 66162 12664 67186
rect 12624 66156 12676 66162
rect 12624 66098 12676 66104
rect 11428 65952 11480 65958
rect 11428 65894 11480 65900
rect 11336 64116 11388 64122
rect 11336 64058 11388 64064
rect 1584 63980 1636 63986
rect 1584 63922 1636 63928
rect 1596 63753 1624 63922
rect 11336 63776 11388 63782
rect 1582 63744 1638 63753
rect 11336 63718 11388 63724
rect 1582 63679 1638 63688
rect 5915 63676 6223 63696
rect 5915 63674 5921 63676
rect 5977 63674 6001 63676
rect 6057 63674 6081 63676
rect 6137 63674 6161 63676
rect 6217 63674 6223 63676
rect 5977 63622 5979 63674
rect 6159 63622 6161 63674
rect 5915 63620 5921 63622
rect 5977 63620 6001 63622
rect 6057 63620 6081 63622
rect 6137 63620 6161 63622
rect 6217 63620 6223 63622
rect 5915 63600 6223 63620
rect 1584 63368 1636 63374
rect 1584 63310 1636 63316
rect 1596 63073 1624 63310
rect 11244 63232 11296 63238
rect 11244 63174 11296 63180
rect 10880 63132 11188 63152
rect 10880 63130 10886 63132
rect 10942 63130 10966 63132
rect 11022 63130 11046 63132
rect 11102 63130 11126 63132
rect 11182 63130 11188 63132
rect 10942 63078 10944 63130
rect 11124 63078 11126 63130
rect 10880 63076 10886 63078
rect 10942 63076 10966 63078
rect 11022 63076 11046 63078
rect 11102 63076 11126 63078
rect 11182 63076 11188 63078
rect 1582 63064 1638 63073
rect 10880 63056 11188 63076
rect 1582 62999 1638 63008
rect 1584 62892 1636 62898
rect 1584 62834 1636 62840
rect 1596 62393 1624 62834
rect 5915 62588 6223 62608
rect 5915 62586 5921 62588
rect 5977 62586 6001 62588
rect 6057 62586 6081 62588
rect 6137 62586 6161 62588
rect 6217 62586 6223 62588
rect 5977 62534 5979 62586
rect 6159 62534 6161 62586
rect 5915 62532 5921 62534
rect 5977 62532 6001 62534
rect 6057 62532 6081 62534
rect 6137 62532 6161 62534
rect 6217 62532 6223 62534
rect 5915 62512 6223 62532
rect 1582 62384 1638 62393
rect 1582 62319 1638 62328
rect 10880 62044 11188 62064
rect 10880 62042 10886 62044
rect 10942 62042 10966 62044
rect 11022 62042 11046 62044
rect 11102 62042 11126 62044
rect 11182 62042 11188 62044
rect 10942 61990 10944 62042
rect 11124 61990 11126 62042
rect 10880 61988 10886 61990
rect 10942 61988 10966 61990
rect 11022 61988 11046 61990
rect 11102 61988 11126 61990
rect 11182 61988 11188 61990
rect 10880 61968 11188 61988
rect 11256 61878 11284 63174
rect 11348 62966 11376 63718
rect 11440 63306 11468 65894
rect 12636 65754 12664 66098
rect 12992 65952 13044 65958
rect 12992 65894 13044 65900
rect 12624 65748 12676 65754
rect 12624 65690 12676 65696
rect 12900 65544 12952 65550
rect 12900 65486 12952 65492
rect 12912 65074 12940 65486
rect 12900 65068 12952 65074
rect 12900 65010 12952 65016
rect 12716 64864 12768 64870
rect 12716 64806 12768 64812
rect 12728 64394 12756 64806
rect 12716 64388 12768 64394
rect 12716 64330 12768 64336
rect 12164 64320 12216 64326
rect 12164 64262 12216 64268
rect 12176 64054 12204 64262
rect 12164 64048 12216 64054
rect 12164 63990 12216 63996
rect 12728 63986 12756 64330
rect 12716 63980 12768 63986
rect 12716 63922 12768 63928
rect 12728 63306 12756 63922
rect 11428 63300 11480 63306
rect 11428 63242 11480 63248
rect 12716 63300 12768 63306
rect 12716 63242 12768 63248
rect 11336 62960 11388 62966
rect 11336 62902 11388 62908
rect 12728 62898 12756 63242
rect 12716 62892 12768 62898
rect 12716 62834 12768 62840
rect 11336 62688 11388 62694
rect 11336 62630 11388 62636
rect 11244 61872 11296 61878
rect 11244 61814 11296 61820
rect 1584 61804 1636 61810
rect 1584 61746 1636 61752
rect 1596 61713 1624 61746
rect 1582 61704 1638 61713
rect 1582 61639 1638 61648
rect 7564 61600 7616 61606
rect 7564 61542 7616 61548
rect 5915 61500 6223 61520
rect 5915 61498 5921 61500
rect 5977 61498 6001 61500
rect 6057 61498 6081 61500
rect 6137 61498 6161 61500
rect 6217 61498 6223 61500
rect 5977 61446 5979 61498
rect 6159 61446 6161 61498
rect 5915 61444 5921 61446
rect 5977 61444 6001 61446
rect 6057 61444 6081 61446
rect 6137 61444 6161 61446
rect 6217 61444 6223 61446
rect 5915 61424 6223 61444
rect 7576 61266 7604 61542
rect 7564 61260 7616 61266
rect 7564 61202 7616 61208
rect 1584 61192 1636 61198
rect 1582 61160 1584 61169
rect 1636 61160 1638 61169
rect 1582 61095 1638 61104
rect 11244 61056 11296 61062
rect 11244 60998 11296 61004
rect 10880 60956 11188 60976
rect 10880 60954 10886 60956
rect 10942 60954 10966 60956
rect 11022 60954 11046 60956
rect 11102 60954 11126 60956
rect 11182 60954 11188 60956
rect 10942 60902 10944 60954
rect 11124 60902 11126 60954
rect 10880 60900 10886 60902
rect 10942 60900 10966 60902
rect 11022 60900 11046 60902
rect 11102 60900 11126 60902
rect 11182 60900 11188 60902
rect 10880 60880 11188 60900
rect 1584 60716 1636 60722
rect 1584 60658 1636 60664
rect 1596 60489 1624 60658
rect 1582 60480 1638 60489
rect 1582 60415 1638 60424
rect 5915 60412 6223 60432
rect 5915 60410 5921 60412
rect 5977 60410 6001 60412
rect 6057 60410 6081 60412
rect 6137 60410 6161 60412
rect 6217 60410 6223 60412
rect 5977 60358 5979 60410
rect 6159 60358 6161 60410
rect 5915 60356 5921 60358
rect 5977 60356 6001 60358
rect 6057 60356 6081 60358
rect 6137 60356 6161 60358
rect 6217 60356 6223 60358
rect 5915 60336 6223 60356
rect 11256 60110 11284 60998
rect 11348 60654 11376 62630
rect 12532 61804 12584 61810
rect 12532 61746 12584 61752
rect 12544 61062 12572 61746
rect 12912 61198 12940 65010
rect 12900 61192 12952 61198
rect 12900 61134 12952 61140
rect 12532 61056 12584 61062
rect 12532 60998 12584 61004
rect 12544 60790 12572 60998
rect 12532 60784 12584 60790
rect 12532 60726 12584 60732
rect 11336 60648 11388 60654
rect 11336 60590 11388 60596
rect 12544 60110 12572 60726
rect 12716 60512 12768 60518
rect 12716 60454 12768 60460
rect 12900 60512 12952 60518
rect 12900 60454 12952 60460
rect 1584 60104 1636 60110
rect 1584 60046 1636 60052
rect 11244 60104 11296 60110
rect 11244 60046 11296 60052
rect 12532 60104 12584 60110
rect 12532 60046 12584 60052
rect 1596 59809 1624 60046
rect 11336 59968 11388 59974
rect 11336 59910 11388 59916
rect 10880 59868 11188 59888
rect 10880 59866 10886 59868
rect 10942 59866 10966 59868
rect 11022 59866 11046 59868
rect 11102 59866 11126 59868
rect 11182 59866 11188 59868
rect 10942 59814 10944 59866
rect 11124 59814 11126 59866
rect 10880 59812 10886 59814
rect 10942 59812 10966 59814
rect 11022 59812 11046 59814
rect 11102 59812 11126 59814
rect 11182 59812 11188 59814
rect 1582 59800 1638 59809
rect 10880 59792 11188 59812
rect 1582 59735 1638 59744
rect 1584 59628 1636 59634
rect 1584 59570 1636 59576
rect 1596 59129 1624 59570
rect 11244 59424 11296 59430
rect 11244 59366 11296 59372
rect 5915 59324 6223 59344
rect 5915 59322 5921 59324
rect 5977 59322 6001 59324
rect 6057 59322 6081 59324
rect 6137 59322 6161 59324
rect 6217 59322 6223 59324
rect 5977 59270 5979 59322
rect 6159 59270 6161 59322
rect 5915 59268 5921 59270
rect 5977 59268 6001 59270
rect 6057 59268 6081 59270
rect 6137 59268 6161 59270
rect 6217 59268 6223 59270
rect 5915 59248 6223 59268
rect 1582 59120 1638 59129
rect 1582 59055 1638 59064
rect 10880 58780 11188 58800
rect 10880 58778 10886 58780
rect 10942 58778 10966 58780
rect 11022 58778 11046 58780
rect 11102 58778 11126 58780
rect 11182 58778 11188 58780
rect 10942 58726 10944 58778
rect 11124 58726 11126 58778
rect 10880 58724 10886 58726
rect 10942 58724 10966 58726
rect 11022 58724 11046 58726
rect 11102 58724 11126 58726
rect 11182 58724 11188 58726
rect 10880 58704 11188 58724
rect 11256 58614 11284 59366
rect 11348 59022 11376 59910
rect 12544 59702 12572 60046
rect 12728 59702 12756 60454
rect 12532 59696 12584 59702
rect 12532 59638 12584 59644
rect 12716 59696 12768 59702
rect 12716 59638 12768 59644
rect 12912 59566 12940 60454
rect 12900 59560 12952 59566
rect 12900 59502 12952 59508
rect 11336 59016 11388 59022
rect 11336 58958 11388 58964
rect 11244 58608 11296 58614
rect 11244 58550 11296 58556
rect 1400 58540 1452 58546
rect 1400 58482 1452 58488
rect 1412 57594 1440 58482
rect 1582 58440 1638 58449
rect 1582 58375 1584 58384
rect 1636 58375 1638 58384
rect 1584 58346 1636 58352
rect 5915 58236 6223 58256
rect 5915 58234 5921 58236
rect 5977 58234 6001 58236
rect 6057 58234 6081 58236
rect 6137 58234 6161 58236
rect 6217 58234 6223 58236
rect 5977 58182 5979 58234
rect 6159 58182 6161 58234
rect 5915 58180 5921 58182
rect 5977 58180 6001 58182
rect 6057 58180 6081 58182
rect 6137 58180 6161 58182
rect 6217 58180 6223 58182
rect 5915 58160 6223 58180
rect 2136 57928 2188 57934
rect 2136 57870 2188 57876
rect 1584 57792 1636 57798
rect 1582 57760 1584 57769
rect 1636 57760 1638 57769
rect 1582 57695 1638 57704
rect 1400 57588 1452 57594
rect 1400 57530 1452 57536
rect 1860 57452 1912 57458
rect 1860 57394 1912 57400
rect 1584 57248 1636 57254
rect 1584 57190 1636 57196
rect 1596 57089 1624 57190
rect 1582 57080 1638 57089
rect 1582 57015 1638 57024
rect 1400 56840 1452 56846
rect 1400 56782 1452 56788
rect 1412 55962 1440 56782
rect 1584 56704 1636 56710
rect 1584 56646 1636 56652
rect 1596 56545 1624 56646
rect 1582 56536 1638 56545
rect 1872 56506 1900 57394
rect 2148 57050 2176 57870
rect 13004 57798 13032 65894
rect 13452 61192 13504 61198
rect 13452 61134 13504 61140
rect 13464 59634 13492 61134
rect 13556 59770 13584 70382
rect 14844 70366 14964 70382
rect 14648 69828 14700 69834
rect 14648 69770 14700 69776
rect 14004 69420 14056 69426
rect 14004 69362 14056 69368
rect 13912 69352 13964 69358
rect 13912 69294 13964 69300
rect 13924 68474 13952 69294
rect 13912 68468 13964 68474
rect 13912 68410 13964 68416
rect 13820 68332 13872 68338
rect 13820 68274 13872 68280
rect 13728 66088 13780 66094
rect 13728 66030 13780 66036
rect 13740 65210 13768 66030
rect 13728 65204 13780 65210
rect 13728 65146 13780 65152
rect 13832 63510 13860 68274
rect 14016 68202 14044 69362
rect 14660 69018 14688 69770
rect 14832 69216 14884 69222
rect 14832 69158 14884 69164
rect 14648 69012 14700 69018
rect 14648 68954 14700 68960
rect 14844 68882 14872 69158
rect 14832 68876 14884 68882
rect 14832 68818 14884 68824
rect 14188 68740 14240 68746
rect 14188 68682 14240 68688
rect 14200 68202 14228 68682
rect 14464 68672 14516 68678
rect 14464 68614 14516 68620
rect 14476 68338 14504 68614
rect 14464 68332 14516 68338
rect 14464 68274 14516 68280
rect 14936 68270 14964 70366
rect 15200 68808 15252 68814
rect 15200 68750 15252 68756
rect 15212 68406 15240 68750
rect 15200 68400 15252 68406
rect 15200 68342 15252 68348
rect 14924 68264 14976 68270
rect 14924 68206 14976 68212
rect 14004 68196 14056 68202
rect 14004 68138 14056 68144
rect 14188 68196 14240 68202
rect 14188 68138 14240 68144
rect 14200 67182 14228 68138
rect 15212 67590 15240 68342
rect 15200 67584 15252 67590
rect 15200 67526 15252 67532
rect 14924 67244 14976 67250
rect 14924 67186 14976 67192
rect 14188 67176 14240 67182
rect 14188 67118 14240 67124
rect 14200 66706 14228 67118
rect 14556 67108 14608 67114
rect 14556 67050 14608 67056
rect 14188 66700 14240 66706
rect 14188 66642 14240 66648
rect 14096 66496 14148 66502
rect 14096 66438 14148 66444
rect 14108 66230 14136 66438
rect 14096 66224 14148 66230
rect 14096 66166 14148 66172
rect 14004 65068 14056 65074
rect 14004 65010 14056 65016
rect 14016 63850 14044 65010
rect 14004 63844 14056 63850
rect 14004 63786 14056 63792
rect 13912 63776 13964 63782
rect 13912 63718 13964 63724
rect 13820 63504 13872 63510
rect 13820 63446 13872 63452
rect 13820 63368 13872 63374
rect 13820 63310 13872 63316
rect 13636 60716 13688 60722
rect 13636 60658 13688 60664
rect 13648 60314 13676 60658
rect 13636 60308 13688 60314
rect 13636 60250 13688 60256
rect 13544 59764 13596 59770
rect 13544 59706 13596 59712
rect 13452 59628 13504 59634
rect 13452 59570 13504 59576
rect 13176 58948 13228 58954
rect 13176 58890 13228 58896
rect 13188 58546 13216 58890
rect 13176 58540 13228 58546
rect 13176 58482 13228 58488
rect 12992 57792 13044 57798
rect 12992 57734 13044 57740
rect 10880 57692 11188 57712
rect 10880 57690 10886 57692
rect 10942 57690 10966 57692
rect 11022 57690 11046 57692
rect 11102 57690 11126 57692
rect 11182 57690 11188 57692
rect 10942 57638 10944 57690
rect 11124 57638 11126 57690
rect 10880 57636 10886 57638
rect 10942 57636 10966 57638
rect 11022 57636 11046 57638
rect 11102 57636 11126 57638
rect 11182 57636 11188 57638
rect 10880 57616 11188 57636
rect 2688 57452 2740 57458
rect 2688 57394 2740 57400
rect 2136 57044 2188 57050
rect 2136 56986 2188 56992
rect 2596 56840 2648 56846
rect 2596 56782 2648 56788
rect 1582 56471 1638 56480
rect 1860 56500 1912 56506
rect 1860 56442 1912 56448
rect 2136 56364 2188 56370
rect 2136 56306 2188 56312
rect 2320 56364 2372 56370
rect 2320 56306 2372 56312
rect 1584 56160 1636 56166
rect 1584 56102 1636 56108
rect 1400 55956 1452 55962
rect 1400 55898 1452 55904
rect 1596 55865 1624 56102
rect 1582 55856 1638 55865
rect 1582 55791 1638 55800
rect 1860 55752 1912 55758
rect 1860 55694 1912 55700
rect 1400 55276 1452 55282
rect 1400 55218 1452 55224
rect 1412 54330 1440 55218
rect 1582 55176 1638 55185
rect 1582 55111 1584 55120
rect 1636 55111 1638 55120
rect 1584 55082 1636 55088
rect 1584 54528 1636 54534
rect 1582 54496 1584 54505
rect 1636 54496 1638 54505
rect 1582 54431 1638 54440
rect 1400 54324 1452 54330
rect 1400 54266 1452 54272
rect 1400 54188 1452 54194
rect 1400 54130 1452 54136
rect 1412 53242 1440 54130
rect 1584 53984 1636 53990
rect 1584 53926 1636 53932
rect 1596 53825 1624 53926
rect 1582 53816 1638 53825
rect 1582 53751 1638 53760
rect 1584 53440 1636 53446
rect 1584 53382 1636 53388
rect 1400 53236 1452 53242
rect 1400 53178 1452 53184
rect 1596 53145 1624 53382
rect 1582 53136 1638 53145
rect 1582 53071 1638 53080
rect 1492 52624 1544 52630
rect 1492 52566 1544 52572
rect 1400 51400 1452 51406
rect 1400 51342 1452 51348
rect 1412 50561 1440 51342
rect 1398 50552 1454 50561
rect 1398 50487 1454 50496
rect 1504 50318 1532 52566
rect 1584 52488 1636 52494
rect 1584 52430 1636 52436
rect 1596 51921 1624 52430
rect 1582 51912 1638 51921
rect 1582 51847 1638 51856
rect 1768 51264 1820 51270
rect 1768 51206 1820 51212
rect 1584 50924 1636 50930
rect 1584 50866 1636 50872
rect 1492 50312 1544 50318
rect 1492 50254 1544 50260
rect 1492 50176 1544 50182
rect 1492 50118 1544 50124
rect 1504 49910 1532 50118
rect 1492 49904 1544 49910
rect 1596 49881 1624 50866
rect 1676 50720 1728 50726
rect 1676 50662 1728 50668
rect 1492 49846 1544 49852
rect 1582 49872 1638 49881
rect 1504 49230 1532 49846
rect 1582 49807 1638 49816
rect 1688 49230 1716 50662
rect 1780 49910 1808 51206
rect 1872 50794 1900 55694
rect 2148 55418 2176 56306
rect 2332 55894 2360 56306
rect 2320 55888 2372 55894
rect 2320 55830 2372 55836
rect 2136 55412 2188 55418
rect 2136 55354 2188 55360
rect 2136 54664 2188 54670
rect 2136 54606 2188 54612
rect 2148 53786 2176 54606
rect 2608 54602 2636 56782
rect 2700 55962 2728 57394
rect 5915 57148 6223 57168
rect 5915 57146 5921 57148
rect 5977 57146 6001 57148
rect 6057 57146 6081 57148
rect 6137 57146 6161 57148
rect 6217 57146 6223 57148
rect 5977 57094 5979 57146
rect 6159 57094 6161 57146
rect 5915 57092 5921 57094
rect 5977 57092 6001 57094
rect 6057 57092 6081 57094
rect 6137 57092 6161 57094
rect 6217 57092 6223 57094
rect 5915 57072 6223 57092
rect 10880 56604 11188 56624
rect 10880 56602 10886 56604
rect 10942 56602 10966 56604
rect 11022 56602 11046 56604
rect 11102 56602 11126 56604
rect 11182 56602 11188 56604
rect 10942 56550 10944 56602
rect 11124 56550 11126 56602
rect 10880 56548 10886 56550
rect 10942 56548 10966 56550
rect 11022 56548 11046 56550
rect 11102 56548 11126 56550
rect 11182 56548 11188 56550
rect 10880 56528 11188 56548
rect 5915 56060 6223 56080
rect 5915 56058 5921 56060
rect 5977 56058 6001 56060
rect 6057 56058 6081 56060
rect 6137 56058 6161 56060
rect 6217 56058 6223 56060
rect 5977 56006 5979 56058
rect 6159 56006 6161 56058
rect 5915 56004 5921 56006
rect 5977 56004 6001 56006
rect 6057 56004 6081 56006
rect 6137 56004 6161 56006
rect 6217 56004 6223 56006
rect 5915 55984 6223 56004
rect 2688 55956 2740 55962
rect 2688 55898 2740 55904
rect 10880 55516 11188 55536
rect 10880 55514 10886 55516
rect 10942 55514 10966 55516
rect 11022 55514 11046 55516
rect 11102 55514 11126 55516
rect 11182 55514 11188 55516
rect 10942 55462 10944 55514
rect 11124 55462 11126 55514
rect 10880 55460 10886 55462
rect 10942 55460 10966 55462
rect 11022 55460 11046 55462
rect 11102 55460 11126 55462
rect 11182 55460 11188 55462
rect 10880 55440 11188 55460
rect 9494 55312 9550 55321
rect 4804 55276 4856 55282
rect 9494 55247 9550 55256
rect 4804 55218 4856 55224
rect 2596 54596 2648 54602
rect 2596 54538 2648 54544
rect 2136 53780 2188 53786
rect 2136 53722 2188 53728
rect 2228 53576 2280 53582
rect 2228 53518 2280 53524
rect 2240 53242 2268 53518
rect 2228 53236 2280 53242
rect 2228 53178 2280 53184
rect 1952 53100 2004 53106
rect 1952 53042 2004 53048
rect 1860 50788 1912 50794
rect 1860 50730 1912 50736
rect 1860 50244 1912 50250
rect 1860 50186 1912 50192
rect 1768 49904 1820 49910
rect 1768 49846 1820 49852
rect 1492 49224 1544 49230
rect 1492 49166 1544 49172
rect 1676 49224 1728 49230
rect 1676 49166 1728 49172
rect 1504 48822 1532 49166
rect 1492 48816 1544 48822
rect 1492 48758 1544 48764
rect 1504 48346 1532 48758
rect 1492 48340 1544 48346
rect 1492 48282 1544 48288
rect 1768 48000 1820 48006
rect 1768 47942 1820 47948
rect 1780 47802 1808 47942
rect 1768 47796 1820 47802
rect 1768 47738 1820 47744
rect 1584 47660 1636 47666
rect 1584 47602 1636 47608
rect 1596 47297 1624 47602
rect 1582 47288 1638 47297
rect 1582 47223 1638 47232
rect 1584 47048 1636 47054
rect 1584 46990 1636 46996
rect 1596 46617 1624 46990
rect 1582 46608 1638 46617
rect 1400 46572 1452 46578
rect 1582 46543 1638 46552
rect 1400 46514 1452 46520
rect 1412 45937 1440 46514
rect 1492 45960 1544 45966
rect 1398 45928 1454 45937
rect 1492 45902 1544 45908
rect 1398 45863 1454 45872
rect 1400 45824 1452 45830
rect 1400 45766 1452 45772
rect 1412 44878 1440 45766
rect 1504 45257 1532 45902
rect 1584 45484 1636 45490
rect 1584 45426 1636 45432
rect 1490 45248 1546 45257
rect 1490 45183 1546 45192
rect 1400 44872 1452 44878
rect 1400 44814 1452 44820
rect 1596 44577 1624 45426
rect 1768 45280 1820 45286
rect 1768 45222 1820 45228
rect 1676 44804 1728 44810
rect 1676 44746 1728 44752
rect 1582 44568 1638 44577
rect 1582 44503 1638 44512
rect 1688 44470 1716 44746
rect 1676 44464 1728 44470
rect 1676 44406 1728 44412
rect 1688 43722 1716 44406
rect 1780 43790 1808 45222
rect 1768 43784 1820 43790
rect 1768 43726 1820 43732
rect 1676 43716 1728 43722
rect 1676 43658 1728 43664
rect 1688 43382 1716 43658
rect 1676 43376 1728 43382
rect 1676 43318 1728 43324
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 1780 42906 1808 43250
rect 1768 42900 1820 42906
rect 1768 42842 1820 42848
rect 1584 42696 1636 42702
rect 1582 42664 1584 42673
rect 1636 42664 1638 42673
rect 1582 42599 1638 42608
rect 1584 42220 1636 42226
rect 1584 42162 1636 42168
rect 1596 41993 1624 42162
rect 1582 41984 1638 41993
rect 1582 41919 1638 41928
rect 1584 41608 1636 41614
rect 1584 41550 1636 41556
rect 1596 41313 1624 41550
rect 1582 41304 1638 41313
rect 1582 41239 1638 41248
rect 1872 41206 1900 50186
rect 1964 48634 1992 53042
rect 2044 52624 2096 52630
rect 2044 52566 2096 52572
rect 2056 52465 2084 52566
rect 2872 52556 2924 52562
rect 2872 52498 2924 52504
rect 2228 52488 2280 52494
rect 2042 52456 2098 52465
rect 2228 52430 2280 52436
rect 2042 52391 2098 52400
rect 2240 52154 2268 52430
rect 2228 52148 2280 52154
rect 2228 52090 2280 52096
rect 2228 51400 2280 51406
rect 2228 51342 2280 51348
rect 2044 51264 2096 51270
rect 2240 51241 2268 51342
rect 2044 51206 2096 51212
rect 2226 51232 2282 51241
rect 2056 50318 2084 51206
rect 2226 51167 2282 51176
rect 2688 50516 2740 50522
rect 2688 50458 2740 50464
rect 2044 50312 2096 50318
rect 2044 50254 2096 50260
rect 2504 49768 2556 49774
rect 2504 49710 2556 49716
rect 2136 49632 2188 49638
rect 2136 49574 2188 49580
rect 2148 48822 2176 49574
rect 2320 49156 2372 49162
rect 2320 49098 2372 49104
rect 2136 48816 2188 48822
rect 2136 48758 2188 48764
rect 2332 48754 2360 49098
rect 2320 48748 2372 48754
rect 2320 48690 2372 48696
rect 1964 48606 2176 48634
rect 1952 48544 2004 48550
rect 1952 48486 2004 48492
rect 1964 48346 1992 48486
rect 1952 48340 2004 48346
rect 1952 48282 2004 48288
rect 1952 43648 2004 43654
rect 1952 43590 2004 43596
rect 1964 43382 1992 43590
rect 1952 43376 2004 43382
rect 1952 43318 2004 43324
rect 1860 41200 1912 41206
rect 1860 41142 1912 41148
rect 1584 41132 1636 41138
rect 1584 41074 1636 41080
rect 1596 40633 1624 41074
rect 1582 40624 1638 40633
rect 1582 40559 1638 40568
rect 1584 40044 1636 40050
rect 1584 39986 1636 39992
rect 1596 39953 1624 39986
rect 1582 39944 1638 39953
rect 1582 39879 1638 39888
rect 1584 39432 1636 39438
rect 1584 39374 1636 39380
rect 1596 39273 1624 39374
rect 1582 39264 1638 39273
rect 1582 39199 1638 39208
rect 1584 38956 1636 38962
rect 1584 38898 1636 38904
rect 1596 38593 1624 38898
rect 1582 38584 1638 38593
rect 1582 38519 1638 38528
rect 1584 38344 1636 38350
rect 1584 38286 1636 38292
rect 1596 37913 1624 38286
rect 1582 37904 1638 37913
rect 1400 37868 1452 37874
rect 1582 37839 1638 37848
rect 1400 37810 1452 37816
rect 1412 37369 1440 37810
rect 1398 37360 1454 37369
rect 1398 37295 1454 37304
rect 1584 36780 1636 36786
rect 1584 36722 1636 36728
rect 1596 36689 1624 36722
rect 1582 36680 1638 36689
rect 1582 36615 1638 36624
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1596 36009 1624 36110
rect 1582 36000 1638 36009
rect 1582 35935 1638 35944
rect 2148 35894 2176 48606
rect 2332 48074 2360 48690
rect 2412 48136 2464 48142
rect 2412 48078 2464 48084
rect 2320 48068 2372 48074
rect 2320 48010 2372 48016
rect 2226 47832 2282 47841
rect 2226 47767 2282 47776
rect 2240 47666 2268 47767
rect 2228 47660 2280 47666
rect 2228 47602 2280 47608
rect 2332 46918 2360 48010
rect 2424 47054 2452 48078
rect 2516 47734 2544 49710
rect 2596 48748 2648 48754
rect 2596 48690 2648 48696
rect 2608 47802 2636 48690
rect 2596 47796 2648 47802
rect 2596 47738 2648 47744
rect 2504 47728 2556 47734
rect 2700 47682 2728 50458
rect 2780 49836 2832 49842
rect 2780 49778 2832 49784
rect 2792 49201 2820 49778
rect 2778 49192 2834 49201
rect 2778 49127 2834 49136
rect 2884 48278 2912 52498
rect 3240 49156 3292 49162
rect 3240 49098 3292 49104
rect 3252 48890 3280 49098
rect 3240 48884 3292 48890
rect 3240 48826 3292 48832
rect 3424 48748 3476 48754
rect 3424 48690 3476 48696
rect 3436 48521 3464 48690
rect 3422 48512 3478 48521
rect 3422 48447 3478 48456
rect 2872 48272 2924 48278
rect 2872 48214 2924 48220
rect 2504 47670 2556 47676
rect 2608 47654 2728 47682
rect 2412 47048 2464 47054
rect 2412 46990 2464 46996
rect 2228 46912 2280 46918
rect 2228 46854 2280 46860
rect 2320 46912 2372 46918
rect 2320 46854 2372 46860
rect 2240 45966 2268 46854
rect 2228 45960 2280 45966
rect 2228 45902 2280 45908
rect 2332 45898 2360 46854
rect 2424 46458 2452 46990
rect 2424 46430 2544 46458
rect 2412 46368 2464 46374
rect 2412 46310 2464 46316
rect 2320 45892 2372 45898
rect 2320 45834 2372 45840
rect 2228 45824 2280 45830
rect 2228 45766 2280 45772
rect 2240 43314 2268 45766
rect 2332 45558 2360 45834
rect 2424 45558 2452 46310
rect 2516 45830 2544 46430
rect 2504 45824 2556 45830
rect 2504 45766 2556 45772
rect 2320 45552 2372 45558
rect 2320 45494 2372 45500
rect 2412 45552 2464 45558
rect 2412 45494 2464 45500
rect 2608 44538 2636 47654
rect 2688 45824 2740 45830
rect 2688 45766 2740 45772
rect 2700 45626 2728 45766
rect 2688 45620 2740 45626
rect 2688 45562 2740 45568
rect 2596 44532 2648 44538
rect 2596 44474 2648 44480
rect 2780 44396 2832 44402
rect 2780 44338 2832 44344
rect 2792 43897 2820 44338
rect 2778 43888 2834 43897
rect 2778 43823 2834 43832
rect 2596 43716 2648 43722
rect 2596 43658 2648 43664
rect 2228 43308 2280 43314
rect 2228 43250 2280 43256
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 2226 43208 2282 43217
rect 2226 43143 2282 43152
rect 2240 42702 2268 43143
rect 2228 42696 2280 42702
rect 2228 42638 2280 42644
rect 2516 37466 2544 43250
rect 2608 42906 2636 43658
rect 2596 42900 2648 42906
rect 2596 42842 2648 42848
rect 2504 37460 2556 37466
rect 2504 37402 2556 37408
rect 2148 35866 2268 35894
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35329 1624 35634
rect 1582 35320 1638 35329
rect 1582 35255 1638 35264
rect 1584 35080 1636 35086
rect 1584 35022 1636 35028
rect 1596 34649 1624 35022
rect 1582 34640 1638 34649
rect 1400 34604 1452 34610
rect 1582 34575 1638 34584
rect 1400 34546 1452 34552
rect 1412 33969 1440 34546
rect 1584 33992 1636 33998
rect 1398 33960 1454 33969
rect 1584 33934 1636 33940
rect 1398 33895 1454 33904
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1412 32745 1440 33458
rect 1596 33289 1624 33934
rect 1582 33280 1638 33289
rect 1582 33215 1638 33224
rect 1492 32904 1544 32910
rect 1492 32846 1544 32852
rect 1398 32736 1454 32745
rect 1398 32671 1454 32680
rect 1504 32065 1532 32846
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1490 32056 1546 32065
rect 1490 31991 1546 32000
rect 1596 31385 1624 32370
rect 1858 31920 1914 31929
rect 1858 31855 1914 31864
rect 1872 31822 1900 31855
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 1676 31680 1728 31686
rect 1676 31622 1728 31628
rect 1582 31376 1638 31385
rect 1582 31311 1638 31320
rect 1400 31136 1452 31142
rect 1400 31078 1452 31084
rect 1412 27470 1440 31078
rect 1582 30696 1638 30705
rect 1582 30631 1638 30640
rect 1596 30598 1624 30631
rect 1584 30592 1636 30598
rect 1584 30534 1636 30540
rect 1688 30258 1716 31622
rect 1860 31340 1912 31346
rect 1860 31282 1912 31288
rect 1872 30870 1900 31282
rect 1860 30864 1912 30870
rect 1860 30806 1912 30812
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1676 30252 1728 30258
rect 1676 30194 1728 30200
rect 1584 30048 1636 30054
rect 1582 30016 1584 30025
rect 1676 30048 1728 30054
rect 1636 30016 1638 30025
rect 1676 29990 1728 29996
rect 1582 29951 1638 29960
rect 1584 29504 1636 29510
rect 1584 29446 1636 29452
rect 1596 29345 1624 29446
rect 1582 29336 1638 29345
rect 1582 29271 1638 29280
rect 1688 29170 1716 29990
rect 1676 29164 1728 29170
rect 1676 29106 1728 29112
rect 1584 29028 1636 29034
rect 1584 28970 1636 28976
rect 1596 28665 1624 28970
rect 1582 28656 1638 28665
rect 1582 28591 1638 28600
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 1596 28121 1624 28358
rect 1582 28112 1638 28121
rect 1582 28047 1638 28056
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 1596 27334 1624 27367
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1584 26784 1636 26790
rect 1582 26752 1584 26761
rect 1636 26752 1638 26761
rect 1582 26687 1638 26696
rect 1584 26240 1636 26246
rect 1780 26234 1808 30670
rect 2136 30592 2188 30598
rect 2136 30534 2188 30540
rect 2148 29646 2176 30534
rect 2136 29640 2188 29646
rect 2136 29582 2188 29588
rect 2136 29504 2188 29510
rect 2136 29446 2188 29452
rect 2148 28558 2176 29446
rect 2136 28552 2188 28558
rect 2136 28494 2188 28500
rect 2240 28490 2268 35866
rect 2320 32224 2372 32230
rect 2320 32166 2372 32172
rect 2332 31346 2360 32166
rect 2516 31822 2544 37402
rect 3976 35488 4028 35494
rect 3976 35430 4028 35436
rect 2596 32768 2648 32774
rect 2596 32710 2648 32716
rect 2608 31822 2636 32710
rect 2504 31816 2556 31822
rect 2504 31758 2556 31764
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2516 31414 2544 31758
rect 3988 31414 4016 35430
rect 4068 34944 4120 34950
rect 4068 34886 4120 34892
rect 4080 31482 4108 34886
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 2504 31408 2556 31414
rect 2504 31350 2556 31356
rect 3976 31408 4028 31414
rect 3976 31350 4028 31356
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 4068 30728 4120 30734
rect 4068 30670 4120 30676
rect 4080 29850 4108 30670
rect 4068 29844 4120 29850
rect 4068 29786 4120 29792
rect 2228 28484 2280 28490
rect 2228 28426 2280 28432
rect 2320 27124 2372 27130
rect 2320 27066 2372 27072
rect 2332 26382 2360 27066
rect 2320 26376 2372 26382
rect 2320 26318 2372 26324
rect 1584 26182 1636 26188
rect 1688 26206 1808 26234
rect 1596 26081 1624 26182
rect 1582 26072 1638 26081
rect 1582 26007 1638 26016
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25401 1624 25638
rect 1688 25498 1716 26206
rect 1676 25492 1728 25498
rect 1676 25434 1728 25440
rect 2320 25492 2372 25498
rect 2320 25434 2372 25440
rect 1582 25392 1638 25401
rect 1582 25327 1638 25336
rect 1860 25288 1912 25294
rect 1860 25230 1912 25236
rect 1872 24886 1900 25230
rect 1860 24880 1912 24886
rect 1860 24822 1912 24828
rect 2332 24818 2360 25434
rect 2320 24812 2372 24818
rect 2320 24754 2372 24760
rect 1582 24712 1638 24721
rect 1582 24647 1584 24656
rect 1636 24647 1638 24656
rect 1584 24618 1636 24624
rect 1584 24064 1636 24070
rect 1582 24032 1584 24041
rect 1636 24032 1638 24041
rect 1582 23967 1638 23976
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1596 22817 1624 22918
rect 1582 22808 1638 22817
rect 2332 22778 2360 23054
rect 1582 22743 1638 22752
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22137 1624 22374
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 1400 21888 1452 21894
rect 1400 21830 1452 21836
rect 1412 21554 1440 21830
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1582 21448 1638 21457
rect 1582 21383 1584 21392
rect 1636 21383 1638 21392
rect 1584 21354 1636 21360
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1412 20942 1440 21286
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1584 20800 1636 20806
rect 1582 20768 1584 20777
rect 1636 20768 1638 20777
rect 1582 20703 1638 20712
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20097 1624 20198
rect 1582 20088 1638 20097
rect 2148 20058 2176 20402
rect 1582 20023 1638 20032
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2332 19854 2360 20538
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2320 19848 2372 19854
rect 2320 19790 2372 19796
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1596 19417 1624 19654
rect 2148 19514 2176 19790
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 1582 19408 1638 19417
rect 1400 19372 1452 19378
rect 1582 19343 1638 19352
rect 1400 19314 1452 19320
rect 1412 18970 1440 19314
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1596 18873 1624 19110
rect 1582 18864 1638 18873
rect 1582 18799 1638 18808
rect 1492 18692 1544 18698
rect 1492 18634 1544 18640
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1412 18290 1440 18566
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17678 1440 18022
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15026 1440 15846
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1412 13938 1440 14554
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11354 1440 11698
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1504 3058 1532 18634
rect 1582 18184 1638 18193
rect 1582 18119 1584 18128
rect 1636 18119 1638 18128
rect 1584 18090 1636 18096
rect 1584 17536 1636 17542
rect 1582 17504 1584 17513
rect 1636 17504 1638 17513
rect 1582 17439 1638 17448
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16833 1624 16934
rect 1582 16824 1638 16833
rect 1582 16759 1638 16768
rect 2700 16522 2728 17138
rect 2688 16516 2740 16522
rect 2688 16458 2740 16464
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16153 1624 16390
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15502 1808 15846
rect 1768 15496 1820 15502
rect 1582 15464 1638 15473
rect 1768 15438 1820 15444
rect 1582 15399 1638 15408
rect 1596 15366 1624 15399
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 1584 14816 1636 14822
rect 1582 14784 1584 14793
rect 1636 14784 1638 14793
rect 1582 14719 1638 14728
rect 2148 14414 2176 15302
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1584 14272 1636 14278
rect 1582 14240 1584 14249
rect 1636 14240 1638 14249
rect 1582 14175 1638 14184
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13569 1624 13670
rect 1582 13560 1638 13569
rect 1582 13495 1638 13504
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12889 1624 13126
rect 2044 12912 2096 12918
rect 1582 12880 1638 12889
rect 2044 12854 2096 12860
rect 1582 12815 1638 12824
rect 2056 12442 2084 12854
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 2056 12238 2084 12378
rect 2044 12232 2096 12238
rect 1582 12200 1638 12209
rect 2044 12174 2096 12180
rect 1582 12135 1638 12144
rect 1596 12102 1624 12135
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1584 11552 1636 11558
rect 1582 11520 1584 11529
rect 1636 11520 1638 11529
rect 1582 11455 1638 11464
rect 2332 11150 2360 12650
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 1596 10849 1624 10950
rect 1582 10840 1638 10849
rect 1582 10775 1638 10784
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10169 1624 10406
rect 1582 10160 1638 10169
rect 1582 10095 1638 10104
rect 2148 10062 2176 10950
rect 2700 10062 2728 12174
rect 4816 11830 4844 55218
rect 5915 54972 6223 54992
rect 5915 54970 5921 54972
rect 5977 54970 6001 54972
rect 6057 54970 6081 54972
rect 6137 54970 6161 54972
rect 6217 54970 6223 54972
rect 5977 54918 5979 54970
rect 6159 54918 6161 54970
rect 5915 54916 5921 54918
rect 5977 54916 6001 54918
rect 6057 54916 6081 54918
rect 6137 54916 6161 54918
rect 6217 54916 6223 54918
rect 5915 54896 6223 54916
rect 7564 54188 7616 54194
rect 7564 54130 7616 54136
rect 5915 53884 6223 53904
rect 5915 53882 5921 53884
rect 5977 53882 6001 53884
rect 6057 53882 6081 53884
rect 6137 53882 6161 53884
rect 6217 53882 6223 53884
rect 5977 53830 5979 53882
rect 6159 53830 6161 53882
rect 5915 53828 5921 53830
rect 5977 53828 6001 53830
rect 6057 53828 6081 53830
rect 6137 53828 6161 53830
rect 6217 53828 6223 53830
rect 5915 53808 6223 53828
rect 6276 53576 6328 53582
rect 6276 53518 6328 53524
rect 5915 52796 6223 52816
rect 5915 52794 5921 52796
rect 5977 52794 6001 52796
rect 6057 52794 6081 52796
rect 6137 52794 6161 52796
rect 6217 52794 6223 52796
rect 5977 52742 5979 52794
rect 6159 52742 6161 52794
rect 5915 52740 5921 52742
rect 5977 52740 6001 52742
rect 6057 52740 6081 52742
rect 6137 52740 6161 52742
rect 6217 52740 6223 52742
rect 5915 52720 6223 52740
rect 5915 51708 6223 51728
rect 5915 51706 5921 51708
rect 5977 51706 6001 51708
rect 6057 51706 6081 51708
rect 6137 51706 6161 51708
rect 6217 51706 6223 51708
rect 5977 51654 5979 51706
rect 6159 51654 6161 51706
rect 5915 51652 5921 51654
rect 5977 51652 6001 51654
rect 6057 51652 6081 51654
rect 6137 51652 6161 51654
rect 6217 51652 6223 51654
rect 5915 51632 6223 51652
rect 5915 50620 6223 50640
rect 5915 50618 5921 50620
rect 5977 50618 6001 50620
rect 6057 50618 6081 50620
rect 6137 50618 6161 50620
rect 6217 50618 6223 50620
rect 5977 50566 5979 50618
rect 6159 50566 6161 50618
rect 5915 50564 5921 50566
rect 5977 50564 6001 50566
rect 6057 50564 6081 50566
rect 6137 50564 6161 50566
rect 6217 50564 6223 50566
rect 5915 50544 6223 50564
rect 5915 49532 6223 49552
rect 5915 49530 5921 49532
rect 5977 49530 6001 49532
rect 6057 49530 6081 49532
rect 6137 49530 6161 49532
rect 6217 49530 6223 49532
rect 5977 49478 5979 49530
rect 6159 49478 6161 49530
rect 5915 49476 5921 49478
rect 5977 49476 6001 49478
rect 6057 49476 6081 49478
rect 6137 49476 6161 49478
rect 6217 49476 6223 49478
rect 5915 49456 6223 49476
rect 5915 48444 6223 48464
rect 5915 48442 5921 48444
rect 5977 48442 6001 48444
rect 6057 48442 6081 48444
rect 6137 48442 6161 48444
rect 6217 48442 6223 48444
rect 5977 48390 5979 48442
rect 6159 48390 6161 48442
rect 5915 48388 5921 48390
rect 5977 48388 6001 48390
rect 6057 48388 6081 48390
rect 6137 48388 6161 48390
rect 6217 48388 6223 48390
rect 5915 48368 6223 48388
rect 5915 47356 6223 47376
rect 5915 47354 5921 47356
rect 5977 47354 6001 47356
rect 6057 47354 6081 47356
rect 6137 47354 6161 47356
rect 6217 47354 6223 47356
rect 5977 47302 5979 47354
rect 6159 47302 6161 47354
rect 5915 47300 5921 47302
rect 5977 47300 6001 47302
rect 6057 47300 6081 47302
rect 6137 47300 6161 47302
rect 6217 47300 6223 47302
rect 5915 47280 6223 47300
rect 5915 46268 6223 46288
rect 5915 46266 5921 46268
rect 5977 46266 6001 46268
rect 6057 46266 6081 46268
rect 6137 46266 6161 46268
rect 6217 46266 6223 46268
rect 5977 46214 5979 46266
rect 6159 46214 6161 46266
rect 5915 46212 5921 46214
rect 5977 46212 6001 46214
rect 6057 46212 6081 46214
rect 6137 46212 6161 46214
rect 6217 46212 6223 46214
rect 5915 46192 6223 46212
rect 5915 45180 6223 45200
rect 5915 45178 5921 45180
rect 5977 45178 6001 45180
rect 6057 45178 6081 45180
rect 6137 45178 6161 45180
rect 6217 45178 6223 45180
rect 5977 45126 5979 45178
rect 6159 45126 6161 45178
rect 5915 45124 5921 45126
rect 5977 45124 6001 45126
rect 6057 45124 6081 45126
rect 6137 45124 6161 45126
rect 6217 45124 6223 45126
rect 5915 45104 6223 45124
rect 5915 44092 6223 44112
rect 5915 44090 5921 44092
rect 5977 44090 6001 44092
rect 6057 44090 6081 44092
rect 6137 44090 6161 44092
rect 6217 44090 6223 44092
rect 5977 44038 5979 44090
rect 6159 44038 6161 44090
rect 5915 44036 5921 44038
rect 5977 44036 6001 44038
rect 6057 44036 6081 44038
rect 6137 44036 6161 44038
rect 6217 44036 6223 44038
rect 5915 44016 6223 44036
rect 5915 43004 6223 43024
rect 5915 43002 5921 43004
rect 5977 43002 6001 43004
rect 6057 43002 6081 43004
rect 6137 43002 6161 43004
rect 6217 43002 6223 43004
rect 5977 42950 5979 43002
rect 6159 42950 6161 43002
rect 5915 42948 5921 42950
rect 5977 42948 6001 42950
rect 6057 42948 6081 42950
rect 6137 42948 6161 42950
rect 6217 42948 6223 42950
rect 5915 42928 6223 42948
rect 5915 41916 6223 41936
rect 5915 41914 5921 41916
rect 5977 41914 6001 41916
rect 6057 41914 6081 41916
rect 6137 41914 6161 41916
rect 6217 41914 6223 41916
rect 5977 41862 5979 41914
rect 6159 41862 6161 41914
rect 5915 41860 5921 41862
rect 5977 41860 6001 41862
rect 6057 41860 6081 41862
rect 6137 41860 6161 41862
rect 6217 41860 6223 41862
rect 5915 41840 6223 41860
rect 5915 40828 6223 40848
rect 5915 40826 5921 40828
rect 5977 40826 6001 40828
rect 6057 40826 6081 40828
rect 6137 40826 6161 40828
rect 6217 40826 6223 40828
rect 5977 40774 5979 40826
rect 6159 40774 6161 40826
rect 5915 40772 5921 40774
rect 5977 40772 6001 40774
rect 6057 40772 6081 40774
rect 6137 40772 6161 40774
rect 6217 40772 6223 40774
rect 5915 40752 6223 40772
rect 5915 39740 6223 39760
rect 5915 39738 5921 39740
rect 5977 39738 6001 39740
rect 6057 39738 6081 39740
rect 6137 39738 6161 39740
rect 6217 39738 6223 39740
rect 5977 39686 5979 39738
rect 6159 39686 6161 39738
rect 5915 39684 5921 39686
rect 5977 39684 6001 39686
rect 6057 39684 6081 39686
rect 6137 39684 6161 39686
rect 6217 39684 6223 39686
rect 5915 39664 6223 39684
rect 5915 38652 6223 38672
rect 5915 38650 5921 38652
rect 5977 38650 6001 38652
rect 6057 38650 6081 38652
rect 6137 38650 6161 38652
rect 6217 38650 6223 38652
rect 5977 38598 5979 38650
rect 6159 38598 6161 38650
rect 5915 38596 5921 38598
rect 5977 38596 6001 38598
rect 6057 38596 6081 38598
rect 6137 38596 6161 38598
rect 6217 38596 6223 38598
rect 5915 38576 6223 38596
rect 5915 37564 6223 37584
rect 5915 37562 5921 37564
rect 5977 37562 6001 37564
rect 6057 37562 6081 37564
rect 6137 37562 6161 37564
rect 6217 37562 6223 37564
rect 5977 37510 5979 37562
rect 6159 37510 6161 37562
rect 5915 37508 5921 37510
rect 5977 37508 6001 37510
rect 6057 37508 6081 37510
rect 6137 37508 6161 37510
rect 6217 37508 6223 37510
rect 5915 37488 6223 37508
rect 5915 36476 6223 36496
rect 5915 36474 5921 36476
rect 5977 36474 6001 36476
rect 6057 36474 6081 36476
rect 6137 36474 6161 36476
rect 6217 36474 6223 36476
rect 5977 36422 5979 36474
rect 6159 36422 6161 36474
rect 5915 36420 5921 36422
rect 5977 36420 6001 36422
rect 6057 36420 6081 36422
rect 6137 36420 6161 36422
rect 6217 36420 6223 36422
rect 5915 36400 6223 36420
rect 5915 35388 6223 35408
rect 5915 35386 5921 35388
rect 5977 35386 6001 35388
rect 6057 35386 6081 35388
rect 6137 35386 6161 35388
rect 6217 35386 6223 35388
rect 5977 35334 5979 35386
rect 6159 35334 6161 35386
rect 5915 35332 5921 35334
rect 5977 35332 6001 35334
rect 6057 35332 6081 35334
rect 6137 35332 6161 35334
rect 6217 35332 6223 35334
rect 5915 35312 6223 35332
rect 5915 34300 6223 34320
rect 5915 34298 5921 34300
rect 5977 34298 6001 34300
rect 6057 34298 6081 34300
rect 6137 34298 6161 34300
rect 6217 34298 6223 34300
rect 5977 34246 5979 34298
rect 6159 34246 6161 34298
rect 5915 34244 5921 34246
rect 5977 34244 6001 34246
rect 6057 34244 6081 34246
rect 6137 34244 6161 34246
rect 6217 34244 6223 34246
rect 5915 34224 6223 34244
rect 5915 33212 6223 33232
rect 5915 33210 5921 33212
rect 5977 33210 6001 33212
rect 6057 33210 6081 33212
rect 6137 33210 6161 33212
rect 6217 33210 6223 33212
rect 5977 33158 5979 33210
rect 6159 33158 6161 33210
rect 5915 33156 5921 33158
rect 5977 33156 6001 33158
rect 6057 33156 6081 33158
rect 6137 33156 6161 33158
rect 6217 33156 6223 33158
rect 5915 33136 6223 33156
rect 5915 32124 6223 32144
rect 5915 32122 5921 32124
rect 5977 32122 6001 32124
rect 6057 32122 6081 32124
rect 6137 32122 6161 32124
rect 6217 32122 6223 32124
rect 5977 32070 5979 32122
rect 6159 32070 6161 32122
rect 5915 32068 5921 32070
rect 5977 32068 6001 32070
rect 6057 32068 6081 32070
rect 6137 32068 6161 32070
rect 6217 32068 6223 32070
rect 5915 32048 6223 32068
rect 5915 31036 6223 31056
rect 5915 31034 5921 31036
rect 5977 31034 6001 31036
rect 6057 31034 6081 31036
rect 6137 31034 6161 31036
rect 6217 31034 6223 31036
rect 5977 30982 5979 31034
rect 6159 30982 6161 31034
rect 5915 30980 5921 30982
rect 5977 30980 6001 30982
rect 6057 30980 6081 30982
rect 6137 30980 6161 30982
rect 6217 30980 6223 30982
rect 5915 30960 6223 30980
rect 5915 29948 6223 29968
rect 5915 29946 5921 29948
rect 5977 29946 6001 29948
rect 6057 29946 6081 29948
rect 6137 29946 6161 29948
rect 6217 29946 6223 29948
rect 5977 29894 5979 29946
rect 6159 29894 6161 29946
rect 5915 29892 5921 29894
rect 5977 29892 6001 29894
rect 6057 29892 6081 29894
rect 6137 29892 6161 29894
rect 6217 29892 6223 29894
rect 5915 29872 6223 29892
rect 5915 28860 6223 28880
rect 5915 28858 5921 28860
rect 5977 28858 6001 28860
rect 6057 28858 6081 28860
rect 6137 28858 6161 28860
rect 6217 28858 6223 28860
rect 5977 28806 5979 28858
rect 6159 28806 6161 28858
rect 5915 28804 5921 28806
rect 5977 28804 6001 28806
rect 6057 28804 6081 28806
rect 6137 28804 6161 28806
rect 6217 28804 6223 28806
rect 5915 28784 6223 28804
rect 5915 27772 6223 27792
rect 5915 27770 5921 27772
rect 5977 27770 6001 27772
rect 6057 27770 6081 27772
rect 6137 27770 6161 27772
rect 6217 27770 6223 27772
rect 5977 27718 5979 27770
rect 6159 27718 6161 27770
rect 5915 27716 5921 27718
rect 5977 27716 6001 27718
rect 6057 27716 6081 27718
rect 6137 27716 6161 27718
rect 6217 27716 6223 27718
rect 5915 27696 6223 27716
rect 5915 26684 6223 26704
rect 5915 26682 5921 26684
rect 5977 26682 6001 26684
rect 6057 26682 6081 26684
rect 6137 26682 6161 26684
rect 6217 26682 6223 26684
rect 5977 26630 5979 26682
rect 6159 26630 6161 26682
rect 5915 26628 5921 26630
rect 5977 26628 6001 26630
rect 6057 26628 6081 26630
rect 6137 26628 6161 26630
rect 6217 26628 6223 26630
rect 5915 26608 6223 26628
rect 5915 25596 6223 25616
rect 5915 25594 5921 25596
rect 5977 25594 6001 25596
rect 6057 25594 6081 25596
rect 6137 25594 6161 25596
rect 6217 25594 6223 25596
rect 5977 25542 5979 25594
rect 6159 25542 6161 25594
rect 5915 25540 5921 25542
rect 5977 25540 6001 25542
rect 6057 25540 6081 25542
rect 6137 25540 6161 25542
rect 6217 25540 6223 25542
rect 5915 25520 6223 25540
rect 5915 24508 6223 24528
rect 5915 24506 5921 24508
rect 5977 24506 6001 24508
rect 6057 24506 6081 24508
rect 6137 24506 6161 24508
rect 6217 24506 6223 24508
rect 5977 24454 5979 24506
rect 6159 24454 6161 24506
rect 5915 24452 5921 24454
rect 5977 24452 6001 24454
rect 6057 24452 6081 24454
rect 6137 24452 6161 24454
rect 6217 24452 6223 24454
rect 5915 24432 6223 24452
rect 5915 23420 6223 23440
rect 5915 23418 5921 23420
rect 5977 23418 6001 23420
rect 6057 23418 6081 23420
rect 6137 23418 6161 23420
rect 6217 23418 6223 23420
rect 5977 23366 5979 23418
rect 6159 23366 6161 23418
rect 5915 23364 5921 23366
rect 5977 23364 6001 23366
rect 6057 23364 6081 23366
rect 6137 23364 6161 23366
rect 6217 23364 6223 23366
rect 5915 23344 6223 23364
rect 5915 22332 6223 22352
rect 5915 22330 5921 22332
rect 5977 22330 6001 22332
rect 6057 22330 6081 22332
rect 6137 22330 6161 22332
rect 6217 22330 6223 22332
rect 5977 22278 5979 22330
rect 6159 22278 6161 22330
rect 5915 22276 5921 22278
rect 5977 22276 6001 22278
rect 6057 22276 6081 22278
rect 6137 22276 6161 22278
rect 6217 22276 6223 22278
rect 5915 22256 6223 22276
rect 5915 21244 6223 21264
rect 5915 21242 5921 21244
rect 5977 21242 6001 21244
rect 6057 21242 6081 21244
rect 6137 21242 6161 21244
rect 6217 21242 6223 21244
rect 5977 21190 5979 21242
rect 6159 21190 6161 21242
rect 5915 21188 5921 21190
rect 5977 21188 6001 21190
rect 6057 21188 6081 21190
rect 6137 21188 6161 21190
rect 6217 21188 6223 21190
rect 5915 21168 6223 21188
rect 5915 20156 6223 20176
rect 5915 20154 5921 20156
rect 5977 20154 6001 20156
rect 6057 20154 6081 20156
rect 6137 20154 6161 20156
rect 6217 20154 6223 20156
rect 5977 20102 5979 20154
rect 6159 20102 6161 20154
rect 5915 20100 5921 20102
rect 5977 20100 6001 20102
rect 6057 20100 6081 20102
rect 6137 20100 6161 20102
rect 6217 20100 6223 20102
rect 5915 20080 6223 20100
rect 5915 19068 6223 19088
rect 5915 19066 5921 19068
rect 5977 19066 6001 19068
rect 6057 19066 6081 19068
rect 6137 19066 6161 19068
rect 6217 19066 6223 19068
rect 5977 19014 5979 19066
rect 6159 19014 6161 19066
rect 5915 19012 5921 19014
rect 5977 19012 6001 19014
rect 6057 19012 6081 19014
rect 6137 19012 6161 19014
rect 6217 19012 6223 19014
rect 5915 18992 6223 19012
rect 5915 17980 6223 18000
rect 5915 17978 5921 17980
rect 5977 17978 6001 17980
rect 6057 17978 6081 17980
rect 6137 17978 6161 17980
rect 6217 17978 6223 17980
rect 5977 17926 5979 17978
rect 6159 17926 6161 17978
rect 5915 17924 5921 17926
rect 5977 17924 6001 17926
rect 6057 17924 6081 17926
rect 6137 17924 6161 17926
rect 6217 17924 6223 17926
rect 5915 17904 6223 17924
rect 5915 16892 6223 16912
rect 5915 16890 5921 16892
rect 5977 16890 6001 16892
rect 6057 16890 6081 16892
rect 6137 16890 6161 16892
rect 6217 16890 6223 16892
rect 5977 16838 5979 16890
rect 6159 16838 6161 16890
rect 5915 16836 5921 16838
rect 5977 16836 6001 16838
rect 6057 16836 6081 16838
rect 6137 16836 6161 16838
rect 6217 16836 6223 16838
rect 5915 16816 6223 16836
rect 6288 16574 6316 53518
rect 7472 45348 7524 45354
rect 7472 45290 7524 45296
rect 7484 45082 7512 45290
rect 7472 45076 7524 45082
rect 7472 45018 7524 45024
rect 6288 16546 6408 16574
rect 5915 15804 6223 15824
rect 5915 15802 5921 15804
rect 5977 15802 6001 15804
rect 6057 15802 6081 15804
rect 6137 15802 6161 15804
rect 6217 15802 6223 15804
rect 5977 15750 5979 15802
rect 6159 15750 6161 15802
rect 5915 15748 5921 15750
rect 5977 15748 6001 15750
rect 6057 15748 6081 15750
rect 6137 15748 6161 15750
rect 6217 15748 6223 15750
rect 5915 15728 6223 15748
rect 5915 14716 6223 14736
rect 5915 14714 5921 14716
rect 5977 14714 6001 14716
rect 6057 14714 6081 14716
rect 6137 14714 6161 14716
rect 6217 14714 6223 14716
rect 5977 14662 5979 14714
rect 6159 14662 6161 14714
rect 5915 14660 5921 14662
rect 5977 14660 6001 14662
rect 6057 14660 6081 14662
rect 6137 14660 6161 14662
rect 6217 14660 6223 14662
rect 5915 14640 6223 14660
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 5915 13628 6223 13648
rect 5915 13626 5921 13628
rect 5977 13626 6001 13628
rect 6057 13626 6081 13628
rect 6137 13626 6161 13628
rect 6217 13626 6223 13628
rect 5977 13574 5979 13626
rect 6159 13574 6161 13626
rect 5915 13572 5921 13574
rect 5977 13572 6001 13574
rect 6057 13572 6081 13574
rect 6137 13572 6161 13574
rect 6217 13572 6223 13574
rect 5915 13552 6223 13572
rect 5915 12540 6223 12560
rect 5915 12538 5921 12540
rect 5977 12538 6001 12540
rect 6057 12538 6081 12540
rect 6137 12538 6161 12540
rect 6217 12538 6223 12540
rect 5977 12486 5979 12538
rect 6159 12486 6161 12538
rect 5915 12484 5921 12486
rect 5977 12484 6001 12486
rect 6057 12484 6081 12486
rect 6137 12484 6161 12486
rect 6217 12484 6223 12486
rect 5915 12464 6223 12484
rect 6288 12238 6316 14486
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 5915 11452 6223 11472
rect 5915 11450 5921 11452
rect 5977 11450 6001 11452
rect 6057 11450 6081 11452
rect 6137 11450 6161 11452
rect 6217 11450 6223 11452
rect 5977 11398 5979 11450
rect 6159 11398 6161 11450
rect 5915 11396 5921 11398
rect 5977 11396 6001 11398
rect 6057 11396 6081 11398
rect 6137 11396 6161 11398
rect 6217 11396 6223 11398
rect 5915 11376 6223 11396
rect 5915 10364 6223 10384
rect 5915 10362 5921 10364
rect 5977 10362 6001 10364
rect 6057 10362 6081 10364
rect 6137 10362 6161 10364
rect 6217 10362 6223 10364
rect 5977 10310 5979 10362
rect 6159 10310 6161 10362
rect 5915 10308 5921 10310
rect 5977 10308 6001 10310
rect 6057 10308 6081 10310
rect 6137 10308 6161 10310
rect 6217 10308 6223 10310
rect 5915 10288 6223 10308
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 1596 9625 1624 9862
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 2148 8974 2176 9862
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2332 8974 2360 9386
rect 5915 9276 6223 9296
rect 5915 9274 5921 9276
rect 5977 9274 6001 9276
rect 6057 9274 6081 9276
rect 6137 9274 6161 9276
rect 6217 9274 6223 9276
rect 5977 9222 5979 9274
rect 6159 9222 6161 9274
rect 5915 9220 5921 9222
rect 5977 9220 6001 9222
rect 6057 9220 6081 9222
rect 6137 9220 6161 9222
rect 6217 9220 6223 9222
rect 5915 9200 6223 9220
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2136 8968 2188 8974
rect 1582 8936 1638 8945
rect 2136 8910 2188 8916
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 1582 8871 1638 8880
rect 1596 8838 1624 8871
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 8498 2176 8774
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 8265 1624 8298
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 2700 7886 2728 9114
rect 5915 8188 6223 8208
rect 5915 8186 5921 8188
rect 5977 8186 6001 8188
rect 6057 8186 6081 8188
rect 6137 8186 6161 8188
rect 6217 8186 6223 8188
rect 5977 8134 5979 8186
rect 6159 8134 6161 8186
rect 5915 8132 5921 8134
rect 5977 8132 6001 8134
rect 6057 8132 6081 8134
rect 6137 8132 6161 8134
rect 6217 8132 6223 8134
rect 5915 8112 6223 8132
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7585 1624 7686
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 2056 6458 2084 7482
rect 6380 7478 6408 16546
rect 7576 9654 7604 54130
rect 9402 43752 9458 43761
rect 9402 43687 9458 43696
rect 9416 43382 9444 43687
rect 9404 43376 9456 43382
rect 9404 43318 9456 43324
rect 8392 42220 8444 42226
rect 8392 42162 8444 42168
rect 8404 41614 8432 42162
rect 8392 41608 8444 41614
rect 8392 41550 8444 41556
rect 8208 40928 8260 40934
rect 8208 40870 8260 40876
rect 8220 40526 8248 40870
rect 8404 40594 8432 41550
rect 8668 40724 8720 40730
rect 8668 40666 8720 40672
rect 8392 40588 8444 40594
rect 8392 40530 8444 40536
rect 8208 40520 8260 40526
rect 8208 40462 8260 40468
rect 8404 40050 8432 40530
rect 8680 40186 8708 40666
rect 8668 40180 8720 40186
rect 8668 40122 8720 40128
rect 8392 40044 8444 40050
rect 8392 39986 8444 39992
rect 8404 39030 8432 39986
rect 8576 39296 8628 39302
rect 8576 39238 8628 39244
rect 8588 39030 8616 39238
rect 8392 39024 8444 39030
rect 8392 38966 8444 38972
rect 8576 39024 8628 39030
rect 8576 38966 8628 38972
rect 8404 38010 8432 38966
rect 9036 38820 9088 38826
rect 9036 38762 9088 38768
rect 8392 38004 8444 38010
rect 8392 37946 8444 37952
rect 9048 37942 9076 38762
rect 9036 37936 9088 37942
rect 9036 37878 9088 37884
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 8220 36378 8248 37198
rect 8312 37194 8340 37810
rect 9128 37664 9180 37670
rect 9128 37606 9180 37612
rect 8300 37188 8352 37194
rect 8300 37130 8352 37136
rect 8208 36372 8260 36378
rect 8208 36314 8260 36320
rect 8312 36174 8340 37130
rect 9140 36854 9168 37606
rect 9128 36848 9180 36854
rect 9508 36825 9536 55247
rect 13360 54800 13412 54806
rect 13360 54742 13412 54748
rect 10880 54428 11188 54448
rect 10880 54426 10886 54428
rect 10942 54426 10966 54428
rect 11022 54426 11046 54428
rect 11102 54426 11126 54428
rect 11182 54426 11188 54428
rect 10942 54374 10944 54426
rect 11124 54374 11126 54426
rect 10880 54372 10886 54374
rect 10942 54372 10966 54374
rect 11022 54372 11046 54374
rect 11102 54372 11126 54374
rect 11182 54372 11188 54374
rect 10880 54352 11188 54372
rect 10880 53340 11188 53360
rect 10880 53338 10886 53340
rect 10942 53338 10966 53340
rect 11022 53338 11046 53340
rect 11102 53338 11126 53340
rect 11182 53338 11188 53340
rect 10942 53286 10944 53338
rect 11124 53286 11126 53338
rect 10880 53284 10886 53286
rect 10942 53284 10966 53286
rect 11022 53284 11046 53286
rect 11102 53284 11126 53286
rect 11182 53284 11188 53286
rect 10880 53264 11188 53284
rect 13372 52698 13400 54742
rect 13360 52692 13412 52698
rect 13360 52634 13412 52640
rect 11796 52488 11848 52494
rect 11796 52430 11848 52436
rect 11888 52488 11940 52494
rect 11888 52430 11940 52436
rect 10880 52252 11188 52272
rect 10880 52250 10886 52252
rect 10942 52250 10966 52252
rect 11022 52250 11046 52252
rect 11102 52250 11126 52252
rect 11182 52250 11188 52252
rect 10942 52198 10944 52250
rect 11124 52198 11126 52250
rect 10880 52196 10886 52198
rect 10942 52196 10966 52198
rect 11022 52196 11046 52198
rect 11102 52196 11126 52198
rect 11182 52196 11188 52198
rect 10880 52176 11188 52196
rect 11808 52154 11836 52430
rect 11796 52148 11848 52154
rect 11796 52090 11848 52096
rect 11612 52012 11664 52018
rect 11612 51954 11664 51960
rect 10880 51164 11188 51184
rect 10880 51162 10886 51164
rect 10942 51162 10966 51164
rect 11022 51162 11046 51164
rect 11102 51162 11126 51164
rect 11182 51162 11188 51164
rect 10942 51110 10944 51162
rect 11124 51110 11126 51162
rect 10880 51108 10886 51110
rect 10942 51108 10966 51110
rect 11022 51108 11046 51110
rect 11102 51108 11126 51110
rect 11182 51108 11188 51110
rect 10880 51088 11188 51108
rect 10508 50244 10560 50250
rect 10508 50186 10560 50192
rect 9956 49224 10008 49230
rect 9956 49166 10008 49172
rect 9588 49156 9640 49162
rect 9588 49098 9640 49104
rect 9600 43450 9628 49098
rect 9864 49088 9916 49094
rect 9864 49030 9916 49036
rect 9772 44804 9824 44810
rect 9772 44746 9824 44752
rect 9680 43920 9732 43926
rect 9680 43862 9732 43868
rect 9588 43444 9640 43450
rect 9588 43386 9640 43392
rect 9692 42770 9720 43862
rect 9784 43722 9812 44746
rect 9772 43716 9824 43722
rect 9772 43658 9824 43664
rect 9876 43450 9904 49030
rect 9968 48890 9996 49166
rect 9956 48884 10008 48890
rect 9956 48826 10008 48832
rect 10048 45824 10100 45830
rect 10048 45766 10100 45772
rect 10060 44946 10088 45766
rect 10048 44940 10100 44946
rect 10048 44882 10100 44888
rect 10416 44736 10468 44742
rect 10416 44678 10468 44684
rect 10428 43858 10456 44678
rect 10416 43852 10468 43858
rect 10416 43794 10468 43800
rect 10140 43781 10192 43787
rect 10140 43723 10192 43729
rect 10324 43784 10376 43790
rect 10324 43726 10376 43732
rect 9956 43648 10008 43654
rect 9956 43590 10008 43596
rect 9968 43450 9996 43590
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9956 43444 10008 43450
rect 9956 43386 10008 43392
rect 9680 42764 9732 42770
rect 9680 42706 9732 42712
rect 9968 42090 9996 43386
rect 10048 43308 10100 43314
rect 10152 43296 10180 43723
rect 10100 43268 10180 43296
rect 10232 43308 10284 43314
rect 10048 43250 10100 43256
rect 10232 43250 10284 43256
rect 10060 42090 10088 43250
rect 10244 42226 10272 43250
rect 10336 43178 10364 43726
rect 10324 43172 10376 43178
rect 10324 43114 10376 43120
rect 10416 42696 10468 42702
rect 10416 42638 10468 42644
rect 10428 42362 10456 42638
rect 10416 42356 10468 42362
rect 10416 42298 10468 42304
rect 10232 42220 10284 42226
rect 10232 42162 10284 42168
rect 9956 42084 10008 42090
rect 9956 42026 10008 42032
rect 10048 42084 10100 42090
rect 10048 42026 10100 42032
rect 10324 42084 10376 42090
rect 10324 42026 10376 42032
rect 9864 40656 9916 40662
rect 9968 40644 9996 42026
rect 10060 41614 10088 42026
rect 10336 41818 10364 42026
rect 10324 41812 10376 41818
rect 10324 41754 10376 41760
rect 10048 41608 10100 41614
rect 10048 41550 10100 41556
rect 9916 40616 9996 40644
rect 9864 40598 9916 40604
rect 9680 40384 9732 40390
rect 9680 40326 9732 40332
rect 9588 37868 9640 37874
rect 9588 37810 9640 37816
rect 9600 37466 9628 37810
rect 9588 37460 9640 37466
rect 9588 37402 9640 37408
rect 9128 36790 9180 36796
rect 9494 36816 9550 36825
rect 8852 36780 8904 36786
rect 9600 36786 9628 37402
rect 9494 36751 9550 36760
rect 9588 36780 9640 36786
rect 8852 36722 8904 36728
rect 9588 36722 9640 36728
rect 8300 36168 8352 36174
rect 8300 36110 8352 36116
rect 8864 35766 8892 36722
rect 9692 36310 9720 40326
rect 9876 39914 9904 40598
rect 10060 40526 10088 41550
rect 10140 40724 10192 40730
rect 10140 40666 10192 40672
rect 10152 40594 10180 40666
rect 10140 40588 10192 40594
rect 10140 40530 10192 40536
rect 10324 40588 10376 40594
rect 10324 40530 10376 40536
rect 10048 40520 10100 40526
rect 10048 40462 10100 40468
rect 10060 39964 10088 40462
rect 10140 40384 10192 40390
rect 10140 40326 10192 40332
rect 10152 40118 10180 40326
rect 10336 40186 10364 40530
rect 10324 40180 10376 40186
rect 10324 40122 10376 40128
rect 10140 40112 10192 40118
rect 10140 40054 10192 40060
rect 10140 39976 10192 39982
rect 10060 39936 10140 39964
rect 10140 39918 10192 39924
rect 9864 39908 9916 39914
rect 9864 39850 9916 39856
rect 9956 39840 10008 39846
rect 9956 39782 10008 39788
rect 9968 38350 9996 39782
rect 10048 39296 10100 39302
rect 10048 39238 10100 39244
rect 9772 38344 9824 38350
rect 9772 38286 9824 38292
rect 9956 38344 10008 38350
rect 9956 38286 10008 38292
rect 9036 36304 9088 36310
rect 9036 36246 9088 36252
rect 9680 36304 9732 36310
rect 9680 36246 9732 36252
rect 9048 35766 9076 36246
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 8852 35760 8904 35766
rect 8852 35702 8904 35708
rect 9036 35760 9088 35766
rect 9036 35702 9088 35708
rect 9692 35290 9720 36110
rect 9680 35284 9732 35290
rect 9680 35226 9732 35232
rect 9784 34746 9812 38286
rect 9864 38208 9916 38214
rect 9864 38150 9916 38156
rect 9876 37942 9904 38150
rect 10060 38010 10088 39238
rect 10048 38004 10100 38010
rect 10048 37946 10100 37952
rect 9864 37936 9916 37942
rect 9864 37878 9916 37884
rect 10414 36680 10470 36689
rect 10414 36615 10470 36624
rect 10048 36100 10100 36106
rect 10048 36042 10100 36048
rect 9772 34740 9824 34746
rect 9772 34682 9824 34688
rect 9680 34604 9732 34610
rect 9680 34546 9732 34552
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 9692 34202 9720 34546
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9680 32836 9732 32842
rect 9680 32778 9732 32784
rect 9692 32434 9720 32778
rect 9784 32502 9812 33254
rect 9876 32910 9904 34546
rect 9956 33856 10008 33862
rect 9956 33798 10008 33804
rect 9864 32904 9916 32910
rect 9864 32846 9916 32852
rect 9772 32496 9824 32502
rect 9772 32438 9824 32444
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9692 31958 9720 32370
rect 9680 31952 9732 31958
rect 9680 31894 9732 31900
rect 9692 31346 9720 31894
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 9692 30734 9720 31282
rect 9680 30728 9732 30734
rect 9680 30670 9732 30676
rect 9784 26234 9812 31758
rect 9968 31754 9996 33798
rect 10060 31822 10088 36042
rect 10324 35080 10376 35086
rect 10324 35022 10376 35028
rect 10336 33386 10364 35022
rect 10324 33380 10376 33386
rect 10324 33322 10376 33328
rect 10428 32570 10456 36615
rect 10416 32564 10468 32570
rect 10416 32506 10468 32512
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 9876 31726 9996 31754
rect 10520 31754 10548 50186
rect 10880 50076 11188 50096
rect 10880 50074 10886 50076
rect 10942 50074 10966 50076
rect 11022 50074 11046 50076
rect 11102 50074 11126 50076
rect 11182 50074 11188 50076
rect 10942 50022 10944 50074
rect 11124 50022 11126 50074
rect 10880 50020 10886 50022
rect 10942 50020 10966 50022
rect 11022 50020 11046 50022
rect 11102 50020 11126 50022
rect 11182 50020 11188 50022
rect 10880 50000 11188 50020
rect 10968 49428 11020 49434
rect 10968 49370 11020 49376
rect 10980 49162 11008 49370
rect 10968 49156 11020 49162
rect 10968 49098 11020 49104
rect 11428 49088 11480 49094
rect 11428 49030 11480 49036
rect 10880 48988 11188 49008
rect 10880 48986 10886 48988
rect 10942 48986 10966 48988
rect 11022 48986 11046 48988
rect 11102 48986 11126 48988
rect 11182 48986 11188 48988
rect 10942 48934 10944 48986
rect 11124 48934 11126 48986
rect 10880 48932 10886 48934
rect 10942 48932 10966 48934
rect 11022 48932 11046 48934
rect 11102 48932 11126 48934
rect 11182 48932 11188 48934
rect 10880 48912 11188 48932
rect 11440 48754 11468 49030
rect 11428 48748 11480 48754
rect 11428 48690 11480 48696
rect 11624 48618 11652 51954
rect 11900 51074 11928 52430
rect 12624 51944 12676 51950
rect 12624 51886 12676 51892
rect 12900 51944 12952 51950
rect 12900 51886 12952 51892
rect 12636 51610 12664 51886
rect 12624 51604 12676 51610
rect 12624 51546 12676 51552
rect 12624 51264 12676 51270
rect 12624 51206 12676 51212
rect 11808 51046 11928 51074
rect 11704 49836 11756 49842
rect 11704 49778 11756 49784
rect 11612 48612 11664 48618
rect 11612 48554 11664 48560
rect 11716 48278 11744 49778
rect 11704 48272 11756 48278
rect 11704 48214 11756 48220
rect 10880 47900 11188 47920
rect 10880 47898 10886 47900
rect 10942 47898 10966 47900
rect 11022 47898 11046 47900
rect 11102 47898 11126 47900
rect 11182 47898 11188 47900
rect 10942 47846 10944 47898
rect 11124 47846 11126 47898
rect 10880 47844 10886 47846
rect 10942 47844 10966 47846
rect 11022 47844 11046 47846
rect 11102 47844 11126 47846
rect 11182 47844 11188 47846
rect 10880 47824 11188 47844
rect 10880 46812 11188 46832
rect 10880 46810 10886 46812
rect 10942 46810 10966 46812
rect 11022 46810 11046 46812
rect 11102 46810 11126 46812
rect 11182 46810 11188 46812
rect 10942 46758 10944 46810
rect 11124 46758 11126 46810
rect 10880 46756 10886 46758
rect 10942 46756 10966 46758
rect 11022 46756 11046 46758
rect 11102 46756 11126 46758
rect 11182 46756 11188 46758
rect 10880 46736 11188 46756
rect 11520 45892 11572 45898
rect 11520 45834 11572 45840
rect 10880 45724 11188 45744
rect 10880 45722 10886 45724
rect 10942 45722 10966 45724
rect 11022 45722 11046 45724
rect 11102 45722 11126 45724
rect 11182 45722 11188 45724
rect 10942 45670 10944 45722
rect 11124 45670 11126 45722
rect 10880 45668 10886 45670
rect 10942 45668 10966 45670
rect 11022 45668 11046 45670
rect 11102 45668 11126 45670
rect 11182 45668 11188 45670
rect 10880 45648 11188 45668
rect 10880 44636 11188 44656
rect 10880 44634 10886 44636
rect 10942 44634 10966 44636
rect 11022 44634 11046 44636
rect 11102 44634 11126 44636
rect 11182 44634 11188 44636
rect 10942 44582 10944 44634
rect 11124 44582 11126 44634
rect 10880 44580 10886 44582
rect 10942 44580 10966 44582
rect 11022 44580 11046 44582
rect 11102 44580 11126 44582
rect 11182 44580 11188 44582
rect 10880 44560 11188 44580
rect 11532 43722 11560 45834
rect 11704 45824 11756 45830
rect 11704 45766 11756 45772
rect 11716 44470 11744 45766
rect 11704 44464 11756 44470
rect 11704 44406 11756 44412
rect 11612 44396 11664 44402
rect 11612 44338 11664 44344
rect 11624 44305 11652 44338
rect 11808 44334 11836 51046
rect 11888 50312 11940 50318
rect 11888 50254 11940 50260
rect 11900 49978 11928 50254
rect 12256 50244 12308 50250
rect 12256 50186 12308 50192
rect 11888 49972 11940 49978
rect 11888 49914 11940 49920
rect 12072 49292 12124 49298
rect 12072 49234 12124 49240
rect 11980 48816 12032 48822
rect 11980 48758 12032 48764
rect 11888 46572 11940 46578
rect 11888 46514 11940 46520
rect 11796 44328 11848 44334
rect 11610 44296 11666 44305
rect 11796 44270 11848 44276
rect 11610 44231 11666 44240
rect 11520 43716 11572 43722
rect 11520 43658 11572 43664
rect 10880 43548 11188 43568
rect 10880 43546 10886 43548
rect 10942 43546 10966 43548
rect 11022 43546 11046 43548
rect 11102 43546 11126 43548
rect 11182 43546 11188 43548
rect 10942 43494 10944 43546
rect 11124 43494 11126 43546
rect 10880 43492 10886 43494
rect 10942 43492 10966 43494
rect 11022 43492 11046 43494
rect 11102 43492 11126 43494
rect 11182 43492 11188 43494
rect 10880 43472 11188 43492
rect 11532 42770 11560 43658
rect 11520 42764 11572 42770
rect 11520 42706 11572 42712
rect 10880 42460 11188 42480
rect 10880 42458 10886 42460
rect 10942 42458 10966 42460
rect 11022 42458 11046 42460
rect 11102 42458 11126 42460
rect 11182 42458 11188 42460
rect 10942 42406 10944 42458
rect 11124 42406 11126 42458
rect 10880 42404 10886 42406
rect 10942 42404 10966 42406
rect 11022 42404 11046 42406
rect 11102 42404 11126 42406
rect 11182 42404 11188 42406
rect 10880 42384 11188 42404
rect 11900 42362 11928 46514
rect 11992 45830 12020 48758
rect 12084 48686 12112 49234
rect 12164 49088 12216 49094
rect 12164 49030 12216 49036
rect 12176 48822 12204 49030
rect 12164 48816 12216 48822
rect 12164 48758 12216 48764
rect 12072 48680 12124 48686
rect 12072 48622 12124 48628
rect 12164 48680 12216 48686
rect 12164 48622 12216 48628
rect 12084 48142 12112 48622
rect 12072 48136 12124 48142
rect 12072 48078 12124 48084
rect 12176 48006 12204 48622
rect 12164 48000 12216 48006
rect 12164 47942 12216 47948
rect 12176 45898 12204 47942
rect 12164 45892 12216 45898
rect 12164 45834 12216 45840
rect 11980 45824 12032 45830
rect 11980 45766 12032 45772
rect 12268 45082 12296 50186
rect 12532 49768 12584 49774
rect 12532 49710 12584 49716
rect 12348 49156 12400 49162
rect 12348 49098 12400 49104
rect 12360 48686 12388 49098
rect 12348 48680 12400 48686
rect 12348 48622 12400 48628
rect 12440 46028 12492 46034
rect 12440 45970 12492 45976
rect 12256 45076 12308 45082
rect 12256 45018 12308 45024
rect 12452 44538 12480 45970
rect 12544 45558 12572 49710
rect 12636 49230 12664 51206
rect 12624 49224 12676 49230
rect 12624 49166 12676 49172
rect 12808 46640 12860 46646
rect 12808 46582 12860 46588
rect 12624 46096 12676 46102
rect 12624 46038 12676 46044
rect 12532 45552 12584 45558
rect 12532 45494 12584 45500
rect 12532 45416 12584 45422
rect 12532 45358 12584 45364
rect 12544 45098 12572 45358
rect 12636 45286 12664 46038
rect 12716 45892 12768 45898
rect 12716 45834 12768 45840
rect 12624 45280 12676 45286
rect 12624 45222 12676 45228
rect 12728 45098 12756 45834
rect 12820 45558 12848 46582
rect 12912 46170 12940 51886
rect 13084 50176 13136 50182
rect 13084 50118 13136 50124
rect 12900 46164 12952 46170
rect 12900 46106 12952 46112
rect 12900 45824 12952 45830
rect 12900 45766 12952 45772
rect 12808 45552 12860 45558
rect 12808 45494 12860 45500
rect 12544 45070 12756 45098
rect 12544 44810 12572 45070
rect 12532 44804 12584 44810
rect 12532 44746 12584 44752
rect 12348 44532 12400 44538
rect 12348 44474 12400 44480
rect 12440 44532 12492 44538
rect 12440 44474 12492 44480
rect 12360 44441 12388 44474
rect 12346 44432 12402 44441
rect 12072 44396 12124 44402
rect 12346 44367 12402 44376
rect 12072 44338 12124 44344
rect 12084 44266 12112 44338
rect 12072 44260 12124 44266
rect 12072 44202 12124 44208
rect 12452 44010 12480 44474
rect 12532 44396 12584 44402
rect 12532 44338 12584 44344
rect 12360 43982 12480 44010
rect 12544 43994 12572 44338
rect 12728 44334 12756 45070
rect 12912 44946 12940 45766
rect 13096 45014 13124 50118
rect 13176 49156 13228 49162
rect 13176 49098 13228 49104
rect 13188 46714 13216 49098
rect 13360 48068 13412 48074
rect 13360 48010 13412 48016
rect 13176 46708 13228 46714
rect 13176 46650 13228 46656
rect 13084 45008 13136 45014
rect 13084 44950 13136 44956
rect 12900 44940 12952 44946
rect 12820 44900 12900 44928
rect 12820 44470 12848 44900
rect 12900 44882 12952 44888
rect 12992 44872 13044 44878
rect 12992 44814 13044 44820
rect 12808 44464 12860 44470
rect 12808 44406 12860 44412
rect 12898 44432 12954 44441
rect 12716 44328 12768 44334
rect 12716 44270 12768 44276
rect 12532 43988 12584 43994
rect 12360 43858 12388 43982
rect 12532 43930 12584 43936
rect 12728 43926 12756 44270
rect 12716 43920 12768 43926
rect 12716 43862 12768 43868
rect 12348 43852 12400 43858
rect 12348 43794 12400 43800
rect 12820 43790 12848 44406
rect 12898 44367 12954 44376
rect 12808 43784 12860 43790
rect 12808 43726 12860 43732
rect 12164 43648 12216 43654
rect 12164 43590 12216 43596
rect 12072 43240 12124 43246
rect 12072 43182 12124 43188
rect 11980 42628 12032 42634
rect 11980 42570 12032 42576
rect 11888 42356 11940 42362
rect 11888 42298 11940 42304
rect 11992 42022 12020 42570
rect 12084 42090 12112 43182
rect 12072 42084 12124 42090
rect 12072 42026 12124 42032
rect 11980 42016 12032 42022
rect 11980 41958 12032 41964
rect 10880 41372 11188 41392
rect 10880 41370 10886 41372
rect 10942 41370 10966 41372
rect 11022 41370 11046 41372
rect 11102 41370 11126 41372
rect 11182 41370 11188 41372
rect 10942 41318 10944 41370
rect 11124 41318 11126 41370
rect 10880 41316 10886 41318
rect 10942 41316 10966 41318
rect 11022 41316 11046 41318
rect 11102 41316 11126 41318
rect 11182 41316 11188 41318
rect 10880 41296 11188 41316
rect 11244 40588 11296 40594
rect 11244 40530 11296 40536
rect 10880 40284 11188 40304
rect 10880 40282 10886 40284
rect 10942 40282 10966 40284
rect 11022 40282 11046 40284
rect 11102 40282 11126 40284
rect 11182 40282 11188 40284
rect 10942 40230 10944 40282
rect 11124 40230 11126 40282
rect 10880 40228 10886 40230
rect 10942 40228 10966 40230
rect 11022 40228 11046 40230
rect 11102 40228 11126 40230
rect 11182 40228 11188 40230
rect 10880 40208 11188 40228
rect 10600 39908 10652 39914
rect 10600 39850 10652 39856
rect 10612 39506 10640 39850
rect 10600 39500 10652 39506
rect 10600 39442 10652 39448
rect 10880 39196 11188 39216
rect 10880 39194 10886 39196
rect 10942 39194 10966 39196
rect 11022 39194 11046 39196
rect 11102 39194 11126 39196
rect 11182 39194 11188 39196
rect 10942 39142 10944 39194
rect 11124 39142 11126 39194
rect 10880 39140 10886 39142
rect 10942 39140 10966 39142
rect 11022 39140 11046 39142
rect 11102 39140 11126 39142
rect 11182 39140 11188 39142
rect 10880 39120 11188 39140
rect 11256 38554 11284 40530
rect 11336 40452 11388 40458
rect 11336 40394 11388 40400
rect 11244 38548 11296 38554
rect 11244 38490 11296 38496
rect 10880 38108 11188 38128
rect 10880 38106 10886 38108
rect 10942 38106 10966 38108
rect 11022 38106 11046 38108
rect 11102 38106 11126 38108
rect 11182 38106 11188 38108
rect 10942 38054 10944 38106
rect 11124 38054 11126 38106
rect 10880 38052 10886 38054
rect 10942 38052 10966 38054
rect 11022 38052 11046 38054
rect 11102 38052 11126 38054
rect 11182 38052 11188 38054
rect 10880 38032 11188 38052
rect 10880 37020 11188 37040
rect 10880 37018 10886 37020
rect 10942 37018 10966 37020
rect 11022 37018 11046 37020
rect 11102 37018 11126 37020
rect 11182 37018 11188 37020
rect 10942 36966 10944 37018
rect 11124 36966 11126 37018
rect 10880 36964 10886 36966
rect 10942 36964 10966 36966
rect 11022 36964 11046 36966
rect 11102 36964 11126 36966
rect 11182 36964 11188 36966
rect 10880 36944 11188 36964
rect 11348 36378 11376 40394
rect 11520 39840 11572 39846
rect 11520 39782 11572 39788
rect 11428 39432 11480 39438
rect 11428 39374 11480 39380
rect 11440 38418 11468 39374
rect 11428 38412 11480 38418
rect 11428 38354 11480 38360
rect 11428 37868 11480 37874
rect 11428 37810 11480 37816
rect 11336 36372 11388 36378
rect 11336 36314 11388 36320
rect 10880 35932 11188 35952
rect 10880 35930 10886 35932
rect 10942 35930 10966 35932
rect 11022 35930 11046 35932
rect 11102 35930 11126 35932
rect 11182 35930 11188 35932
rect 10942 35878 10944 35930
rect 11124 35878 11126 35930
rect 10880 35876 10886 35878
rect 10942 35876 10966 35878
rect 11022 35876 11046 35878
rect 11102 35876 11126 35878
rect 11182 35876 11188 35878
rect 10880 35856 11188 35876
rect 10600 35012 10652 35018
rect 10600 34954 10652 34960
rect 10612 33114 10640 34954
rect 10880 34844 11188 34864
rect 10880 34842 10886 34844
rect 10942 34842 10966 34844
rect 11022 34842 11046 34844
rect 11102 34842 11126 34844
rect 11182 34842 11188 34844
rect 10942 34790 10944 34842
rect 11124 34790 11126 34842
rect 10880 34788 10886 34790
rect 10942 34788 10966 34790
rect 11022 34788 11046 34790
rect 11102 34788 11126 34790
rect 11182 34788 11188 34790
rect 10880 34768 11188 34788
rect 10784 34468 10836 34474
rect 10784 34410 10836 34416
rect 10796 33998 10824 34410
rect 11244 34060 11296 34066
rect 11244 34002 11296 34008
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10796 33454 10824 33934
rect 10880 33756 11188 33776
rect 10880 33754 10886 33756
rect 10942 33754 10966 33756
rect 11022 33754 11046 33756
rect 11102 33754 11126 33756
rect 11182 33754 11188 33756
rect 10942 33702 10944 33754
rect 11124 33702 11126 33754
rect 10880 33700 10886 33702
rect 10942 33700 10966 33702
rect 11022 33700 11046 33702
rect 11102 33700 11126 33702
rect 11182 33700 11188 33702
rect 10880 33680 11188 33700
rect 11256 33522 11284 34002
rect 11244 33516 11296 33522
rect 11244 33458 11296 33464
rect 10784 33448 10836 33454
rect 10784 33390 10836 33396
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 11256 33046 11284 33458
rect 11336 33108 11388 33114
rect 11336 33050 11388 33056
rect 11244 33040 11296 33046
rect 11244 32982 11296 32988
rect 10880 32668 11188 32688
rect 10880 32666 10886 32668
rect 10942 32666 10966 32668
rect 11022 32666 11046 32668
rect 11102 32666 11126 32668
rect 11182 32666 11188 32668
rect 10942 32614 10944 32666
rect 11124 32614 11126 32666
rect 10880 32612 10886 32614
rect 10942 32612 10966 32614
rect 11022 32612 11046 32614
rect 11102 32612 11126 32614
rect 11182 32612 11188 32614
rect 10880 32592 11188 32612
rect 11152 32496 11204 32502
rect 11152 32438 11204 32444
rect 11060 32292 11112 32298
rect 11060 32234 11112 32240
rect 11072 31822 11100 32234
rect 11060 31816 11112 31822
rect 11060 31758 11112 31764
rect 11164 31754 11192 32438
rect 11256 32298 11284 32982
rect 11244 32292 11296 32298
rect 11244 32234 11296 32240
rect 11244 31952 11296 31958
rect 11244 31894 11296 31900
rect 10520 31726 10640 31754
rect 9876 30734 9904 31726
rect 9956 31204 10008 31210
rect 9956 31146 10008 31152
rect 9968 30802 9996 31146
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 10612 28966 10640 31726
rect 11152 31748 11204 31754
rect 11152 31690 11204 31696
rect 10880 31580 11188 31600
rect 10880 31578 10886 31580
rect 10942 31578 10966 31580
rect 11022 31578 11046 31580
rect 11102 31578 11126 31580
rect 11182 31578 11188 31580
rect 10942 31526 10944 31578
rect 11124 31526 11126 31578
rect 10880 31524 10886 31526
rect 10942 31524 10966 31526
rect 11022 31524 11046 31526
rect 11102 31524 11126 31526
rect 11182 31524 11188 31526
rect 10880 31504 11188 31524
rect 11256 30734 11284 31894
rect 11348 31890 11376 33050
rect 11440 32026 11468 37810
rect 11532 33862 11560 39782
rect 11888 39636 11940 39642
rect 11888 39578 11940 39584
rect 11612 39432 11664 39438
rect 11612 39374 11664 39380
rect 11624 38010 11652 39374
rect 11704 39364 11756 39370
rect 11704 39306 11756 39312
rect 11716 39098 11744 39306
rect 11900 39098 11928 39578
rect 11704 39092 11756 39098
rect 11704 39034 11756 39040
rect 11888 39092 11940 39098
rect 11888 39034 11940 39040
rect 11796 38752 11848 38758
rect 11796 38694 11848 38700
rect 11612 38004 11664 38010
rect 11612 37946 11664 37952
rect 11612 37800 11664 37806
rect 11612 37742 11664 37748
rect 11624 35290 11652 37742
rect 11808 37398 11836 38694
rect 11796 37392 11848 37398
rect 11796 37334 11848 37340
rect 11704 37120 11756 37126
rect 11704 37062 11756 37068
rect 11612 35284 11664 35290
rect 11612 35226 11664 35232
rect 11520 33856 11572 33862
rect 11520 33798 11572 33804
rect 11612 33856 11664 33862
rect 11612 33798 11664 33804
rect 11520 33584 11572 33590
rect 11520 33526 11572 33532
rect 11532 32774 11560 33526
rect 11624 33522 11652 33798
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11612 33380 11664 33386
rect 11612 33322 11664 33328
rect 11624 32910 11652 33322
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11532 32502 11560 32710
rect 11520 32496 11572 32502
rect 11520 32438 11572 32444
rect 11428 32020 11480 32026
rect 11428 31962 11480 31968
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 11716 31754 11744 37062
rect 11992 36106 12020 41958
rect 12084 41682 12112 42026
rect 12072 41676 12124 41682
rect 12072 41618 12124 41624
rect 12176 39846 12204 43590
rect 12820 43382 12848 43726
rect 12808 43376 12860 43382
rect 12808 43318 12860 43324
rect 12808 43240 12860 43246
rect 12808 43182 12860 43188
rect 12820 42906 12848 43182
rect 12808 42900 12860 42906
rect 12808 42842 12860 42848
rect 12912 41818 12940 44367
rect 13004 44198 13032 44814
rect 13188 44470 13216 46650
rect 13268 46096 13320 46102
rect 13268 46038 13320 46044
rect 13280 45966 13308 46038
rect 13268 45960 13320 45966
rect 13268 45902 13320 45908
rect 13268 45824 13320 45830
rect 13268 45766 13320 45772
rect 13280 45558 13308 45766
rect 13268 45552 13320 45558
rect 13268 45494 13320 45500
rect 13372 45354 13400 48010
rect 13360 45348 13412 45354
rect 13360 45290 13412 45296
rect 13372 44878 13400 45290
rect 13360 44872 13412 44878
rect 13360 44814 13412 44820
rect 13268 44736 13320 44742
rect 13268 44678 13320 44684
rect 13176 44464 13228 44470
rect 13176 44406 13228 44412
rect 12992 44192 13044 44198
rect 12992 44134 13044 44140
rect 12992 43920 13044 43926
rect 12992 43862 13044 43868
rect 13004 42566 13032 43862
rect 13084 43784 13136 43790
rect 13082 43752 13084 43761
rect 13136 43752 13138 43761
rect 13082 43687 13138 43696
rect 13084 43648 13136 43654
rect 13084 43590 13136 43596
rect 13096 43314 13124 43590
rect 13084 43308 13136 43314
rect 13084 43250 13136 43256
rect 13280 43246 13308 44678
rect 13268 43240 13320 43246
rect 13268 43182 13320 43188
rect 12992 42560 13044 42566
rect 12992 42502 13044 42508
rect 12900 41812 12952 41818
rect 12900 41754 12952 41760
rect 12348 41540 12400 41546
rect 12348 41482 12400 41488
rect 12164 39840 12216 39846
rect 12164 39782 12216 39788
rect 12164 39296 12216 39302
rect 12164 39238 12216 39244
rect 12176 38962 12204 39238
rect 12164 38956 12216 38962
rect 12164 38898 12216 38904
rect 12164 38820 12216 38826
rect 12164 38762 12216 38768
rect 12070 38720 12126 38729
rect 12070 38655 12126 38664
rect 11980 36100 12032 36106
rect 11980 36042 12032 36048
rect 11796 34400 11848 34406
rect 11796 34342 11848 34348
rect 11888 34400 11940 34406
rect 11888 34342 11940 34348
rect 11808 32502 11836 34342
rect 11900 34066 11928 34342
rect 11888 34060 11940 34066
rect 11888 34002 11940 34008
rect 12084 33658 12112 38655
rect 12176 38350 12204 38762
rect 12164 38344 12216 38350
rect 12164 38286 12216 38292
rect 12176 37942 12204 38286
rect 12164 37936 12216 37942
rect 12164 37878 12216 37884
rect 12176 37466 12204 37878
rect 12256 37664 12308 37670
rect 12256 37606 12308 37612
rect 12164 37460 12216 37466
rect 12164 37402 12216 37408
rect 12268 37194 12296 37606
rect 12256 37188 12308 37194
rect 12256 37130 12308 37136
rect 12360 35290 12388 41482
rect 12912 40118 12940 41754
rect 12900 40112 12952 40118
rect 12900 40054 12952 40060
rect 12716 39296 12768 39302
rect 12716 39238 12768 39244
rect 12532 39024 12584 39030
rect 12532 38966 12584 38972
rect 12440 37868 12492 37874
rect 12440 37810 12492 37816
rect 12452 37466 12480 37810
rect 12440 37460 12492 37466
rect 12440 37402 12492 37408
rect 12544 37398 12572 38966
rect 12728 38706 12756 39238
rect 13464 39114 13492 59570
rect 13556 59022 13584 59706
rect 13544 59016 13596 59022
rect 13544 58958 13596 58964
rect 13544 58336 13596 58342
rect 13544 58278 13596 58284
rect 13556 58070 13584 58278
rect 13544 58064 13596 58070
rect 13544 58006 13596 58012
rect 13832 57934 13860 63310
rect 13924 60734 13952 63718
rect 14200 63374 14228 66642
rect 14568 66638 14596 67050
rect 14740 67040 14792 67046
rect 14740 66982 14792 66988
rect 14752 66638 14780 66982
rect 14936 66842 14964 67186
rect 15212 67114 15240 67526
rect 15200 67108 15252 67114
rect 15200 67050 15252 67056
rect 15384 67040 15436 67046
rect 15384 66982 15436 66988
rect 14924 66836 14976 66842
rect 14924 66778 14976 66784
rect 15396 66638 15424 66982
rect 14556 66632 14608 66638
rect 14556 66574 14608 66580
rect 14740 66632 14792 66638
rect 14740 66574 14792 66580
rect 15292 66632 15344 66638
rect 15292 66574 15344 66580
rect 15384 66632 15436 66638
rect 15384 66574 15436 66580
rect 14832 66564 14884 66570
rect 14832 66506 14884 66512
rect 14844 65958 14872 66506
rect 14832 65952 14884 65958
rect 14832 65894 14884 65900
rect 14556 65000 14608 65006
rect 14556 64942 14608 64948
rect 14568 63918 14596 64942
rect 14648 64048 14700 64054
rect 14648 63990 14700 63996
rect 14556 63912 14608 63918
rect 14556 63854 14608 63860
rect 14188 63368 14240 63374
rect 14188 63310 14240 63316
rect 14568 63306 14596 63854
rect 14556 63300 14608 63306
rect 14556 63242 14608 63248
rect 14096 61940 14148 61946
rect 14096 61882 14148 61888
rect 13924 60722 14044 60734
rect 13924 60716 14056 60722
rect 13924 60706 14004 60716
rect 14004 60658 14056 60664
rect 14004 60580 14056 60586
rect 14108 60568 14136 61882
rect 14280 60648 14332 60654
rect 14280 60590 14332 60596
rect 14056 60540 14136 60568
rect 14004 60522 14056 60528
rect 13820 57928 13872 57934
rect 13820 57870 13872 57876
rect 13636 57452 13688 57458
rect 13636 57394 13688 57400
rect 13648 57050 13676 57394
rect 13832 57322 13860 57870
rect 14016 57440 14044 60522
rect 14096 60240 14148 60246
rect 14096 60182 14148 60188
rect 14108 59634 14136 60182
rect 14292 59770 14320 60590
rect 14464 60036 14516 60042
rect 14464 59978 14516 59984
rect 14280 59764 14332 59770
rect 14280 59706 14332 59712
rect 14096 59628 14148 59634
rect 14096 59570 14148 59576
rect 14476 58886 14504 59978
rect 14568 59922 14596 63242
rect 14660 63238 14688 63990
rect 14648 63232 14700 63238
rect 14648 63174 14700 63180
rect 14660 62150 14688 63174
rect 14648 62144 14700 62150
rect 14648 62086 14700 62092
rect 14660 60042 14688 62086
rect 14740 61600 14792 61606
rect 14740 61542 14792 61548
rect 14752 60518 14780 61542
rect 14740 60512 14792 60518
rect 14740 60454 14792 60460
rect 14648 60036 14700 60042
rect 14648 59978 14700 59984
rect 14740 60036 14792 60042
rect 14740 59978 14792 59984
rect 14752 59922 14780 59978
rect 14568 59894 14780 59922
rect 14464 58880 14516 58886
rect 14464 58822 14516 58828
rect 14188 57792 14240 57798
rect 14188 57734 14240 57740
rect 14200 57458 14228 57734
rect 14096 57452 14148 57458
rect 14016 57412 14096 57440
rect 14096 57394 14148 57400
rect 14188 57452 14240 57458
rect 14188 57394 14240 57400
rect 13820 57316 13872 57322
rect 13820 57258 13872 57264
rect 13636 57044 13688 57050
rect 13636 56986 13688 56992
rect 14004 56840 14056 56846
rect 14004 56782 14056 56788
rect 14016 56234 14044 56782
rect 14004 56228 14056 56234
rect 14004 56170 14056 56176
rect 14108 56166 14136 57394
rect 14188 57248 14240 57254
rect 14188 57190 14240 57196
rect 14200 56846 14228 57190
rect 14188 56840 14240 56846
rect 14188 56782 14240 56788
rect 14476 56302 14504 58822
rect 14752 56370 14780 59894
rect 14844 59430 14872 65894
rect 15304 65754 15332 66574
rect 15292 65748 15344 65754
rect 15292 65690 15344 65696
rect 15292 65544 15344 65550
rect 15292 65486 15344 65492
rect 15304 65210 15332 65486
rect 15292 65204 15344 65210
rect 15292 65146 15344 65152
rect 15488 64870 15516 70518
rect 15580 70514 15608 70790
rect 15568 70508 15620 70514
rect 15568 70450 15620 70456
rect 15752 70304 15804 70310
rect 15752 70246 15804 70252
rect 15764 69902 15792 70246
rect 15846 70204 16154 70224
rect 15846 70202 15852 70204
rect 15908 70202 15932 70204
rect 15988 70202 16012 70204
rect 16068 70202 16092 70204
rect 16148 70202 16154 70204
rect 15908 70150 15910 70202
rect 16090 70150 16092 70202
rect 15846 70148 15852 70150
rect 15908 70148 15932 70150
rect 15988 70148 16012 70150
rect 16068 70148 16092 70150
rect 16148 70148 16154 70150
rect 15846 70128 16154 70148
rect 15752 69896 15804 69902
rect 15752 69838 15804 69844
rect 16212 69760 16264 69766
rect 16212 69702 16264 69708
rect 15846 69116 16154 69136
rect 15846 69114 15852 69116
rect 15908 69114 15932 69116
rect 15988 69114 16012 69116
rect 16068 69114 16092 69116
rect 16148 69114 16154 69116
rect 15908 69062 15910 69114
rect 16090 69062 16092 69114
rect 15846 69060 15852 69062
rect 15908 69060 15932 69062
rect 15988 69060 16012 69062
rect 16068 69060 16092 69062
rect 16148 69060 16154 69062
rect 15846 69040 16154 69060
rect 16224 68950 16252 69702
rect 16304 69216 16356 69222
rect 16304 69158 16356 69164
rect 16212 68944 16264 68950
rect 16212 68886 16264 68892
rect 16316 68474 16344 69158
rect 16304 68468 16356 68474
rect 16304 68410 16356 68416
rect 15846 68028 16154 68048
rect 15846 68026 15852 68028
rect 15908 68026 15932 68028
rect 15988 68026 16012 68028
rect 16068 68026 16092 68028
rect 16148 68026 16154 68028
rect 15908 67974 15910 68026
rect 16090 67974 16092 68026
rect 15846 67972 15852 67974
rect 15908 67972 15932 67974
rect 15988 67972 16012 67974
rect 16068 67972 16092 67974
rect 16148 67972 16154 67974
rect 15846 67952 16154 67972
rect 15846 66940 16154 66960
rect 15846 66938 15852 66940
rect 15908 66938 15932 66940
rect 15988 66938 16012 66940
rect 16068 66938 16092 66940
rect 16148 66938 16154 66940
rect 15908 66886 15910 66938
rect 16090 66886 16092 66938
rect 15846 66884 15852 66886
rect 15908 66884 15932 66886
rect 15988 66884 16012 66886
rect 16068 66884 16092 66886
rect 16148 66884 16154 66886
rect 15846 66864 16154 66884
rect 16316 66586 16344 68410
rect 16408 66706 16436 71130
rect 16500 71058 16528 72694
rect 16488 71052 16540 71058
rect 16488 70994 16540 71000
rect 16592 70990 16620 74122
rect 16684 73914 16712 75210
rect 16776 74730 16804 75890
rect 17040 75744 17092 75750
rect 17040 75686 17092 75692
rect 17052 75410 17080 75686
rect 17040 75404 17092 75410
rect 17040 75346 17092 75352
rect 16856 75268 16908 75274
rect 16856 75210 16908 75216
rect 16764 74724 16816 74730
rect 16764 74666 16816 74672
rect 16672 73908 16724 73914
rect 16672 73850 16724 73856
rect 16868 73098 16896 75210
rect 16948 75200 17000 75206
rect 16948 75142 17000 75148
rect 17040 75200 17092 75206
rect 17040 75142 17092 75148
rect 16960 73778 16988 75142
rect 16948 73772 17000 73778
rect 16948 73714 17000 73720
rect 16960 73302 16988 73714
rect 16948 73296 17000 73302
rect 16948 73238 17000 73244
rect 16856 73092 16908 73098
rect 16856 73034 16908 73040
rect 17052 73030 17080 75142
rect 17224 74928 17276 74934
rect 17224 74870 17276 74876
rect 17236 74118 17264 74870
rect 17960 74860 18012 74866
rect 17960 74802 18012 74808
rect 17224 74112 17276 74118
rect 17224 74054 17276 74060
rect 17040 73024 17092 73030
rect 17040 72966 17092 72972
rect 16948 71936 17000 71942
rect 16948 71878 17000 71884
rect 16580 70984 16632 70990
rect 16580 70926 16632 70932
rect 16960 70514 16988 71878
rect 16948 70508 17000 70514
rect 16948 70450 17000 70456
rect 16764 70440 16816 70446
rect 16764 70382 16816 70388
rect 16672 69352 16724 69358
rect 16672 69294 16724 69300
rect 16684 67726 16712 69294
rect 16776 69018 16804 70382
rect 16764 69012 16816 69018
rect 16764 68954 16816 68960
rect 16672 67720 16724 67726
rect 16672 67662 16724 67668
rect 17052 67182 17080 72966
rect 17132 72684 17184 72690
rect 17132 72626 17184 72632
rect 17144 69766 17172 72626
rect 17236 72486 17264 74054
rect 17972 73914 18000 74802
rect 18236 74792 18288 74798
rect 18236 74734 18288 74740
rect 18248 74458 18276 74734
rect 18236 74452 18288 74458
rect 18236 74394 18288 74400
rect 19076 74390 19104 75890
rect 19892 75812 19944 75818
rect 19892 75754 19944 75760
rect 19616 75744 19668 75750
rect 19616 75686 19668 75692
rect 19708 75744 19760 75750
rect 19708 75686 19760 75692
rect 19628 75410 19656 75686
rect 19616 75404 19668 75410
rect 19616 75346 19668 75352
rect 19720 75342 19748 75686
rect 19708 75336 19760 75342
rect 19708 75278 19760 75284
rect 19904 75274 19932 75754
rect 19892 75268 19944 75274
rect 19892 75210 19944 75216
rect 20180 74934 20208 75890
rect 21192 75546 21220 76230
rect 21548 75880 21600 75886
rect 21548 75822 21600 75828
rect 21180 75540 21232 75546
rect 21180 75482 21232 75488
rect 21192 75206 21220 75482
rect 21272 75268 21324 75274
rect 21272 75210 21324 75216
rect 21180 75200 21232 75206
rect 21180 75142 21232 75148
rect 20811 75100 21119 75120
rect 20811 75098 20817 75100
rect 20873 75098 20897 75100
rect 20953 75098 20977 75100
rect 21033 75098 21057 75100
rect 21113 75098 21119 75100
rect 20873 75046 20875 75098
rect 21055 75046 21057 75098
rect 20811 75044 20817 75046
rect 20873 75044 20897 75046
rect 20953 75044 20977 75046
rect 21033 75044 21057 75046
rect 21113 75044 21119 75046
rect 20811 75024 21119 75044
rect 20168 74928 20220 74934
rect 20168 74870 20220 74876
rect 20720 74928 20772 74934
rect 20720 74870 20772 74876
rect 20076 74656 20128 74662
rect 20076 74598 20128 74604
rect 19892 74452 19944 74458
rect 19892 74394 19944 74400
rect 19064 74384 19116 74390
rect 19064 74326 19116 74332
rect 18420 74316 18472 74322
rect 18420 74258 18472 74264
rect 17960 73908 18012 73914
rect 17960 73850 18012 73856
rect 17868 73840 17920 73846
rect 17868 73782 17920 73788
rect 17500 73772 17552 73778
rect 17500 73714 17552 73720
rect 17316 73636 17368 73642
rect 17316 73578 17368 73584
rect 17328 73234 17356 73578
rect 17512 73370 17540 73714
rect 17500 73364 17552 73370
rect 17500 73306 17552 73312
rect 17316 73228 17368 73234
rect 17316 73170 17368 73176
rect 17224 72480 17276 72486
rect 17224 72422 17276 72428
rect 17236 70854 17264 72422
rect 17328 72078 17356 73170
rect 17408 73160 17460 73166
rect 17406 73128 17408 73137
rect 17460 73128 17462 73137
rect 17406 73063 17462 73072
rect 17880 73030 17908 73782
rect 18236 73772 18288 73778
rect 18236 73714 18288 73720
rect 18248 73574 18276 73714
rect 18432 73642 18460 74258
rect 19904 74186 19932 74394
rect 19524 74180 19576 74186
rect 19524 74122 19576 74128
rect 19892 74180 19944 74186
rect 19892 74122 19944 74128
rect 19536 73846 19564 74122
rect 19708 74112 19760 74118
rect 19708 74054 19760 74060
rect 19720 73914 19748 74054
rect 19708 73908 19760 73914
rect 19708 73850 19760 73856
rect 19524 73840 19576 73846
rect 19524 73782 19576 73788
rect 18420 73636 18472 73642
rect 18420 73578 18472 73584
rect 18236 73568 18288 73574
rect 18236 73510 18288 73516
rect 19536 73370 19564 73782
rect 19720 73370 19748 73850
rect 19904 73710 19932 74122
rect 19892 73704 19944 73710
rect 19892 73646 19944 73652
rect 19524 73364 19576 73370
rect 19524 73306 19576 73312
rect 19708 73364 19760 73370
rect 19708 73306 19760 73312
rect 19708 73092 19760 73098
rect 19708 73034 19760 73040
rect 17868 73024 17920 73030
rect 17868 72966 17920 72972
rect 17880 72146 17908 72966
rect 18236 72616 18288 72622
rect 18236 72558 18288 72564
rect 17960 72548 18012 72554
rect 17960 72490 18012 72496
rect 17868 72140 17920 72146
rect 17868 72082 17920 72088
rect 17316 72072 17368 72078
rect 17316 72014 17368 72020
rect 17328 71738 17356 72014
rect 17316 71732 17368 71738
rect 17316 71674 17368 71680
rect 17224 70848 17276 70854
rect 17224 70790 17276 70796
rect 17132 69760 17184 69766
rect 17132 69702 17184 69708
rect 17328 69426 17356 71674
rect 17500 71596 17552 71602
rect 17500 71538 17552 71544
rect 17512 71505 17540 71538
rect 17880 71534 17908 72082
rect 17972 71602 18000 72490
rect 18144 72276 18196 72282
rect 18144 72218 18196 72224
rect 17960 71596 18012 71602
rect 17960 71538 18012 71544
rect 17868 71528 17920 71534
rect 17498 71496 17554 71505
rect 17868 71470 17920 71476
rect 17498 71431 17554 71440
rect 17408 70984 17460 70990
rect 17408 70926 17460 70932
rect 17420 69850 17448 70926
rect 17420 69822 17540 69850
rect 17408 69760 17460 69766
rect 17408 69702 17460 69708
rect 17316 69420 17368 69426
rect 17316 69362 17368 69368
rect 17316 68740 17368 68746
rect 17316 68682 17368 68688
rect 17328 68134 17356 68682
rect 17316 68128 17368 68134
rect 17316 68070 17368 68076
rect 17040 67176 17092 67182
rect 17040 67118 17092 67124
rect 16396 66700 16448 66706
rect 16396 66642 16448 66648
rect 16316 66558 16436 66586
rect 15846 65852 16154 65872
rect 15846 65850 15852 65852
rect 15908 65850 15932 65852
rect 15988 65850 16012 65852
rect 16068 65850 16092 65852
rect 16148 65850 16154 65852
rect 15908 65798 15910 65850
rect 16090 65798 16092 65850
rect 15846 65796 15852 65798
rect 15908 65796 15932 65798
rect 15988 65796 16012 65798
rect 16068 65796 16092 65798
rect 16148 65796 16154 65798
rect 15846 65776 16154 65796
rect 15568 65068 15620 65074
rect 15568 65010 15620 65016
rect 15476 64864 15528 64870
rect 15476 64806 15528 64812
rect 15108 64320 15160 64326
rect 15108 64262 15160 64268
rect 15016 63232 15068 63238
rect 15016 63174 15068 63180
rect 14924 61600 14976 61606
rect 14924 61542 14976 61548
rect 14832 59424 14884 59430
rect 14832 59366 14884 59372
rect 14936 57526 14964 61542
rect 14924 57520 14976 57526
rect 14924 57462 14976 57468
rect 14740 56364 14792 56370
rect 14740 56306 14792 56312
rect 14464 56296 14516 56302
rect 14464 56238 14516 56244
rect 14096 56160 14148 56166
rect 14096 56102 14148 56108
rect 14648 55072 14700 55078
rect 14648 55014 14700 55020
rect 14188 53100 14240 53106
rect 14188 53042 14240 53048
rect 13912 53032 13964 53038
rect 13912 52974 13964 52980
rect 13924 52698 13952 52974
rect 13544 52692 13596 52698
rect 13544 52634 13596 52640
rect 13912 52692 13964 52698
rect 13912 52634 13964 52640
rect 13556 44266 13584 52634
rect 14200 52630 14228 53042
rect 14280 52896 14332 52902
rect 14280 52838 14332 52844
rect 14188 52624 14240 52630
rect 14188 52566 14240 52572
rect 14292 52494 14320 52838
rect 14280 52488 14332 52494
rect 14280 52430 14332 52436
rect 14372 52352 14424 52358
rect 14372 52294 14424 52300
rect 14004 52080 14056 52086
rect 14004 52022 14056 52028
rect 13728 50856 13780 50862
rect 13728 50798 13780 50804
rect 13740 48890 13768 50798
rect 13728 48884 13780 48890
rect 13728 48826 13780 48832
rect 13912 48000 13964 48006
rect 13912 47942 13964 47948
rect 13924 47802 13952 47942
rect 13912 47796 13964 47802
rect 13912 47738 13964 47744
rect 14016 46374 14044 52022
rect 14384 51338 14412 52294
rect 14660 52086 14688 55014
rect 14832 52488 14884 52494
rect 14832 52430 14884 52436
rect 14648 52080 14700 52086
rect 14648 52022 14700 52028
rect 14464 52012 14516 52018
rect 14464 51954 14516 51960
rect 14476 51610 14504 51954
rect 14740 51944 14792 51950
rect 14740 51886 14792 51892
rect 14752 51610 14780 51886
rect 14464 51604 14516 51610
rect 14464 51546 14516 51552
rect 14740 51604 14792 51610
rect 14740 51546 14792 51552
rect 14648 51400 14700 51406
rect 14554 51368 14610 51377
rect 14372 51332 14424 51338
rect 14648 51342 14700 51348
rect 14554 51303 14610 51312
rect 14372 51274 14424 51280
rect 14384 50998 14412 51274
rect 14372 50992 14424 50998
rect 14372 50934 14424 50940
rect 14280 49836 14332 49842
rect 14280 49778 14332 49784
rect 14188 49768 14240 49774
rect 14188 49710 14240 49716
rect 14096 49700 14148 49706
rect 14096 49642 14148 49648
rect 14108 49434 14136 49642
rect 14096 49428 14148 49434
rect 14096 49370 14148 49376
rect 14096 49224 14148 49230
rect 14096 49166 14148 49172
rect 14108 47530 14136 49166
rect 14096 47524 14148 47530
rect 14096 47466 14148 47472
rect 14200 46714 14228 49710
rect 14292 49434 14320 49778
rect 14280 49428 14332 49434
rect 14280 49370 14332 49376
rect 14384 49314 14412 50934
rect 14568 49774 14596 51303
rect 14556 49768 14608 49774
rect 14556 49710 14608 49716
rect 14292 49286 14412 49314
rect 14292 48142 14320 49286
rect 14280 48136 14332 48142
rect 14280 48078 14332 48084
rect 14372 48136 14424 48142
rect 14372 48078 14424 48084
rect 14188 46708 14240 46714
rect 14188 46650 14240 46656
rect 13820 46368 13872 46374
rect 13820 46310 13872 46316
rect 14004 46368 14056 46374
rect 14004 46310 14056 46316
rect 13832 46034 13860 46310
rect 13820 46028 13872 46034
rect 13820 45970 13872 45976
rect 14004 45620 14056 45626
rect 14004 45562 14056 45568
rect 13728 45484 13780 45490
rect 13728 45426 13780 45432
rect 13544 44260 13596 44266
rect 13544 44202 13596 44208
rect 13556 39574 13584 44202
rect 13740 43994 13768 45426
rect 13912 44872 13964 44878
rect 13912 44814 13964 44820
rect 13728 43988 13780 43994
rect 13728 43930 13780 43936
rect 13924 39642 13952 44814
rect 14016 42838 14044 45562
rect 14188 45484 14240 45490
rect 14188 45426 14240 45432
rect 14200 44470 14228 45426
rect 14188 44464 14240 44470
rect 14188 44406 14240 44412
rect 14200 43790 14228 44406
rect 14188 43784 14240 43790
rect 14188 43726 14240 43732
rect 14096 43716 14148 43722
rect 14096 43658 14148 43664
rect 14108 43110 14136 43658
rect 14292 43178 14320 48078
rect 14384 47258 14412 48078
rect 14464 47660 14516 47666
rect 14464 47602 14516 47608
rect 14372 47252 14424 47258
rect 14372 47194 14424 47200
rect 14372 47048 14424 47054
rect 14372 46990 14424 46996
rect 14384 46102 14412 46990
rect 14476 46646 14504 47602
rect 14556 47592 14608 47598
rect 14556 47534 14608 47540
rect 14464 46640 14516 46646
rect 14464 46582 14516 46588
rect 14568 46510 14596 47534
rect 14660 47530 14688 51342
rect 14740 48612 14792 48618
rect 14740 48554 14792 48560
rect 14752 47734 14780 48554
rect 14740 47728 14792 47734
rect 14740 47670 14792 47676
rect 14648 47524 14700 47530
rect 14648 47466 14700 47472
rect 14648 47048 14700 47054
rect 14648 46990 14700 46996
rect 14556 46504 14608 46510
rect 14556 46446 14608 46452
rect 14372 46096 14424 46102
rect 14372 46038 14424 46044
rect 14568 43858 14596 46446
rect 14660 46170 14688 46990
rect 14740 46980 14792 46986
rect 14740 46922 14792 46928
rect 14752 46646 14780 46922
rect 14740 46640 14792 46646
rect 14740 46582 14792 46588
rect 14648 46164 14700 46170
rect 14648 46106 14700 46112
rect 14648 44736 14700 44742
rect 14648 44678 14700 44684
rect 14372 43852 14424 43858
rect 14372 43794 14424 43800
rect 14556 43852 14608 43858
rect 14556 43794 14608 43800
rect 14280 43172 14332 43178
rect 14280 43114 14332 43120
rect 14096 43104 14148 43110
rect 14096 43046 14148 43052
rect 14004 42832 14056 42838
rect 14004 42774 14056 42780
rect 14384 42702 14412 43794
rect 14464 43716 14516 43722
rect 14464 43658 14516 43664
rect 14372 42696 14424 42702
rect 14372 42638 14424 42644
rect 14476 42294 14504 43658
rect 14568 43382 14596 43794
rect 14660 43722 14688 44678
rect 14752 44538 14780 46582
rect 14844 46442 14872 52430
rect 14924 52420 14976 52426
rect 14924 52362 14976 52368
rect 14936 51406 14964 52362
rect 14924 51400 14976 51406
rect 14924 51342 14976 51348
rect 14936 51066 14964 51342
rect 14924 51060 14976 51066
rect 14924 51002 14976 51008
rect 14924 50924 14976 50930
rect 14924 50866 14976 50872
rect 14936 50182 14964 50866
rect 14924 50176 14976 50182
rect 14924 50118 14976 50124
rect 14924 48000 14976 48006
rect 14924 47942 14976 47948
rect 14936 47054 14964 47942
rect 14924 47048 14976 47054
rect 14924 46990 14976 46996
rect 14832 46436 14884 46442
rect 14832 46378 14884 46384
rect 15028 46186 15056 63174
rect 15120 62694 15148 64262
rect 15580 63986 15608 65010
rect 15846 64764 16154 64784
rect 15846 64762 15852 64764
rect 15908 64762 15932 64764
rect 15988 64762 16012 64764
rect 16068 64762 16092 64764
rect 16148 64762 16154 64764
rect 15908 64710 15910 64762
rect 16090 64710 16092 64762
rect 15846 64708 15852 64710
rect 15908 64708 15932 64710
rect 15988 64708 16012 64710
rect 16068 64708 16092 64710
rect 16148 64708 16154 64710
rect 15846 64688 16154 64708
rect 15568 63980 15620 63986
rect 15568 63922 15620 63928
rect 15580 63510 15608 63922
rect 15846 63676 16154 63696
rect 15846 63674 15852 63676
rect 15908 63674 15932 63676
rect 15988 63674 16012 63676
rect 16068 63674 16092 63676
rect 16148 63674 16154 63676
rect 15908 63622 15910 63674
rect 16090 63622 16092 63674
rect 15846 63620 15852 63622
rect 15908 63620 15932 63622
rect 15988 63620 16012 63622
rect 16068 63620 16092 63622
rect 16148 63620 16154 63622
rect 15846 63600 16154 63620
rect 15568 63504 15620 63510
rect 15568 63446 15620 63452
rect 15568 63368 15620 63374
rect 15568 63310 15620 63316
rect 15384 63300 15436 63306
rect 15384 63242 15436 63248
rect 15200 62756 15252 62762
rect 15200 62698 15252 62704
rect 15108 62688 15160 62694
rect 15108 62630 15160 62636
rect 15212 61810 15240 62698
rect 15200 61804 15252 61810
rect 15200 61746 15252 61752
rect 15212 61266 15240 61746
rect 15396 61402 15424 63242
rect 15580 61810 15608 63310
rect 15846 62588 16154 62608
rect 15846 62586 15852 62588
rect 15908 62586 15932 62588
rect 15988 62586 16012 62588
rect 16068 62586 16092 62588
rect 16148 62586 16154 62588
rect 15908 62534 15910 62586
rect 16090 62534 16092 62586
rect 15846 62532 15852 62534
rect 15908 62532 15932 62534
rect 15988 62532 16012 62534
rect 16068 62532 16092 62534
rect 16148 62532 16154 62534
rect 15846 62512 16154 62532
rect 16028 62416 16080 62422
rect 16028 62358 16080 62364
rect 16040 62286 16068 62358
rect 16028 62280 16080 62286
rect 16028 62222 16080 62228
rect 16212 62280 16264 62286
rect 16212 62222 16264 62228
rect 15568 61804 15620 61810
rect 15568 61746 15620 61752
rect 16224 61742 16252 62222
rect 16408 61826 16436 66558
rect 17132 66496 17184 66502
rect 17132 66438 17184 66444
rect 17144 66230 17172 66438
rect 17132 66224 17184 66230
rect 17132 66166 17184 66172
rect 16856 66156 16908 66162
rect 16856 66098 16908 66104
rect 16868 65754 16896 66098
rect 16856 65748 16908 65754
rect 16856 65690 16908 65696
rect 17328 65618 17356 68070
rect 17420 67726 17448 69702
rect 17512 68882 17540 69822
rect 17500 68876 17552 68882
rect 17500 68818 17552 68824
rect 17408 67720 17460 67726
rect 17408 67662 17460 67668
rect 17512 65618 17540 68818
rect 17592 67652 17644 67658
rect 17592 67594 17644 67600
rect 17316 65612 17368 65618
rect 17316 65554 17368 65560
rect 17500 65612 17552 65618
rect 17500 65554 17552 65560
rect 17512 65142 17540 65554
rect 17604 65414 17632 67594
rect 17684 67584 17736 67590
rect 17684 67526 17736 67532
rect 17696 66638 17724 67526
rect 17684 66632 17736 66638
rect 17684 66574 17736 66580
rect 17880 66570 17908 71470
rect 17960 71392 18012 71398
rect 17960 71334 18012 71340
rect 17972 69494 18000 71334
rect 18156 70650 18184 72218
rect 18248 71194 18276 72558
rect 18420 71528 18472 71534
rect 18418 71496 18420 71505
rect 19340 71528 19392 71534
rect 18472 71496 18474 71505
rect 19340 71470 19392 71476
rect 18418 71431 18474 71440
rect 18236 71188 18288 71194
rect 18236 71130 18288 71136
rect 18144 70644 18196 70650
rect 18144 70586 18196 70592
rect 18052 69828 18104 69834
rect 18052 69770 18104 69776
rect 17960 69488 18012 69494
rect 17960 69430 18012 69436
rect 17868 66564 17920 66570
rect 17868 66506 17920 66512
rect 17592 65408 17644 65414
rect 17592 65350 17644 65356
rect 17604 65210 17632 65350
rect 17592 65204 17644 65210
rect 17592 65146 17644 65152
rect 17500 65136 17552 65142
rect 17500 65078 17552 65084
rect 17132 65068 17184 65074
rect 17132 65010 17184 65016
rect 17144 63986 17172 65010
rect 17880 64874 17908 66506
rect 18064 65754 18092 69770
rect 18144 69352 18196 69358
rect 18144 69294 18196 69300
rect 18156 67930 18184 69294
rect 18248 68406 18276 71130
rect 18420 70916 18472 70922
rect 18420 70858 18472 70864
rect 18328 70644 18380 70650
rect 18328 70586 18380 70592
rect 18236 68400 18288 68406
rect 18236 68342 18288 68348
rect 18144 67924 18196 67930
rect 18144 67866 18196 67872
rect 18340 66706 18368 70586
rect 18432 66842 18460 70858
rect 18512 70100 18564 70106
rect 18512 70042 18564 70048
rect 18420 66836 18472 66842
rect 18420 66778 18472 66784
rect 18328 66700 18380 66706
rect 18328 66642 18380 66648
rect 18420 66496 18472 66502
rect 18420 66438 18472 66444
rect 18432 65958 18460 66438
rect 18524 66201 18552 70042
rect 19352 69222 19380 71470
rect 19524 71120 19576 71126
rect 19524 71062 19576 71068
rect 19536 70514 19564 71062
rect 19616 70916 19668 70922
rect 19616 70858 19668 70864
rect 19432 70508 19484 70514
rect 19432 70450 19484 70456
rect 19524 70508 19576 70514
rect 19524 70450 19576 70456
rect 19340 69216 19392 69222
rect 19340 69158 19392 69164
rect 18604 68740 18656 68746
rect 18604 68682 18656 68688
rect 18616 67386 18644 68682
rect 18696 67720 18748 67726
rect 18696 67662 18748 67668
rect 18604 67380 18656 67386
rect 18604 67322 18656 67328
rect 18708 67114 18736 67662
rect 18696 67108 18748 67114
rect 18696 67050 18748 67056
rect 18604 66632 18656 66638
rect 18604 66574 18656 66580
rect 18510 66192 18566 66201
rect 18510 66127 18566 66136
rect 18420 65952 18472 65958
rect 18420 65894 18472 65900
rect 18052 65748 18104 65754
rect 18052 65690 18104 65696
rect 18616 65074 18644 66574
rect 18696 66156 18748 66162
rect 18696 66098 18748 66104
rect 18708 65210 18736 66098
rect 19444 65754 19472 70450
rect 19524 69828 19576 69834
rect 19524 69770 19576 69776
rect 19536 68406 19564 69770
rect 19524 68400 19576 68406
rect 19524 68342 19576 68348
rect 19536 67318 19564 68342
rect 19524 67312 19576 67318
rect 19524 67254 19576 67260
rect 19628 66842 19656 70858
rect 19720 70650 19748 73034
rect 19800 71392 19852 71398
rect 19800 71334 19852 71340
rect 19708 70644 19760 70650
rect 19708 70586 19760 70592
rect 19708 70508 19760 70514
rect 19708 70450 19760 70456
rect 19720 69358 19748 70450
rect 19812 69834 19840 71334
rect 19904 69834 19932 73646
rect 20088 73574 20116 74598
rect 20444 74248 20496 74254
rect 20444 74190 20496 74196
rect 20456 73642 20484 74190
rect 20732 73760 20760 74870
rect 21284 74866 21312 75210
rect 21456 74996 21508 75002
rect 21456 74938 21508 74944
rect 21272 74860 21324 74866
rect 21272 74802 21324 74808
rect 21364 74860 21416 74866
rect 21364 74802 21416 74808
rect 21272 74656 21324 74662
rect 21272 74598 21324 74604
rect 21284 74254 21312 74598
rect 21180 74248 21232 74254
rect 21180 74190 21232 74196
rect 21272 74248 21324 74254
rect 21272 74190 21324 74196
rect 20811 74012 21119 74032
rect 20811 74010 20817 74012
rect 20873 74010 20897 74012
rect 20953 74010 20977 74012
rect 21033 74010 21057 74012
rect 21113 74010 21119 74012
rect 20873 73958 20875 74010
rect 21055 73958 21057 74010
rect 20811 73956 20817 73958
rect 20873 73956 20897 73958
rect 20953 73956 20977 73958
rect 21033 73956 21057 73958
rect 21113 73956 21119 73958
rect 20811 73936 21119 73956
rect 21088 73772 21140 73778
rect 20640 73732 21088 73760
rect 20444 73636 20496 73642
rect 20444 73578 20496 73584
rect 20076 73568 20128 73574
rect 20076 73510 20128 73516
rect 19984 70644 20036 70650
rect 19984 70586 20036 70592
rect 19800 69828 19852 69834
rect 19800 69770 19852 69776
rect 19892 69828 19944 69834
rect 19892 69770 19944 69776
rect 19708 69352 19760 69358
rect 19708 69294 19760 69300
rect 19708 69216 19760 69222
rect 19708 69158 19760 69164
rect 19720 67250 19748 69158
rect 19812 68746 19840 69770
rect 19800 68740 19852 68746
rect 19800 68682 19852 68688
rect 19708 67244 19760 67250
rect 19708 67186 19760 67192
rect 19904 67182 19932 69770
rect 19996 68814 20024 70586
rect 20088 70394 20116 73510
rect 20536 73160 20588 73166
rect 20536 73102 20588 73108
rect 20088 70366 20208 70394
rect 19984 68808 20036 68814
rect 19984 68750 20036 68756
rect 20076 68808 20128 68814
rect 20076 68750 20128 68756
rect 20088 68202 20116 68750
rect 20076 68196 20128 68202
rect 20076 68138 20128 68144
rect 19984 67652 20036 67658
rect 19984 67594 20036 67600
rect 19892 67176 19944 67182
rect 19892 67118 19944 67124
rect 19616 66836 19668 66842
rect 19616 66778 19668 66784
rect 19432 65748 19484 65754
rect 19432 65690 19484 65696
rect 19340 65544 19392 65550
rect 19340 65486 19392 65492
rect 18696 65204 18748 65210
rect 18696 65146 18748 65152
rect 18604 65068 18656 65074
rect 18604 65010 18656 65016
rect 17788 64846 17908 64874
rect 17132 63980 17184 63986
rect 17132 63922 17184 63928
rect 16580 63300 16632 63306
rect 16580 63242 16632 63248
rect 16488 62688 16540 62694
rect 16488 62630 16540 62636
rect 16500 62286 16528 62630
rect 16488 62280 16540 62286
rect 16488 62222 16540 62228
rect 16316 61798 16436 61826
rect 16592 61810 16620 63242
rect 16856 62348 16908 62354
rect 16856 62290 16908 62296
rect 16764 62212 16816 62218
rect 16764 62154 16816 62160
rect 16672 62144 16724 62150
rect 16672 62086 16724 62092
rect 16580 61804 16632 61810
rect 16212 61736 16264 61742
rect 16212 61678 16264 61684
rect 15846 61500 16154 61520
rect 15846 61498 15852 61500
rect 15908 61498 15932 61500
rect 15988 61498 16012 61500
rect 16068 61498 16092 61500
rect 16148 61498 16154 61500
rect 15908 61446 15910 61498
rect 16090 61446 16092 61498
rect 15846 61444 15852 61446
rect 15908 61444 15932 61446
rect 15988 61444 16012 61446
rect 16068 61444 16092 61446
rect 16148 61444 16154 61446
rect 15846 61424 16154 61444
rect 15384 61396 15436 61402
rect 16224 61384 16252 61678
rect 15384 61338 15436 61344
rect 16132 61356 16252 61384
rect 15200 61260 15252 61266
rect 15200 61202 15252 61208
rect 15660 61260 15712 61266
rect 15660 61202 15712 61208
rect 15476 60036 15528 60042
rect 15476 59978 15528 59984
rect 15108 57996 15160 58002
rect 15108 57938 15160 57944
rect 15120 51377 15148 57938
rect 15292 57860 15344 57866
rect 15292 57802 15344 57808
rect 15304 57594 15332 57802
rect 15292 57588 15344 57594
rect 15292 57530 15344 57536
rect 15384 57248 15436 57254
rect 15384 57190 15436 57196
rect 15396 56506 15424 57190
rect 15384 56500 15436 56506
rect 15384 56442 15436 56448
rect 15384 55956 15436 55962
rect 15384 55898 15436 55904
rect 15200 55888 15252 55894
rect 15200 55830 15252 55836
rect 15106 51368 15162 51377
rect 15106 51303 15162 51312
rect 15108 50924 15160 50930
rect 15108 50866 15160 50872
rect 15120 48074 15148 50866
rect 15212 48890 15240 55830
rect 15396 54754 15424 55898
rect 15488 54874 15516 59978
rect 15568 57792 15620 57798
rect 15568 57734 15620 57740
rect 15580 56370 15608 57734
rect 15672 57254 15700 61202
rect 16132 60858 16160 61356
rect 16212 61124 16264 61130
rect 16212 61066 16264 61072
rect 16120 60852 16172 60858
rect 16120 60794 16172 60800
rect 15752 60512 15804 60518
rect 15752 60454 15804 60460
rect 15764 60314 15792 60454
rect 15846 60412 16154 60432
rect 15846 60410 15852 60412
rect 15908 60410 15932 60412
rect 15988 60410 16012 60412
rect 16068 60410 16092 60412
rect 16148 60410 16154 60412
rect 15908 60358 15910 60410
rect 16090 60358 16092 60410
rect 15846 60356 15852 60358
rect 15908 60356 15932 60358
rect 15988 60356 16012 60358
rect 16068 60356 16092 60358
rect 16148 60356 16154 60358
rect 15846 60336 16154 60356
rect 15752 60308 15804 60314
rect 15752 60250 15804 60256
rect 15764 60042 15792 60250
rect 15752 60036 15804 60042
rect 15752 59978 15804 59984
rect 15846 59324 16154 59344
rect 15846 59322 15852 59324
rect 15908 59322 15932 59324
rect 15988 59322 16012 59324
rect 16068 59322 16092 59324
rect 16148 59322 16154 59324
rect 15908 59270 15910 59322
rect 16090 59270 16092 59322
rect 15846 59268 15852 59270
rect 15908 59268 15932 59270
rect 15988 59268 16012 59270
rect 16068 59268 16092 59270
rect 16148 59268 16154 59270
rect 15846 59248 16154 59268
rect 15846 58236 16154 58256
rect 15846 58234 15852 58236
rect 15908 58234 15932 58236
rect 15988 58234 16012 58236
rect 16068 58234 16092 58236
rect 16148 58234 16154 58236
rect 15908 58182 15910 58234
rect 16090 58182 16092 58234
rect 15846 58180 15852 58182
rect 15908 58180 15932 58182
rect 15988 58180 16012 58182
rect 16068 58180 16092 58182
rect 16148 58180 16154 58182
rect 15846 58160 16154 58180
rect 15660 57248 15712 57254
rect 15660 57190 15712 57196
rect 15568 56364 15620 56370
rect 15568 56306 15620 56312
rect 15476 54868 15528 54874
rect 15476 54810 15528 54816
rect 15396 54726 15516 54754
rect 15384 51400 15436 51406
rect 15384 51342 15436 51348
rect 15200 48884 15252 48890
rect 15200 48826 15252 48832
rect 15108 48068 15160 48074
rect 15108 48010 15160 48016
rect 14936 46158 15056 46186
rect 14740 44532 14792 44538
rect 14740 44474 14792 44480
rect 14648 43716 14700 43722
rect 14648 43658 14700 43664
rect 14556 43376 14608 43382
rect 14556 43318 14608 43324
rect 14464 42288 14516 42294
rect 14464 42230 14516 42236
rect 14568 42158 14596 43318
rect 14660 42362 14688 43658
rect 14648 42356 14700 42362
rect 14648 42298 14700 42304
rect 14280 42152 14332 42158
rect 14280 42094 14332 42100
rect 14556 42152 14608 42158
rect 14556 42094 14608 42100
rect 14096 42016 14148 42022
rect 14096 41958 14148 41964
rect 14108 41614 14136 41958
rect 14096 41608 14148 41614
rect 14096 41550 14148 41556
rect 14004 40384 14056 40390
rect 14004 40326 14056 40332
rect 13912 39636 13964 39642
rect 13912 39578 13964 39584
rect 13544 39568 13596 39574
rect 13544 39510 13596 39516
rect 13464 39086 13584 39114
rect 12992 38956 13044 38962
rect 12992 38898 13044 38904
rect 13004 38758 13032 38898
rect 13452 38820 13504 38826
rect 13452 38762 13504 38768
rect 12636 38678 12756 38706
rect 12992 38752 13044 38758
rect 12992 38694 13044 38700
rect 12636 38418 12664 38678
rect 12624 38412 12676 38418
rect 12624 38354 12676 38360
rect 12532 37392 12584 37398
rect 12532 37334 12584 37340
rect 12544 37262 12572 37334
rect 12532 37256 12584 37262
rect 12532 37198 12584 37204
rect 12636 37074 12664 38354
rect 12992 38276 13044 38282
rect 12992 38218 13044 38224
rect 13004 38010 13032 38218
rect 12716 38004 12768 38010
rect 12716 37946 12768 37952
rect 12992 38004 13044 38010
rect 12992 37946 13044 37952
rect 12728 37262 12756 37946
rect 12716 37256 12768 37262
rect 12716 37198 12768 37204
rect 12808 37120 12860 37126
rect 12636 37046 12756 37074
rect 12808 37062 12860 37068
rect 12348 35284 12400 35290
rect 12348 35226 12400 35232
rect 12624 35080 12676 35086
rect 12624 35022 12676 35028
rect 12348 33856 12400 33862
rect 12348 33798 12400 33804
rect 12072 33652 12124 33658
rect 12072 33594 12124 33600
rect 11796 32496 11848 32502
rect 11796 32438 11848 32444
rect 12360 32230 12388 33798
rect 12636 33386 12664 35022
rect 12624 33380 12676 33386
rect 12624 33322 12676 33328
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 11624 31726 11744 31754
rect 11428 30932 11480 30938
rect 11428 30874 11480 30880
rect 11244 30728 11296 30734
rect 11244 30670 11296 30676
rect 11244 30592 11296 30598
rect 11244 30534 11296 30540
rect 10880 30492 11188 30512
rect 10880 30490 10886 30492
rect 10942 30490 10966 30492
rect 11022 30490 11046 30492
rect 11102 30490 11126 30492
rect 11182 30490 11188 30492
rect 10942 30438 10944 30490
rect 11124 30438 11126 30490
rect 10880 30436 10886 30438
rect 10942 30436 10966 30438
rect 11022 30436 11046 30438
rect 11102 30436 11126 30438
rect 11182 30436 11188 30438
rect 10880 30416 11188 30436
rect 11256 30258 11284 30534
rect 11244 30252 11296 30258
rect 11244 30194 11296 30200
rect 11440 30190 11468 30874
rect 11624 30326 11652 31726
rect 12084 31482 12112 31826
rect 12360 31754 12388 32166
rect 12176 31726 12388 31754
rect 12176 31686 12204 31726
rect 12164 31680 12216 31686
rect 12164 31622 12216 31628
rect 12072 31476 12124 31482
rect 12072 31418 12124 31424
rect 11612 30320 11664 30326
rect 11612 30262 11664 30268
rect 11428 30184 11480 30190
rect 11428 30126 11480 30132
rect 12728 29646 12756 37046
rect 12820 31686 12848 37062
rect 13464 36922 13492 38762
rect 13556 37466 13584 39086
rect 14016 37942 14044 40326
rect 14292 39642 14320 42094
rect 14280 39636 14332 39642
rect 14280 39578 14332 39584
rect 14188 39364 14240 39370
rect 14188 39306 14240 39312
rect 14096 38888 14148 38894
rect 14096 38830 14148 38836
rect 14108 38729 14136 38830
rect 14094 38720 14150 38729
rect 14094 38655 14150 38664
rect 14096 38344 14148 38350
rect 14096 38286 14148 38292
rect 14004 37936 14056 37942
rect 14004 37878 14056 37884
rect 13728 37732 13780 37738
rect 13728 37674 13780 37680
rect 13544 37460 13596 37466
rect 13544 37402 13596 37408
rect 13740 37330 13768 37674
rect 13728 37324 13780 37330
rect 13728 37266 13780 37272
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13556 36786 13584 37062
rect 13740 36786 13768 37266
rect 13544 36780 13596 36786
rect 13544 36722 13596 36728
rect 13728 36780 13780 36786
rect 13728 36722 13780 36728
rect 13360 35488 13412 35494
rect 13360 35430 13412 35436
rect 13176 34672 13228 34678
rect 13176 34614 13228 34620
rect 12992 34604 13044 34610
rect 12992 34546 13044 34552
rect 13004 34134 13032 34546
rect 12992 34128 13044 34134
rect 12992 34070 13044 34076
rect 13084 34060 13136 34066
rect 13084 34002 13136 34008
rect 12992 33924 13044 33930
rect 12992 33866 13044 33872
rect 13004 33522 13032 33866
rect 12992 33516 13044 33522
rect 12992 33458 13044 33464
rect 12808 31680 12860 31686
rect 12808 31622 12860 31628
rect 12820 30394 12848 31622
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 10880 29404 11188 29424
rect 10880 29402 10886 29404
rect 10942 29402 10966 29404
rect 11022 29402 11046 29404
rect 11102 29402 11126 29404
rect 11182 29402 11188 29404
rect 10942 29350 10944 29402
rect 11124 29350 11126 29402
rect 10880 29348 10886 29350
rect 10942 29348 10966 29350
rect 11022 29348 11046 29350
rect 11102 29348 11126 29350
rect 11182 29348 11188 29350
rect 10880 29328 11188 29348
rect 12624 29164 12676 29170
rect 12624 29106 12676 29112
rect 12636 29073 12664 29106
rect 12622 29064 12678 29073
rect 12348 29028 12400 29034
rect 12622 28999 12678 29008
rect 12348 28970 12400 28976
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 9692 26206 9812 26234
rect 9692 19990 9720 26206
rect 10796 23866 10824 28426
rect 10880 28316 11188 28336
rect 10880 28314 10886 28316
rect 10942 28314 10966 28316
rect 11022 28314 11046 28316
rect 11102 28314 11126 28316
rect 11182 28314 11188 28316
rect 10942 28262 10944 28314
rect 11124 28262 11126 28314
rect 10880 28260 10886 28262
rect 10942 28260 10966 28262
rect 11022 28260 11046 28262
rect 11102 28260 11126 28262
rect 11182 28260 11188 28262
rect 10880 28240 11188 28260
rect 12360 27470 12388 28970
rect 12072 27464 12124 27470
rect 12072 27406 12124 27412
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 10880 27228 11188 27248
rect 10880 27226 10886 27228
rect 10942 27226 10966 27228
rect 11022 27226 11046 27228
rect 11102 27226 11126 27228
rect 11182 27226 11188 27228
rect 10942 27174 10944 27226
rect 11124 27174 11126 27226
rect 10880 27172 10886 27174
rect 10942 27172 10966 27174
rect 11022 27172 11046 27174
rect 11102 27172 11126 27174
rect 11182 27172 11188 27174
rect 10880 27152 11188 27172
rect 12084 27130 12112 27406
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 10880 26140 11188 26160
rect 10880 26138 10886 26140
rect 10942 26138 10966 26140
rect 11022 26138 11046 26140
rect 11102 26138 11126 26140
rect 11182 26138 11188 26140
rect 10942 26086 10944 26138
rect 11124 26086 11126 26138
rect 10880 26084 10886 26086
rect 10942 26084 10966 26086
rect 11022 26084 11046 26086
rect 11102 26084 11126 26086
rect 11182 26084 11188 26086
rect 10880 26064 11188 26084
rect 12544 25770 12572 26930
rect 12532 25764 12584 25770
rect 12532 25706 12584 25712
rect 10880 25052 11188 25072
rect 10880 25050 10886 25052
rect 10942 25050 10966 25052
rect 11022 25050 11046 25052
rect 11102 25050 11126 25052
rect 11182 25050 11188 25052
rect 10942 24998 10944 25050
rect 11124 24998 11126 25050
rect 10880 24996 10886 24998
rect 10942 24996 10966 24998
rect 11022 24996 11046 24998
rect 11102 24996 11126 24998
rect 11182 24996 11188 24998
rect 10880 24976 11188 24996
rect 10880 23964 11188 23984
rect 10880 23962 10886 23964
rect 10942 23962 10966 23964
rect 11022 23962 11046 23964
rect 11102 23962 11126 23964
rect 11182 23962 11188 23964
rect 10942 23910 10944 23962
rect 11124 23910 11126 23962
rect 10880 23908 10886 23910
rect 10942 23908 10966 23910
rect 11022 23908 11046 23910
rect 11102 23908 11126 23910
rect 11182 23908 11188 23910
rect 10880 23888 11188 23908
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10880 22876 11188 22896
rect 10880 22874 10886 22876
rect 10942 22874 10966 22876
rect 11022 22874 11046 22876
rect 11102 22874 11126 22876
rect 11182 22874 11188 22876
rect 10942 22822 10944 22874
rect 11124 22822 11126 22874
rect 10880 22820 10886 22822
rect 10942 22820 10966 22822
rect 11022 22820 11046 22822
rect 11102 22820 11126 22822
rect 11182 22820 11188 22822
rect 10880 22800 11188 22820
rect 10880 21788 11188 21808
rect 10880 21786 10886 21788
rect 10942 21786 10966 21788
rect 11022 21786 11046 21788
rect 11102 21786 11126 21788
rect 11182 21786 11188 21788
rect 10942 21734 10944 21786
rect 11124 21734 11126 21786
rect 10880 21732 10886 21734
rect 10942 21732 10966 21734
rect 11022 21732 11046 21734
rect 11102 21732 11126 21734
rect 11182 21732 11188 21734
rect 10880 21712 11188 21732
rect 12728 21146 12756 29582
rect 12806 29064 12862 29073
rect 12806 28999 12862 29008
rect 12820 27334 12848 28999
rect 12808 27328 12860 27334
rect 12808 27270 12860 27276
rect 13004 26602 13032 33458
rect 13096 33454 13124 34002
rect 13084 33448 13136 33454
rect 13084 33390 13136 33396
rect 13096 32026 13124 33390
rect 13188 32570 13216 34614
rect 13268 33584 13320 33590
rect 13268 33526 13320 33532
rect 13176 32564 13228 32570
rect 13176 32506 13228 32512
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 13188 31754 13216 32506
rect 13096 31726 13216 31754
rect 13096 31414 13124 31726
rect 13280 31482 13308 33526
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 13084 31408 13136 31414
rect 13084 31350 13136 31356
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13096 29646 13124 30126
rect 13084 29640 13136 29646
rect 13084 29582 13136 29588
rect 13096 29238 13124 29582
rect 13084 29232 13136 29238
rect 13084 29174 13136 29180
rect 13372 29170 13400 35430
rect 14108 35290 14136 38286
rect 14200 38010 14228 39306
rect 14188 38004 14240 38010
rect 14188 37946 14240 37952
rect 14556 38004 14608 38010
rect 14556 37946 14608 37952
rect 14096 35284 14148 35290
rect 14096 35226 14148 35232
rect 14568 35086 14596 37946
rect 14936 36582 14964 46158
rect 15016 43308 15068 43314
rect 15016 43250 15068 43256
rect 15028 42770 15056 43250
rect 15016 42764 15068 42770
rect 15016 42706 15068 42712
rect 15028 39438 15056 42706
rect 15120 42634 15148 48010
rect 15200 45892 15252 45898
rect 15200 45834 15252 45840
rect 15212 43994 15240 45834
rect 15292 44804 15344 44810
rect 15292 44746 15344 44752
rect 15200 43988 15252 43994
rect 15200 43930 15252 43936
rect 15200 43172 15252 43178
rect 15200 43114 15252 43120
rect 15212 42770 15240 43114
rect 15200 42764 15252 42770
rect 15200 42706 15252 42712
rect 15108 42628 15160 42634
rect 15108 42570 15160 42576
rect 15120 42362 15148 42570
rect 15108 42356 15160 42362
rect 15108 42298 15160 42304
rect 15304 41274 15332 44746
rect 15396 44266 15424 51342
rect 15488 51074 15516 54726
rect 15672 51074 15700 57190
rect 15846 57148 16154 57168
rect 15846 57146 15852 57148
rect 15908 57146 15932 57148
rect 15988 57146 16012 57148
rect 16068 57146 16092 57148
rect 16148 57146 16154 57148
rect 15908 57094 15910 57146
rect 16090 57094 16092 57146
rect 15846 57092 15852 57094
rect 15908 57092 15932 57094
rect 15988 57092 16012 57094
rect 16068 57092 16092 57094
rect 16148 57092 16154 57094
rect 15846 57072 16154 57092
rect 16224 57050 16252 61066
rect 16316 59702 16344 61798
rect 16580 61746 16632 61752
rect 16396 61396 16448 61402
rect 16396 61338 16448 61344
rect 16304 59696 16356 59702
rect 16304 59638 16356 59644
rect 16408 59022 16436 61338
rect 16684 60722 16712 62086
rect 16672 60716 16724 60722
rect 16672 60658 16724 60664
rect 16776 60058 16804 62154
rect 16868 61946 16896 62290
rect 16856 61940 16908 61946
rect 16856 61882 16908 61888
rect 16868 61266 16896 61882
rect 16856 61260 16908 61266
rect 16856 61202 16908 61208
rect 16948 61056 17000 61062
rect 16948 60998 17000 61004
rect 16856 60648 16908 60654
rect 16856 60590 16908 60596
rect 16684 60030 16804 60058
rect 16684 59974 16712 60030
rect 16672 59968 16724 59974
rect 16672 59910 16724 59916
rect 16396 59016 16448 59022
rect 16396 58958 16448 58964
rect 16684 58614 16712 59910
rect 16868 59770 16896 60590
rect 16856 59764 16908 59770
rect 16856 59706 16908 59712
rect 16764 59628 16816 59634
rect 16764 59570 16816 59576
rect 16672 58608 16724 58614
rect 16672 58550 16724 58556
rect 16776 58410 16804 59570
rect 16488 58404 16540 58410
rect 16488 58346 16540 58352
rect 16764 58404 16816 58410
rect 16764 58346 16816 58352
rect 16304 57860 16356 57866
rect 16304 57802 16356 57808
rect 16212 57044 16264 57050
rect 16212 56986 16264 56992
rect 16316 56250 16344 57802
rect 16500 57798 16528 58346
rect 16488 57792 16540 57798
rect 16488 57734 16540 57740
rect 16500 56438 16528 57734
rect 16488 56432 16540 56438
rect 16488 56374 16540 56380
rect 16960 56352 16988 60998
rect 16224 56222 16344 56250
rect 16868 56324 16988 56352
rect 15846 56060 16154 56080
rect 15846 56058 15852 56060
rect 15908 56058 15932 56060
rect 15988 56058 16012 56060
rect 16068 56058 16092 56060
rect 16148 56058 16154 56060
rect 15908 56006 15910 56058
rect 16090 56006 16092 56058
rect 15846 56004 15852 56006
rect 15908 56004 15932 56006
rect 15988 56004 16012 56006
rect 16068 56004 16092 56006
rect 16148 56004 16154 56006
rect 15846 55984 16154 56004
rect 16224 55826 16252 56222
rect 16304 55888 16356 55894
rect 16304 55830 16356 55836
rect 16212 55820 16264 55826
rect 16212 55762 16264 55768
rect 16224 55350 16252 55762
rect 16212 55344 16264 55350
rect 16212 55286 16264 55292
rect 15846 54972 16154 54992
rect 15846 54970 15852 54972
rect 15908 54970 15932 54972
rect 15988 54970 16012 54972
rect 16068 54970 16092 54972
rect 16148 54970 16154 54972
rect 15908 54918 15910 54970
rect 16090 54918 16092 54970
rect 15846 54916 15852 54918
rect 15908 54916 15932 54918
rect 15988 54916 16012 54918
rect 16068 54916 16092 54918
rect 16148 54916 16154 54918
rect 15846 54896 16154 54916
rect 16316 54670 16344 55830
rect 16580 55684 16632 55690
rect 16580 55626 16632 55632
rect 16592 55418 16620 55626
rect 16580 55412 16632 55418
rect 16580 55354 16632 55360
rect 16304 54664 16356 54670
rect 16304 54606 16356 54612
rect 16672 54528 16724 54534
rect 16672 54470 16724 54476
rect 16684 54194 16712 54470
rect 16868 54262 16896 56324
rect 16948 55684 17000 55690
rect 16948 55626 17000 55632
rect 16856 54256 16908 54262
rect 16856 54198 16908 54204
rect 16672 54188 16724 54194
rect 16672 54130 16724 54136
rect 15846 53884 16154 53904
rect 15846 53882 15852 53884
rect 15908 53882 15932 53884
rect 15988 53882 16012 53884
rect 16068 53882 16092 53884
rect 16148 53882 16154 53884
rect 15908 53830 15910 53882
rect 16090 53830 16092 53882
rect 15846 53828 15852 53830
rect 15908 53828 15932 53830
rect 15988 53828 16012 53830
rect 16068 53828 16092 53830
rect 16148 53828 16154 53830
rect 15846 53808 16154 53828
rect 15846 52796 16154 52816
rect 15846 52794 15852 52796
rect 15908 52794 15932 52796
rect 15988 52794 16012 52796
rect 16068 52794 16092 52796
rect 16148 52794 16154 52796
rect 15908 52742 15910 52794
rect 16090 52742 16092 52794
rect 15846 52740 15852 52742
rect 15908 52740 15932 52742
rect 15988 52740 16012 52742
rect 16068 52740 16092 52742
rect 16148 52740 16154 52742
rect 15846 52720 16154 52740
rect 16960 52154 16988 55626
rect 17144 55264 17172 63922
rect 17788 63510 17816 64846
rect 17960 63844 18012 63850
rect 17960 63786 18012 63792
rect 17776 63504 17828 63510
rect 17776 63446 17828 63452
rect 17868 63028 17920 63034
rect 17868 62970 17920 62976
rect 17880 62898 17908 62970
rect 17408 62892 17460 62898
rect 17868 62892 17920 62898
rect 17460 62852 17540 62880
rect 17408 62834 17460 62840
rect 17224 62824 17276 62830
rect 17224 62766 17276 62772
rect 17236 61742 17264 62766
rect 17316 62756 17368 62762
rect 17316 62698 17368 62704
rect 17328 62393 17356 62698
rect 17408 62688 17460 62694
rect 17408 62630 17460 62636
rect 17314 62384 17370 62393
rect 17314 62319 17370 62328
rect 17420 62286 17448 62630
rect 17316 62280 17368 62286
rect 17316 62222 17368 62228
rect 17408 62280 17460 62286
rect 17408 62222 17460 62228
rect 17224 61736 17276 61742
rect 17224 61678 17276 61684
rect 17328 60314 17356 62222
rect 17512 62150 17540 62852
rect 17868 62834 17920 62840
rect 17500 62144 17552 62150
rect 17500 62086 17552 62092
rect 17500 61736 17552 61742
rect 17500 61678 17552 61684
rect 17408 61192 17460 61198
rect 17408 61134 17460 61140
rect 17316 60308 17368 60314
rect 17316 60250 17368 60256
rect 17224 58880 17276 58886
rect 17224 58822 17276 58828
rect 17236 58478 17264 58822
rect 17224 58472 17276 58478
rect 17224 58414 17276 58420
rect 17316 58472 17368 58478
rect 17316 58414 17368 58420
rect 17236 57934 17264 58414
rect 17224 57928 17276 57934
rect 17224 57870 17276 57876
rect 17236 56914 17264 57870
rect 17328 57866 17356 58414
rect 17316 57860 17368 57866
rect 17316 57802 17368 57808
rect 17224 56908 17276 56914
rect 17224 56850 17276 56856
rect 17328 56778 17356 57802
rect 17316 56772 17368 56778
rect 17316 56714 17368 56720
rect 17328 55418 17356 56714
rect 17316 55412 17368 55418
rect 17316 55354 17368 55360
rect 17224 55276 17276 55282
rect 17144 55236 17224 55264
rect 17224 55218 17276 55224
rect 17040 54596 17092 54602
rect 17040 54538 17092 54544
rect 16948 52148 17000 52154
rect 16948 52090 17000 52096
rect 17052 52018 17080 54538
rect 17040 52012 17092 52018
rect 17040 51954 17092 51960
rect 15752 51808 15804 51814
rect 15752 51750 15804 51756
rect 15764 51474 15792 51750
rect 15846 51708 16154 51728
rect 15846 51706 15852 51708
rect 15908 51706 15932 51708
rect 15988 51706 16012 51708
rect 16068 51706 16092 51708
rect 16148 51706 16154 51708
rect 15908 51654 15910 51706
rect 16090 51654 16092 51706
rect 15846 51652 15852 51654
rect 15908 51652 15932 51654
rect 15988 51652 16012 51654
rect 16068 51652 16092 51654
rect 16148 51652 16154 51654
rect 15846 51632 16154 51652
rect 15752 51468 15804 51474
rect 15752 51410 15804 51416
rect 15488 51046 15608 51074
rect 15672 51046 16436 51074
rect 15476 50856 15528 50862
rect 15476 50798 15528 50804
rect 15488 50318 15516 50798
rect 15580 50794 15608 51046
rect 15568 50788 15620 50794
rect 15568 50730 15620 50736
rect 15752 50720 15804 50726
rect 15752 50662 15804 50668
rect 15476 50312 15528 50318
rect 15476 50254 15528 50260
rect 15660 50312 15712 50318
rect 15764 50300 15792 50662
rect 15846 50620 16154 50640
rect 15846 50618 15852 50620
rect 15908 50618 15932 50620
rect 15988 50618 16012 50620
rect 16068 50618 16092 50620
rect 16148 50618 16154 50620
rect 15908 50566 15910 50618
rect 16090 50566 16092 50618
rect 15846 50564 15852 50566
rect 15908 50564 15932 50566
rect 15988 50564 16012 50566
rect 16068 50564 16092 50566
rect 16148 50564 16154 50566
rect 15846 50544 16154 50564
rect 15844 50312 15896 50318
rect 15764 50272 15844 50300
rect 15660 50254 15712 50260
rect 15844 50254 15896 50260
rect 15672 49978 15700 50254
rect 15660 49972 15712 49978
rect 15660 49914 15712 49920
rect 15476 49836 15528 49842
rect 15476 49778 15528 49784
rect 15488 46442 15516 49778
rect 15846 49532 16154 49552
rect 15846 49530 15852 49532
rect 15908 49530 15932 49532
rect 15988 49530 16012 49532
rect 16068 49530 16092 49532
rect 16148 49530 16154 49532
rect 15908 49478 15910 49530
rect 16090 49478 16092 49530
rect 15846 49476 15852 49478
rect 15908 49476 15932 49478
rect 15988 49476 16012 49478
rect 16068 49476 16092 49478
rect 16148 49476 16154 49478
rect 15846 49456 16154 49476
rect 15752 48748 15804 48754
rect 15752 48690 15804 48696
rect 15568 46640 15620 46646
rect 15568 46582 15620 46588
rect 15476 46436 15528 46442
rect 15476 46378 15528 46384
rect 15476 44464 15528 44470
rect 15476 44406 15528 44412
rect 15384 44260 15436 44266
rect 15384 44202 15436 44208
rect 15488 43314 15516 44406
rect 15580 43722 15608 46582
rect 15660 46572 15712 46578
rect 15660 46514 15712 46520
rect 15672 44470 15700 46514
rect 15764 46050 15792 48690
rect 15846 48444 16154 48464
rect 15846 48442 15852 48444
rect 15908 48442 15932 48444
rect 15988 48442 16012 48444
rect 16068 48442 16092 48444
rect 16148 48442 16154 48444
rect 15908 48390 15910 48442
rect 16090 48390 16092 48442
rect 15846 48388 15852 48390
rect 15908 48388 15932 48390
rect 15988 48388 16012 48390
rect 16068 48388 16092 48390
rect 16148 48388 16154 48390
rect 15846 48368 16154 48388
rect 16212 48000 16264 48006
rect 16212 47942 16264 47948
rect 15846 47356 16154 47376
rect 15846 47354 15852 47356
rect 15908 47354 15932 47356
rect 15988 47354 16012 47356
rect 16068 47354 16092 47356
rect 16148 47354 16154 47356
rect 15908 47302 15910 47354
rect 16090 47302 16092 47354
rect 15846 47300 15852 47302
rect 15908 47300 15932 47302
rect 15988 47300 16012 47302
rect 16068 47300 16092 47302
rect 16148 47300 16154 47302
rect 15846 47280 16154 47300
rect 16224 46578 16252 47942
rect 16212 46572 16264 46578
rect 16212 46514 16264 46520
rect 16304 46504 16356 46510
rect 16304 46446 16356 46452
rect 15846 46268 16154 46288
rect 15846 46266 15852 46268
rect 15908 46266 15932 46268
rect 15988 46266 16012 46268
rect 16068 46266 16092 46268
rect 16148 46266 16154 46268
rect 15908 46214 15910 46266
rect 16090 46214 16092 46266
rect 15846 46212 15852 46214
rect 15908 46212 15932 46214
rect 15988 46212 16012 46214
rect 16068 46212 16092 46214
rect 16148 46212 16154 46214
rect 15846 46192 16154 46212
rect 15764 46022 15884 46050
rect 15752 45892 15804 45898
rect 15752 45834 15804 45840
rect 15764 45626 15792 45834
rect 15752 45620 15804 45626
rect 15752 45562 15804 45568
rect 15856 45506 15884 46022
rect 15764 45478 15884 45506
rect 15764 44742 15792 45478
rect 15846 45180 16154 45200
rect 15846 45178 15852 45180
rect 15908 45178 15932 45180
rect 15988 45178 16012 45180
rect 16068 45178 16092 45180
rect 16148 45178 16154 45180
rect 15908 45126 15910 45178
rect 16090 45126 16092 45178
rect 15846 45124 15852 45126
rect 15908 45124 15932 45126
rect 15988 45124 16012 45126
rect 16068 45124 16092 45126
rect 16148 45124 16154 45126
rect 15846 45104 16154 45124
rect 15752 44736 15804 44742
rect 15752 44678 15804 44684
rect 15660 44464 15712 44470
rect 15660 44406 15712 44412
rect 15568 43716 15620 43722
rect 15568 43658 15620 43664
rect 15476 43308 15528 43314
rect 15476 43250 15528 43256
rect 15488 42702 15516 43250
rect 15476 42696 15528 42702
rect 15476 42638 15528 42644
rect 15660 42696 15712 42702
rect 15660 42638 15712 42644
rect 15384 42560 15436 42566
rect 15384 42502 15436 42508
rect 15396 41614 15424 42502
rect 15672 41818 15700 42638
rect 15764 42294 15792 44678
rect 16316 44470 16344 46446
rect 16304 44464 16356 44470
rect 16304 44406 16356 44412
rect 15846 44092 16154 44112
rect 15846 44090 15852 44092
rect 15908 44090 15932 44092
rect 15988 44090 16012 44092
rect 16068 44090 16092 44092
rect 16148 44090 16154 44092
rect 15908 44038 15910 44090
rect 16090 44038 16092 44090
rect 15846 44036 15852 44038
rect 15908 44036 15932 44038
rect 15988 44036 16012 44038
rect 16068 44036 16092 44038
rect 16148 44036 16154 44038
rect 15846 44016 16154 44036
rect 16316 43790 16344 44406
rect 16408 43790 16436 51046
rect 16854 47832 16910 47841
rect 16854 47767 16910 47776
rect 16764 47660 16816 47666
rect 16764 47602 16816 47608
rect 16488 46708 16540 46714
rect 16488 46650 16540 46656
rect 16304 43784 16356 43790
rect 16304 43726 16356 43732
rect 16396 43784 16448 43790
rect 16396 43726 16448 43732
rect 16304 43308 16356 43314
rect 16304 43250 16356 43256
rect 16212 43104 16264 43110
rect 16212 43046 16264 43052
rect 15846 43004 16154 43024
rect 15846 43002 15852 43004
rect 15908 43002 15932 43004
rect 15988 43002 16012 43004
rect 16068 43002 16092 43004
rect 16148 43002 16154 43004
rect 15908 42950 15910 43002
rect 16090 42950 16092 43002
rect 15846 42948 15852 42950
rect 15908 42948 15932 42950
rect 15988 42948 16012 42950
rect 16068 42948 16092 42950
rect 16148 42948 16154 42950
rect 15846 42928 16154 42948
rect 15752 42288 15804 42294
rect 15752 42230 15804 42236
rect 15846 41916 16154 41936
rect 15846 41914 15852 41916
rect 15908 41914 15932 41916
rect 15988 41914 16012 41916
rect 16068 41914 16092 41916
rect 16148 41914 16154 41916
rect 15908 41862 15910 41914
rect 16090 41862 16092 41914
rect 15846 41860 15852 41862
rect 15908 41860 15932 41862
rect 15988 41860 16012 41862
rect 16068 41860 16092 41862
rect 16148 41860 16154 41862
rect 15846 41840 16154 41860
rect 15660 41812 15712 41818
rect 15660 41754 15712 41760
rect 15384 41608 15436 41614
rect 15384 41550 15436 41556
rect 15292 41268 15344 41274
rect 15292 41210 15344 41216
rect 15752 41064 15804 41070
rect 15752 41006 15804 41012
rect 15764 40526 15792 41006
rect 15846 40828 16154 40848
rect 15846 40826 15852 40828
rect 15908 40826 15932 40828
rect 15988 40826 16012 40828
rect 16068 40826 16092 40828
rect 16148 40826 16154 40828
rect 15908 40774 15910 40826
rect 16090 40774 16092 40826
rect 15846 40772 15852 40774
rect 15908 40772 15932 40774
rect 15988 40772 16012 40774
rect 16068 40772 16092 40774
rect 16148 40772 16154 40774
rect 15846 40752 16154 40772
rect 15752 40520 15804 40526
rect 15752 40462 15804 40468
rect 15752 40112 15804 40118
rect 15752 40054 15804 40060
rect 15016 39432 15068 39438
rect 15016 39374 15068 39380
rect 15384 39364 15436 39370
rect 15384 39306 15436 39312
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 15016 37188 15068 37194
rect 15016 37130 15068 37136
rect 15028 36922 15056 37130
rect 15016 36916 15068 36922
rect 15016 36858 15068 36864
rect 14924 36576 14976 36582
rect 14924 36518 14976 36524
rect 15212 36378 15240 37198
rect 15396 36961 15424 39306
rect 15660 39296 15712 39302
rect 15660 39238 15712 39244
rect 15568 38752 15620 38758
rect 15568 38694 15620 38700
rect 15476 38208 15528 38214
rect 15476 38150 15528 38156
rect 15488 37942 15516 38150
rect 15476 37936 15528 37942
rect 15476 37878 15528 37884
rect 15580 37194 15608 38694
rect 15672 38214 15700 39238
rect 15660 38208 15712 38214
rect 15660 38150 15712 38156
rect 15660 37664 15712 37670
rect 15660 37606 15712 37612
rect 15568 37188 15620 37194
rect 15568 37130 15620 37136
rect 15382 36952 15438 36961
rect 15382 36887 15438 36896
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15016 36168 15068 36174
rect 15016 36110 15068 36116
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14096 35012 14148 35018
rect 14096 34954 14148 34960
rect 13912 34740 13964 34746
rect 13912 34682 13964 34688
rect 13820 34468 13872 34474
rect 13820 34410 13872 34416
rect 13728 34128 13780 34134
rect 13728 34070 13780 34076
rect 13740 33930 13768 34070
rect 13832 33998 13860 34410
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 13728 33924 13780 33930
rect 13728 33866 13780 33872
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 13452 31136 13504 31142
rect 13452 31078 13504 31084
rect 13464 30394 13492 31078
rect 13452 30388 13504 30394
rect 13452 30330 13504 30336
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13556 28150 13584 33798
rect 13740 33658 13768 33866
rect 13728 33652 13780 33658
rect 13728 33594 13780 33600
rect 13636 32904 13688 32910
rect 13636 32846 13688 32852
rect 13648 32502 13676 32846
rect 13636 32496 13688 32502
rect 13636 32438 13688 32444
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 13636 30660 13688 30666
rect 13636 30602 13688 30608
rect 13648 28801 13676 30602
rect 13728 30320 13780 30326
rect 13728 30262 13780 30268
rect 13740 29170 13768 30262
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13634 28792 13690 28801
rect 13634 28727 13690 28736
rect 13832 28218 13860 31826
rect 13924 29238 13952 34682
rect 14108 34610 14136 34954
rect 14004 34604 14056 34610
rect 14004 34546 14056 34552
rect 14096 34604 14148 34610
rect 14096 34546 14148 34552
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14016 34202 14044 34546
rect 14004 34196 14056 34202
rect 14004 34138 14056 34144
rect 14108 31822 14136 34546
rect 14752 33386 14780 34546
rect 14924 34400 14976 34406
rect 14924 34342 14976 34348
rect 14740 33380 14792 33386
rect 14740 33322 14792 33328
rect 14372 33108 14424 33114
rect 14372 33050 14424 33056
rect 14280 32836 14332 32842
rect 14280 32778 14332 32784
rect 14292 32026 14320 32778
rect 14384 32434 14412 33050
rect 14936 32910 14964 34342
rect 15028 33386 15056 36110
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 15120 33998 15148 35022
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15016 33380 15068 33386
rect 15016 33322 15068 33328
rect 14924 32904 14976 32910
rect 14924 32846 14976 32852
rect 14464 32836 14516 32842
rect 14464 32778 14516 32784
rect 14476 32570 14504 32778
rect 14740 32768 14792 32774
rect 14740 32710 14792 32716
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14752 32434 14780 32710
rect 15120 32434 15148 33934
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 14372 32428 14424 32434
rect 14556 32428 14608 32434
rect 14372 32370 14424 32376
rect 14464 32412 14516 32418
rect 14556 32370 14608 32376
rect 14740 32428 14792 32434
rect 14740 32370 14792 32376
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 14464 32354 14516 32360
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14096 31816 14148 31822
rect 14096 31758 14148 31764
rect 14004 31476 14056 31482
rect 14004 31418 14056 31424
rect 14016 30258 14044 31418
rect 14188 31136 14240 31142
rect 14188 31078 14240 31084
rect 14200 30258 14228 31078
rect 14476 30326 14504 32354
rect 14568 31482 14596 32370
rect 15016 31748 15068 31754
rect 15016 31690 15068 31696
rect 15028 31482 15056 31690
rect 14556 31476 14608 31482
rect 14556 31418 14608 31424
rect 15016 31476 15068 31482
rect 15016 31418 15068 31424
rect 15108 31340 15160 31346
rect 15108 31282 15160 31288
rect 14740 30388 14792 30394
rect 14740 30330 14792 30336
rect 14464 30320 14516 30326
rect 14464 30262 14516 30268
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 14004 30048 14056 30054
rect 14004 29990 14056 29996
rect 13912 29232 13964 29238
rect 13912 29174 13964 29180
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 13544 28144 13596 28150
rect 13544 28086 13596 28092
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13004 26574 13124 26602
rect 12992 26240 13044 26246
rect 12992 26182 13044 26188
rect 13004 25838 13032 26182
rect 13096 25906 13124 26574
rect 13648 26042 13676 26726
rect 13832 26382 13860 28154
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 13636 26036 13688 26042
rect 13636 25978 13688 25984
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 13004 24886 13032 25774
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 13004 24206 13032 24822
rect 13096 24750 13124 25842
rect 13280 24954 13308 25978
rect 13268 24948 13320 24954
rect 13268 24890 13320 24896
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13188 23730 13216 24278
rect 13280 24138 13308 24890
rect 14016 24818 14044 29990
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14188 29504 14240 29510
rect 14188 29446 14240 29452
rect 14004 24812 14056 24818
rect 14004 24754 14056 24760
rect 13452 24744 13504 24750
rect 13452 24686 13504 24692
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13464 24206 13492 24686
rect 13924 24410 13952 24686
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 14108 24206 14136 24550
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13004 23322 13032 23666
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 14108 23186 14136 23462
rect 14096 23180 14148 23186
rect 14096 23122 14148 23128
rect 14200 23118 14228 29446
rect 14384 28257 14412 29582
rect 14476 29510 14504 30262
rect 14648 30184 14700 30190
rect 14648 30126 14700 30132
rect 14660 29646 14688 30126
rect 14752 29646 14780 30330
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14476 28694 14504 29446
rect 14660 29102 14688 29582
rect 15120 29306 15148 31282
rect 15212 31142 15240 33390
rect 15292 31680 15344 31686
rect 15292 31622 15344 31628
rect 15200 31136 15252 31142
rect 15200 31078 15252 31084
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15108 29300 15160 29306
rect 15108 29242 15160 29248
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14464 28688 14516 28694
rect 14464 28630 14516 28636
rect 14660 28626 14688 29038
rect 14738 28792 14794 28801
rect 14738 28727 14794 28736
rect 14648 28620 14700 28626
rect 14648 28562 14700 28568
rect 14752 28558 14780 28727
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14370 28248 14426 28257
rect 14370 28183 14426 28192
rect 15016 27056 15068 27062
rect 15120 27044 15148 29242
rect 15068 27016 15148 27044
rect 15016 26998 15068 27004
rect 15212 26382 15240 30534
rect 15304 28994 15332 31622
rect 15396 31414 15424 36887
rect 15476 36780 15528 36786
rect 15528 36740 15608 36768
rect 15476 36722 15528 36728
rect 15476 35624 15528 35630
rect 15476 35566 15528 35572
rect 15384 31408 15436 31414
rect 15384 31350 15436 31356
rect 15488 30598 15516 35566
rect 15580 32026 15608 36740
rect 15568 32020 15620 32026
rect 15568 31962 15620 31968
rect 15672 31754 15700 37606
rect 15764 36378 15792 40054
rect 15846 39740 16154 39760
rect 15846 39738 15852 39740
rect 15908 39738 15932 39740
rect 15988 39738 16012 39740
rect 16068 39738 16092 39740
rect 16148 39738 16154 39740
rect 15908 39686 15910 39738
rect 16090 39686 16092 39738
rect 15846 39684 15852 39686
rect 15908 39684 15932 39686
rect 15988 39684 16012 39686
rect 16068 39684 16092 39686
rect 16148 39684 16154 39686
rect 15846 39664 16154 39684
rect 16224 38842 16252 43046
rect 16316 38962 16344 43250
rect 16396 42560 16448 42566
rect 16396 42502 16448 42508
rect 16408 41206 16436 42502
rect 16396 41200 16448 41206
rect 16396 41142 16448 41148
rect 16304 38956 16356 38962
rect 16304 38898 16356 38904
rect 16224 38814 16344 38842
rect 15846 38652 16154 38672
rect 15846 38650 15852 38652
rect 15908 38650 15932 38652
rect 15988 38650 16012 38652
rect 16068 38650 16092 38652
rect 16148 38650 16154 38652
rect 15908 38598 15910 38650
rect 16090 38598 16092 38650
rect 15846 38596 15852 38598
rect 15908 38596 15932 38598
rect 15988 38596 16012 38598
rect 16068 38596 16092 38598
rect 16148 38596 16154 38598
rect 15846 38576 16154 38596
rect 16212 38412 16264 38418
rect 16212 38354 16264 38360
rect 16224 37670 16252 38354
rect 16212 37664 16264 37670
rect 16212 37606 16264 37612
rect 15846 37564 16154 37584
rect 15846 37562 15852 37564
rect 15908 37562 15932 37564
rect 15988 37562 16012 37564
rect 16068 37562 16092 37564
rect 16148 37562 16154 37564
rect 15908 37510 15910 37562
rect 16090 37510 16092 37562
rect 15846 37508 15852 37510
rect 15908 37508 15932 37510
rect 15988 37508 16012 37510
rect 16068 37508 16092 37510
rect 16148 37508 16154 37510
rect 15846 37488 16154 37508
rect 15934 36952 15990 36961
rect 15934 36887 15990 36896
rect 15948 36854 15976 36887
rect 15936 36848 15988 36854
rect 15936 36790 15988 36796
rect 15844 36780 15896 36786
rect 15844 36722 15896 36728
rect 15856 36689 15884 36722
rect 16316 36718 16344 38814
rect 16500 38486 16528 46650
rect 16776 45082 16804 47602
rect 16764 45076 16816 45082
rect 16764 45018 16816 45024
rect 16580 44260 16632 44266
rect 16580 44202 16632 44208
rect 16592 43994 16620 44202
rect 16868 44146 16896 47767
rect 17052 47190 17080 51954
rect 17236 51338 17264 55218
rect 17420 54806 17448 61134
rect 17512 61130 17540 61678
rect 17972 61198 18000 63786
rect 18420 62824 18472 62830
rect 18420 62766 18472 62772
rect 18328 62484 18380 62490
rect 18328 62426 18380 62432
rect 18340 61266 18368 62426
rect 18328 61260 18380 61266
rect 18328 61202 18380 61208
rect 17960 61192 18012 61198
rect 17960 61134 18012 61140
rect 17500 61124 17552 61130
rect 17500 61066 17552 61072
rect 18340 60858 18368 61202
rect 18328 60852 18380 60858
rect 18328 60794 18380 60800
rect 17868 60784 17920 60790
rect 17868 60726 17920 60732
rect 17684 60104 17736 60110
rect 17684 60046 17736 60052
rect 17592 58608 17644 58614
rect 17592 58550 17644 58556
rect 17604 57798 17632 58550
rect 17592 57792 17644 57798
rect 17592 57734 17644 57740
rect 17500 56908 17552 56914
rect 17500 56850 17552 56856
rect 17512 56352 17540 56850
rect 17604 56710 17632 57734
rect 17696 57050 17724 60046
rect 17880 58002 17908 60726
rect 18432 60654 18460 62766
rect 18512 61736 18564 61742
rect 18512 61678 18564 61684
rect 18524 61402 18552 61678
rect 18512 61396 18564 61402
rect 18512 61338 18564 61344
rect 18512 61192 18564 61198
rect 18512 61134 18564 61140
rect 18420 60648 18472 60654
rect 18420 60590 18472 60596
rect 18328 58948 18380 58954
rect 18328 58890 18380 58896
rect 17868 57996 17920 58002
rect 17868 57938 17920 57944
rect 17868 57860 17920 57866
rect 17868 57802 17920 57808
rect 18236 57860 18288 57866
rect 18236 57802 18288 57808
rect 17684 57044 17736 57050
rect 17684 56986 17736 56992
rect 17880 56914 17908 57802
rect 17960 57452 18012 57458
rect 17960 57394 18012 57400
rect 17868 56908 17920 56914
rect 17868 56850 17920 56856
rect 17684 56840 17736 56846
rect 17684 56782 17736 56788
rect 17592 56704 17644 56710
rect 17592 56646 17644 56652
rect 17592 56364 17644 56370
rect 17512 56324 17592 56352
rect 17408 54800 17460 54806
rect 17408 54742 17460 54748
rect 17420 54330 17448 54742
rect 17408 54324 17460 54330
rect 17408 54266 17460 54272
rect 17224 51332 17276 51338
rect 17224 51274 17276 51280
rect 17512 51074 17540 56324
rect 17592 56306 17644 56312
rect 17696 55282 17724 56782
rect 17776 55616 17828 55622
rect 17776 55558 17828 55564
rect 17684 55276 17736 55282
rect 17684 55218 17736 55224
rect 17696 51406 17724 55218
rect 17788 53242 17816 55558
rect 17972 55418 18000 57394
rect 18052 56160 18104 56166
rect 18052 56102 18104 56108
rect 17960 55412 18012 55418
rect 17960 55354 18012 55360
rect 18064 53786 18092 56102
rect 18248 55622 18276 57802
rect 18340 57254 18368 58890
rect 18524 58138 18552 61134
rect 18616 59226 18644 65010
rect 19352 64462 19380 65486
rect 19996 64666 20024 67594
rect 20076 67176 20128 67182
rect 20076 67118 20128 67124
rect 20088 64666 20116 67118
rect 20180 66706 20208 70366
rect 20444 69420 20496 69426
rect 20444 69362 20496 69368
rect 20260 69352 20312 69358
rect 20260 69294 20312 69300
rect 20272 68218 20300 69294
rect 20456 68921 20484 69362
rect 20548 69018 20576 73102
rect 20640 69494 20668 73732
rect 21088 73714 21140 73720
rect 21192 73370 21220 74190
rect 21376 73914 21404 74802
rect 21364 73908 21416 73914
rect 21364 73850 21416 73856
rect 21468 73778 21496 74938
rect 21560 74798 21588 75822
rect 25776 75644 26084 75664
rect 25776 75642 25782 75644
rect 25838 75642 25862 75644
rect 25918 75642 25942 75644
rect 25998 75642 26022 75644
rect 26078 75642 26084 75644
rect 25838 75590 25840 75642
rect 26020 75590 26022 75642
rect 25776 75588 25782 75590
rect 25838 75588 25862 75590
rect 25918 75588 25942 75590
rect 25998 75588 26022 75590
rect 26078 75588 26084 75590
rect 25776 75568 26084 75588
rect 22376 75472 22428 75478
rect 22376 75414 22428 75420
rect 21548 74792 21600 74798
rect 21548 74734 21600 74740
rect 21824 74792 21876 74798
rect 21824 74734 21876 74740
rect 21456 73772 21508 73778
rect 21456 73714 21508 73720
rect 21560 73710 21588 74734
rect 21836 74458 21864 74734
rect 21824 74452 21876 74458
rect 21824 74394 21876 74400
rect 21364 73704 21416 73710
rect 21364 73646 21416 73652
rect 21548 73704 21600 73710
rect 21548 73646 21600 73652
rect 21180 73364 21232 73370
rect 21180 73306 21232 73312
rect 20720 73024 20772 73030
rect 20720 72966 20772 72972
rect 20732 71194 20760 72966
rect 20811 72924 21119 72944
rect 20811 72922 20817 72924
rect 20873 72922 20897 72924
rect 20953 72922 20977 72924
rect 21033 72922 21057 72924
rect 21113 72922 21119 72924
rect 20873 72870 20875 72922
rect 21055 72870 21057 72922
rect 20811 72868 20817 72870
rect 20873 72868 20897 72870
rect 20953 72868 20977 72870
rect 21033 72868 21057 72870
rect 21113 72868 21119 72870
rect 20811 72848 21119 72868
rect 20811 71836 21119 71856
rect 20811 71834 20817 71836
rect 20873 71834 20897 71836
rect 20953 71834 20977 71836
rect 21033 71834 21057 71836
rect 21113 71834 21119 71836
rect 20873 71782 20875 71834
rect 21055 71782 21057 71834
rect 20811 71780 20817 71782
rect 20873 71780 20897 71782
rect 20953 71780 20977 71782
rect 21033 71780 21057 71782
rect 21113 71780 21119 71782
rect 20811 71760 21119 71780
rect 21272 71664 21324 71670
rect 21272 71606 21324 71612
rect 20720 71188 20772 71194
rect 20720 71130 20772 71136
rect 20628 69488 20680 69494
rect 20628 69430 20680 69436
rect 20536 69012 20588 69018
rect 20536 68954 20588 68960
rect 20442 68912 20498 68921
rect 20352 68876 20404 68882
rect 20442 68847 20498 68856
rect 20352 68818 20404 68824
rect 20364 68406 20392 68818
rect 20444 68740 20496 68746
rect 20444 68682 20496 68688
rect 20536 68740 20588 68746
rect 20536 68682 20588 68688
rect 20456 68474 20484 68682
rect 20444 68468 20496 68474
rect 20444 68410 20496 68416
rect 20352 68400 20404 68406
rect 20352 68342 20404 68348
rect 20442 68368 20498 68377
rect 20442 68303 20498 68312
rect 20272 68190 20392 68218
rect 20168 66700 20220 66706
rect 20168 66642 20220 66648
rect 20260 65476 20312 65482
rect 20260 65418 20312 65424
rect 20272 65074 20300 65418
rect 20260 65068 20312 65074
rect 20260 65010 20312 65016
rect 19984 64660 20036 64666
rect 19984 64602 20036 64608
rect 20076 64660 20128 64666
rect 20076 64602 20128 64608
rect 19340 64456 19392 64462
rect 19340 64398 19392 64404
rect 18696 62144 18748 62150
rect 18696 62086 18748 62092
rect 18880 62144 18932 62150
rect 18880 62086 18932 62092
rect 18708 60586 18736 62086
rect 18788 61804 18840 61810
rect 18788 61746 18840 61752
rect 18800 60858 18828 61746
rect 18788 60852 18840 60858
rect 18788 60794 18840 60800
rect 18892 60734 18920 62086
rect 19156 61600 19208 61606
rect 19156 61542 19208 61548
rect 18970 61160 19026 61169
rect 18970 61095 19026 61104
rect 18984 60790 19012 61095
rect 18800 60706 18920 60734
rect 18972 60784 19024 60790
rect 18972 60726 19024 60732
rect 19064 60716 19116 60722
rect 18696 60580 18748 60586
rect 18696 60522 18748 60528
rect 18604 59220 18656 59226
rect 18604 59162 18656 59168
rect 18512 58132 18564 58138
rect 18512 58074 18564 58080
rect 18328 57248 18380 57254
rect 18328 57190 18380 57196
rect 18420 57248 18472 57254
rect 18420 57190 18472 57196
rect 18236 55616 18288 55622
rect 18236 55558 18288 55564
rect 18052 53780 18104 53786
rect 18052 53722 18104 53728
rect 17868 53576 17920 53582
rect 17868 53518 17920 53524
rect 17776 53236 17828 53242
rect 17776 53178 17828 53184
rect 17788 52426 17816 53178
rect 17880 52698 17908 53518
rect 18248 53174 18276 55558
rect 18340 55350 18368 57190
rect 18432 56438 18460 57190
rect 18420 56432 18472 56438
rect 18420 56374 18472 56380
rect 18696 55752 18748 55758
rect 18696 55694 18748 55700
rect 18328 55344 18380 55350
rect 18328 55286 18380 55292
rect 18708 53786 18736 55694
rect 18800 55078 18828 60706
rect 19168 60704 19196 61542
rect 19116 60676 19196 60704
rect 19064 60658 19116 60664
rect 19352 60636 19380 64398
rect 20272 64054 20300 65010
rect 20364 64530 20392 68190
rect 20456 65634 20484 68303
rect 20548 68270 20576 68682
rect 20628 68672 20680 68678
rect 20628 68614 20680 68620
rect 20536 68264 20588 68270
rect 20536 68206 20588 68212
rect 20536 66632 20588 66638
rect 20536 66574 20588 66580
rect 20548 65754 20576 66574
rect 20640 66026 20668 68614
rect 20732 68338 20760 71130
rect 20811 70748 21119 70768
rect 20811 70746 20817 70748
rect 20873 70746 20897 70748
rect 20953 70746 20977 70748
rect 21033 70746 21057 70748
rect 21113 70746 21119 70748
rect 20873 70694 20875 70746
rect 21055 70694 21057 70746
rect 20811 70692 20817 70694
rect 20873 70692 20897 70694
rect 20953 70692 20977 70694
rect 21033 70692 21057 70694
rect 21113 70692 21119 70694
rect 20811 70672 21119 70692
rect 20812 70508 20864 70514
rect 20812 70450 20864 70456
rect 20824 70106 20852 70450
rect 21088 70304 21140 70310
rect 21088 70246 21140 70252
rect 20812 70100 20864 70106
rect 20812 70042 20864 70048
rect 21100 69902 21128 70246
rect 21088 69896 21140 69902
rect 21088 69838 21140 69844
rect 20811 69660 21119 69680
rect 20811 69658 20817 69660
rect 20873 69658 20897 69660
rect 20953 69658 20977 69660
rect 21033 69658 21057 69660
rect 21113 69658 21119 69660
rect 20873 69606 20875 69658
rect 21055 69606 21057 69658
rect 20811 69604 20817 69606
rect 20873 69604 20897 69606
rect 20953 69604 20977 69606
rect 21033 69604 21057 69606
rect 21113 69604 21119 69606
rect 20811 69584 21119 69604
rect 20811 68572 21119 68592
rect 20811 68570 20817 68572
rect 20873 68570 20897 68572
rect 20953 68570 20977 68572
rect 21033 68570 21057 68572
rect 21113 68570 21119 68572
rect 20873 68518 20875 68570
rect 21055 68518 21057 68570
rect 20811 68516 20817 68518
rect 20873 68516 20897 68518
rect 20953 68516 20977 68518
rect 21033 68516 21057 68518
rect 21113 68516 21119 68518
rect 20811 68496 21119 68516
rect 20720 68332 20772 68338
rect 20720 68274 20772 68280
rect 21180 68264 21232 68270
rect 21180 68206 21232 68212
rect 20811 67484 21119 67504
rect 20811 67482 20817 67484
rect 20873 67482 20897 67484
rect 20953 67482 20977 67484
rect 21033 67482 21057 67484
rect 21113 67482 21119 67484
rect 20873 67430 20875 67482
rect 21055 67430 21057 67482
rect 20811 67428 20817 67430
rect 20873 67428 20897 67430
rect 20953 67428 20977 67430
rect 21033 67428 21057 67430
rect 21113 67428 21119 67430
rect 20811 67408 21119 67428
rect 20720 66496 20772 66502
rect 20720 66438 20772 66444
rect 20628 66020 20680 66026
rect 20628 65962 20680 65968
rect 20536 65748 20588 65754
rect 20536 65690 20588 65696
rect 20456 65606 20576 65634
rect 20444 65408 20496 65414
rect 20444 65350 20496 65356
rect 20456 65142 20484 65350
rect 20444 65136 20496 65142
rect 20444 65078 20496 65084
rect 20548 64954 20576 65606
rect 20456 64926 20576 64954
rect 20352 64524 20404 64530
rect 20352 64466 20404 64472
rect 20260 64048 20312 64054
rect 20260 63990 20312 63996
rect 20272 63442 20300 63990
rect 20456 63866 20484 64926
rect 20536 64388 20588 64394
rect 20536 64330 20588 64336
rect 20548 63986 20576 64330
rect 20640 64122 20668 65962
rect 20732 65618 20760 66438
rect 20811 66396 21119 66416
rect 20811 66394 20817 66396
rect 20873 66394 20897 66396
rect 20953 66394 20977 66396
rect 21033 66394 21057 66396
rect 21113 66394 21119 66396
rect 20873 66342 20875 66394
rect 21055 66342 21057 66394
rect 20811 66340 20817 66342
rect 20873 66340 20897 66342
rect 20953 66340 20977 66342
rect 21033 66340 21057 66342
rect 21113 66340 21119 66342
rect 20811 66320 21119 66340
rect 21192 65686 21220 68206
rect 21284 67862 21312 71606
rect 21376 71398 21404 73646
rect 21456 71596 21508 71602
rect 21456 71538 21508 71544
rect 21364 71392 21416 71398
rect 21364 71334 21416 71340
rect 21376 70446 21404 71334
rect 21364 70440 21416 70446
rect 21364 70382 21416 70388
rect 21468 69426 21496 71538
rect 22388 70582 22416 75414
rect 24952 75200 25004 75206
rect 24952 75142 25004 75148
rect 22560 74656 22612 74662
rect 22560 74598 22612 74604
rect 22836 74656 22888 74662
rect 22836 74598 22888 74604
rect 22572 74534 22600 74598
rect 22572 74506 22692 74534
rect 22664 74118 22692 74506
rect 22652 74112 22704 74118
rect 22652 74054 22704 74060
rect 22468 71460 22520 71466
rect 22468 71402 22520 71408
rect 22376 70576 22428 70582
rect 22376 70518 22428 70524
rect 22008 70508 22060 70514
rect 22008 70450 22060 70456
rect 22284 70508 22336 70514
rect 22284 70450 22336 70456
rect 21824 70304 21876 70310
rect 21824 70246 21876 70252
rect 21836 69834 21864 70246
rect 22020 70106 22048 70450
rect 22296 70394 22324 70450
rect 22296 70366 22416 70394
rect 22008 70100 22060 70106
rect 22008 70042 22060 70048
rect 22284 69896 22336 69902
rect 22284 69838 22336 69844
rect 21824 69828 21876 69834
rect 21824 69770 21876 69776
rect 21916 69828 21968 69834
rect 21916 69770 21968 69776
rect 21928 69562 21956 69770
rect 22100 69760 22152 69766
rect 22100 69702 22152 69708
rect 21916 69556 21968 69562
rect 21916 69498 21968 69504
rect 22112 69426 22140 69702
rect 21456 69420 21508 69426
rect 21456 69362 21508 69368
rect 22100 69420 22152 69426
rect 22100 69362 22152 69368
rect 21272 67856 21324 67862
rect 21272 67798 21324 67804
rect 20812 65680 20864 65686
rect 20812 65622 20864 65628
rect 21180 65680 21232 65686
rect 21180 65622 21232 65628
rect 20720 65612 20772 65618
rect 20720 65554 20772 65560
rect 20824 65498 20852 65622
rect 20732 65470 20852 65498
rect 21180 65476 21232 65482
rect 20732 65142 20760 65470
rect 21180 65418 21232 65424
rect 20811 65308 21119 65328
rect 20811 65306 20817 65308
rect 20873 65306 20897 65308
rect 20953 65306 20977 65308
rect 21033 65306 21057 65308
rect 21113 65306 21119 65308
rect 20873 65254 20875 65306
rect 21055 65254 21057 65306
rect 20811 65252 20817 65254
rect 20873 65252 20897 65254
rect 20953 65252 20977 65254
rect 21033 65252 21057 65254
rect 21113 65252 21119 65254
rect 20811 65232 21119 65252
rect 20720 65136 20772 65142
rect 20720 65078 20772 65084
rect 20628 64116 20680 64122
rect 20628 64058 20680 64064
rect 20732 64054 20760 65078
rect 21192 64666 21220 65418
rect 21284 65210 21312 67798
rect 21468 66254 21496 69362
rect 22192 69284 22244 69290
rect 22192 69226 22244 69232
rect 21376 66226 21496 66254
rect 21272 65204 21324 65210
rect 21272 65146 21324 65152
rect 21180 64660 21232 64666
rect 21180 64602 21232 64608
rect 20811 64220 21119 64240
rect 20811 64218 20817 64220
rect 20873 64218 20897 64220
rect 20953 64218 20977 64220
rect 21033 64218 21057 64220
rect 21113 64218 21119 64220
rect 20873 64166 20875 64218
rect 21055 64166 21057 64218
rect 20811 64164 20817 64166
rect 20873 64164 20897 64166
rect 20953 64164 20977 64166
rect 21033 64164 21057 64166
rect 21113 64164 21119 64166
rect 20811 64144 21119 64164
rect 20720 64048 20772 64054
rect 20720 63990 20772 63996
rect 20536 63980 20588 63986
rect 20536 63922 20588 63928
rect 20456 63838 20576 63866
rect 20352 63504 20404 63510
rect 20352 63446 20404 63452
rect 20260 63436 20312 63442
rect 20260 63378 20312 63384
rect 20364 62898 20392 63446
rect 19432 62892 19484 62898
rect 19432 62834 19484 62840
rect 20352 62892 20404 62898
rect 20352 62834 20404 62840
rect 19260 60608 19380 60636
rect 18970 60072 19026 60081
rect 18970 60007 18972 60016
rect 19024 60007 19026 60016
rect 18972 59978 19024 59984
rect 19156 59968 19208 59974
rect 19156 59910 19208 59916
rect 19168 59702 19196 59910
rect 19156 59696 19208 59702
rect 19156 59638 19208 59644
rect 19064 59628 19116 59634
rect 19064 59570 19116 59576
rect 18880 59492 18932 59498
rect 18880 59434 18932 59440
rect 18892 55418 18920 59434
rect 19076 58698 19104 59570
rect 19076 58682 19196 58698
rect 19076 58676 19208 58682
rect 19076 58670 19156 58676
rect 19156 58618 19208 58624
rect 19260 58614 19288 60608
rect 19338 60208 19394 60217
rect 19338 60143 19340 60152
rect 19392 60143 19394 60152
rect 19340 60114 19392 60120
rect 19248 58608 19300 58614
rect 19248 58550 19300 58556
rect 19340 57452 19392 57458
rect 19340 57394 19392 57400
rect 19248 56840 19300 56846
rect 19248 56782 19300 56788
rect 19064 56364 19116 56370
rect 19064 56306 19116 56312
rect 18880 55412 18932 55418
rect 18880 55354 18932 55360
rect 18788 55072 18840 55078
rect 18788 55014 18840 55020
rect 18696 53780 18748 53786
rect 18696 53722 18748 53728
rect 18236 53168 18288 53174
rect 18236 53110 18288 53116
rect 18328 53100 18380 53106
rect 18328 53042 18380 53048
rect 18340 52698 18368 53042
rect 17868 52692 17920 52698
rect 17868 52634 17920 52640
rect 18328 52692 18380 52698
rect 18328 52634 18380 52640
rect 18512 52624 18564 52630
rect 18512 52566 18564 52572
rect 18052 52488 18104 52494
rect 18052 52430 18104 52436
rect 18328 52488 18380 52494
rect 18328 52430 18380 52436
rect 17776 52420 17828 52426
rect 17776 52362 17828 52368
rect 18064 52086 18092 52430
rect 18052 52080 18104 52086
rect 18052 52022 18104 52028
rect 17960 52012 18012 52018
rect 17960 51954 18012 51960
rect 17972 51610 18000 51954
rect 18340 51950 18368 52430
rect 18328 51944 18380 51950
rect 18328 51886 18380 51892
rect 17960 51604 18012 51610
rect 17960 51546 18012 51552
rect 18340 51474 18368 51886
rect 18328 51468 18380 51474
rect 18328 51410 18380 51416
rect 17684 51400 17736 51406
rect 17684 51342 17736 51348
rect 17328 51046 17540 51074
rect 17328 50930 17356 51046
rect 17316 50924 17368 50930
rect 17316 50866 17368 50872
rect 17132 49768 17184 49774
rect 17132 49710 17184 49716
rect 17040 47184 17092 47190
rect 17040 47126 17092 47132
rect 16948 45824 17000 45830
rect 16948 45766 17000 45772
rect 16960 45558 16988 45766
rect 16948 45552 17000 45558
rect 16948 45494 17000 45500
rect 16948 45076 17000 45082
rect 16948 45018 17000 45024
rect 16776 44118 16896 44146
rect 16580 43988 16632 43994
rect 16580 43930 16632 43936
rect 16672 42220 16724 42226
rect 16672 42162 16724 42168
rect 16684 42022 16712 42162
rect 16672 42016 16724 42022
rect 16672 41958 16724 41964
rect 16684 41138 16712 41958
rect 16672 41132 16724 41138
rect 16672 41074 16724 41080
rect 16580 39840 16632 39846
rect 16580 39782 16632 39788
rect 16592 39506 16620 39782
rect 16580 39500 16632 39506
rect 16580 39442 16632 39448
rect 16592 39030 16620 39442
rect 16580 39024 16632 39030
rect 16580 38966 16632 38972
rect 16488 38480 16540 38486
rect 16488 38422 16540 38428
rect 16672 38276 16724 38282
rect 16672 38218 16724 38224
rect 16684 38010 16712 38218
rect 16672 38004 16724 38010
rect 16672 37946 16724 37952
rect 16672 37256 16724 37262
rect 16672 37198 16724 37204
rect 16488 37120 16540 37126
rect 16488 37062 16540 37068
rect 16500 36922 16528 37062
rect 16488 36916 16540 36922
rect 16488 36858 16540 36864
rect 16580 36848 16632 36854
rect 16580 36790 16632 36796
rect 16304 36712 16356 36718
rect 15842 36680 15898 36689
rect 16304 36654 16356 36660
rect 15842 36615 15898 36624
rect 16592 36582 16620 36790
rect 16580 36576 16632 36582
rect 16580 36518 16632 36524
rect 15846 36476 16154 36496
rect 15846 36474 15852 36476
rect 15908 36474 15932 36476
rect 15988 36474 16012 36476
rect 16068 36474 16092 36476
rect 16148 36474 16154 36476
rect 15908 36422 15910 36474
rect 16090 36422 16092 36474
rect 15846 36420 15852 36422
rect 15908 36420 15932 36422
rect 15988 36420 16012 36422
rect 16068 36420 16092 36422
rect 16148 36420 16154 36422
rect 15846 36400 16154 36420
rect 15752 36372 15804 36378
rect 15752 36314 15804 36320
rect 15764 34678 15792 36314
rect 16684 35766 16712 37198
rect 16672 35760 16724 35766
rect 16672 35702 16724 35708
rect 15846 35388 16154 35408
rect 15846 35386 15852 35388
rect 15908 35386 15932 35388
rect 15988 35386 16012 35388
rect 16068 35386 16092 35388
rect 16148 35386 16154 35388
rect 15908 35334 15910 35386
rect 16090 35334 16092 35386
rect 15846 35332 15852 35334
rect 15908 35332 15932 35334
rect 15988 35332 16012 35334
rect 16068 35332 16092 35334
rect 16148 35332 16154 35334
rect 15846 35312 16154 35332
rect 16396 35216 16448 35222
rect 16396 35158 16448 35164
rect 15752 34672 15804 34678
rect 15752 34614 15804 34620
rect 15846 34300 16154 34320
rect 15846 34298 15852 34300
rect 15908 34298 15932 34300
rect 15988 34298 16012 34300
rect 16068 34298 16092 34300
rect 16148 34298 16154 34300
rect 15908 34246 15910 34298
rect 16090 34246 16092 34298
rect 15846 34244 15852 34246
rect 15908 34244 15932 34246
rect 15988 34244 16012 34246
rect 16068 34244 16092 34246
rect 16148 34244 16154 34246
rect 15846 34224 16154 34244
rect 16212 33516 16264 33522
rect 16212 33458 16264 33464
rect 15846 33212 16154 33232
rect 15846 33210 15852 33212
rect 15908 33210 15932 33212
rect 15988 33210 16012 33212
rect 16068 33210 16092 33212
rect 16148 33210 16154 33212
rect 15908 33158 15910 33210
rect 16090 33158 16092 33210
rect 15846 33156 15852 33158
rect 15908 33156 15932 33158
rect 15988 33156 16012 33158
rect 16068 33156 16092 33158
rect 16148 33156 16154 33158
rect 15846 33136 16154 33156
rect 16224 33114 16252 33458
rect 16212 33108 16264 33114
rect 16212 33050 16264 33056
rect 15752 32224 15804 32230
rect 15752 32166 15804 32172
rect 16304 32224 16356 32230
rect 16304 32166 16356 32172
rect 15580 31726 15700 31754
rect 15580 31686 15608 31726
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15660 31680 15712 31686
rect 15660 31622 15712 31628
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 15580 30734 15608 31350
rect 15672 31346 15700 31622
rect 15660 31340 15712 31346
rect 15660 31282 15712 31288
rect 15660 31136 15712 31142
rect 15660 31078 15712 31084
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15476 30592 15528 30598
rect 15476 30534 15528 30540
rect 15488 29594 15516 30534
rect 15488 29566 15608 29594
rect 15304 28966 15424 28994
rect 15396 28422 15424 28966
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15304 27402 15332 28358
rect 15396 27674 15424 28358
rect 15488 27946 15516 28494
rect 15476 27940 15528 27946
rect 15476 27882 15528 27888
rect 15474 27840 15530 27849
rect 15474 27775 15530 27784
rect 15384 27668 15436 27674
rect 15384 27610 15436 27616
rect 15382 27568 15438 27577
rect 15382 27503 15438 27512
rect 15292 27396 15344 27402
rect 15292 27338 15344 27344
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15396 24682 15424 27503
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 10880 20700 11188 20720
rect 10880 20698 10886 20700
rect 10942 20698 10966 20700
rect 11022 20698 11046 20700
rect 11102 20698 11126 20700
rect 11182 20698 11188 20700
rect 10942 20646 10944 20698
rect 11124 20646 11126 20698
rect 10880 20644 10886 20646
rect 10942 20644 10966 20646
rect 11022 20644 11046 20646
rect 11102 20644 11126 20646
rect 11182 20644 11188 20646
rect 10880 20624 11188 20644
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 10880 19612 11188 19632
rect 10880 19610 10886 19612
rect 10942 19610 10966 19612
rect 11022 19610 11046 19612
rect 11102 19610 11126 19612
rect 11182 19610 11188 19612
rect 10942 19558 10944 19610
rect 11124 19558 11126 19610
rect 10880 19556 10886 19558
rect 10942 19556 10966 19558
rect 11022 19556 11046 19558
rect 11102 19556 11126 19558
rect 11182 19556 11188 19558
rect 10880 19536 11188 19556
rect 10880 18524 11188 18544
rect 10880 18522 10886 18524
rect 10942 18522 10966 18524
rect 11022 18522 11046 18524
rect 11102 18522 11126 18524
rect 11182 18522 11188 18524
rect 10942 18470 10944 18522
rect 11124 18470 11126 18522
rect 10880 18468 10886 18470
rect 10942 18468 10966 18470
rect 11022 18468 11046 18470
rect 11102 18468 11126 18470
rect 11182 18468 11188 18470
rect 10880 18448 11188 18468
rect 10880 17436 11188 17456
rect 10880 17434 10886 17436
rect 10942 17434 10966 17436
rect 11022 17434 11046 17436
rect 11102 17434 11126 17436
rect 11182 17434 11188 17436
rect 10942 17382 10944 17434
rect 11124 17382 11126 17434
rect 10880 17380 10886 17382
rect 10942 17380 10966 17382
rect 11022 17380 11046 17382
rect 11102 17380 11126 17382
rect 11182 17380 11188 17382
rect 10880 17360 11188 17380
rect 10880 16348 11188 16368
rect 10880 16346 10886 16348
rect 10942 16346 10966 16348
rect 11022 16346 11046 16348
rect 11102 16346 11126 16348
rect 11182 16346 11188 16348
rect 10942 16294 10944 16346
rect 11124 16294 11126 16346
rect 10880 16292 10886 16294
rect 10942 16292 10966 16294
rect 11022 16292 11046 16294
rect 11102 16292 11126 16294
rect 11182 16292 11188 16294
rect 10880 16272 11188 16292
rect 10880 15260 11188 15280
rect 10880 15258 10886 15260
rect 10942 15258 10966 15260
rect 11022 15258 11046 15260
rect 11102 15258 11126 15260
rect 11182 15258 11188 15260
rect 10942 15206 10944 15258
rect 11124 15206 11126 15258
rect 10880 15204 10886 15206
rect 10942 15204 10966 15206
rect 11022 15204 11046 15206
rect 11102 15204 11126 15206
rect 11182 15204 11188 15206
rect 10880 15184 11188 15204
rect 10880 14172 11188 14192
rect 10880 14170 10886 14172
rect 10942 14170 10966 14172
rect 11022 14170 11046 14172
rect 11102 14170 11126 14172
rect 11182 14170 11188 14172
rect 10942 14118 10944 14170
rect 11124 14118 11126 14170
rect 10880 14116 10886 14118
rect 10942 14116 10966 14118
rect 11022 14116 11046 14118
rect 11102 14116 11126 14118
rect 11182 14116 11188 14118
rect 10880 14096 11188 14116
rect 10880 13084 11188 13104
rect 10880 13082 10886 13084
rect 10942 13082 10966 13084
rect 11022 13082 11046 13084
rect 11102 13082 11126 13084
rect 11182 13082 11188 13084
rect 10942 13030 10944 13082
rect 11124 13030 11126 13082
rect 10880 13028 10886 13030
rect 10942 13028 10966 13030
rect 11022 13028 11046 13030
rect 11102 13028 11126 13030
rect 11182 13028 11188 13030
rect 10880 13008 11188 13028
rect 10880 11996 11188 12016
rect 10880 11994 10886 11996
rect 10942 11994 10966 11996
rect 11022 11994 11046 11996
rect 11102 11994 11126 11996
rect 11182 11994 11188 11996
rect 10942 11942 10944 11994
rect 11124 11942 11126 11994
rect 10880 11940 10886 11942
rect 10942 11940 10966 11942
rect 11022 11940 11046 11942
rect 11102 11940 11126 11942
rect 11182 11940 11188 11942
rect 10880 11920 11188 11940
rect 10880 10908 11188 10928
rect 10880 10906 10886 10908
rect 10942 10906 10966 10908
rect 11022 10906 11046 10908
rect 11102 10906 11126 10908
rect 11182 10906 11188 10908
rect 10942 10854 10944 10906
rect 11124 10854 11126 10906
rect 10880 10852 10886 10854
rect 10942 10852 10966 10854
rect 11022 10852 11046 10854
rect 11102 10852 11126 10854
rect 11182 10852 11188 10854
rect 10880 10832 11188 10852
rect 10880 9820 11188 9840
rect 10880 9818 10886 9820
rect 10942 9818 10966 9820
rect 11022 9818 11046 9820
rect 11102 9818 11126 9820
rect 11182 9818 11188 9820
rect 10942 9766 10944 9818
rect 11124 9766 11126 9818
rect 10880 9764 10886 9766
rect 10942 9764 10966 9766
rect 11022 9764 11046 9766
rect 11102 9764 11126 9766
rect 11182 9764 11188 9766
rect 10880 9744 11188 9764
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 10880 8732 11188 8752
rect 10880 8730 10886 8732
rect 10942 8730 10966 8732
rect 11022 8730 11046 8732
rect 11102 8730 11126 8732
rect 11182 8730 11188 8732
rect 10942 8678 10944 8730
rect 11124 8678 11126 8730
rect 10880 8676 10886 8678
rect 10942 8676 10966 8678
rect 11022 8676 11046 8678
rect 11102 8676 11126 8678
rect 11182 8676 11188 8678
rect 10880 8656 11188 8676
rect 14292 8362 14320 23802
rect 15488 23254 15516 27775
rect 15580 26586 15608 29566
rect 15672 28082 15700 31078
rect 15764 29646 15792 32166
rect 15846 32124 16154 32144
rect 15846 32122 15852 32124
rect 15908 32122 15932 32124
rect 15988 32122 16012 32124
rect 16068 32122 16092 32124
rect 16148 32122 16154 32124
rect 15908 32070 15910 32122
rect 16090 32070 16092 32122
rect 15846 32068 15852 32070
rect 15908 32068 15932 32070
rect 15988 32068 16012 32070
rect 16068 32068 16092 32070
rect 16148 32068 16154 32070
rect 15846 32048 16154 32068
rect 15936 31952 15988 31958
rect 15936 31894 15988 31900
rect 15948 31346 15976 31894
rect 15936 31340 15988 31346
rect 15988 31300 16252 31328
rect 15936 31282 15988 31288
rect 15846 31036 16154 31056
rect 15846 31034 15852 31036
rect 15908 31034 15932 31036
rect 15988 31034 16012 31036
rect 16068 31034 16092 31036
rect 16148 31034 16154 31036
rect 15908 30982 15910 31034
rect 16090 30982 16092 31034
rect 15846 30980 15852 30982
rect 15908 30980 15932 30982
rect 15988 30980 16012 30982
rect 16068 30980 16092 30982
rect 16148 30980 16154 30982
rect 15846 30960 16154 30980
rect 16224 30666 16252 31300
rect 16212 30660 16264 30666
rect 16212 30602 16264 30608
rect 15846 29948 16154 29968
rect 15846 29946 15852 29948
rect 15908 29946 15932 29948
rect 15988 29946 16012 29948
rect 16068 29946 16092 29948
rect 16148 29946 16154 29948
rect 15908 29894 15910 29946
rect 16090 29894 16092 29946
rect 15846 29892 15852 29894
rect 15908 29892 15932 29894
rect 15988 29892 16012 29894
rect 16068 29892 16092 29894
rect 16148 29892 16154 29894
rect 15846 29872 16154 29892
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15764 28121 15792 29106
rect 15846 28860 16154 28880
rect 15846 28858 15852 28860
rect 15908 28858 15932 28860
rect 15988 28858 16012 28860
rect 16068 28858 16092 28860
rect 16148 28858 16154 28860
rect 15908 28806 15910 28858
rect 16090 28806 16092 28858
rect 15846 28804 15852 28806
rect 15908 28804 15932 28806
rect 15988 28804 16012 28806
rect 16068 28804 16092 28806
rect 16148 28804 16154 28806
rect 15846 28784 16154 28804
rect 15842 28248 15898 28257
rect 15842 28183 15844 28192
rect 15896 28183 15898 28192
rect 15844 28154 15896 28160
rect 15750 28112 15806 28121
rect 15660 28076 15712 28082
rect 15750 28047 15806 28056
rect 15660 28018 15712 28024
rect 15672 26874 15700 28018
rect 15752 28008 15804 28014
rect 15752 27950 15804 27956
rect 15764 27402 15792 27950
rect 15846 27772 16154 27792
rect 15846 27770 15852 27772
rect 15908 27770 15932 27772
rect 15988 27770 16012 27772
rect 16068 27770 16092 27772
rect 16148 27770 16154 27772
rect 15908 27718 15910 27770
rect 16090 27718 16092 27770
rect 15846 27716 15852 27718
rect 15908 27716 15932 27718
rect 15988 27716 16012 27718
rect 16068 27716 16092 27718
rect 16148 27716 16154 27718
rect 15846 27696 16154 27716
rect 15752 27396 15804 27402
rect 15752 27338 15804 27344
rect 15764 27062 15792 27338
rect 15752 27056 15804 27062
rect 16224 27033 16252 30602
rect 15752 26998 15804 27004
rect 16210 27024 16266 27033
rect 16210 26959 16266 26968
rect 15752 26920 15804 26926
rect 15672 26868 15752 26874
rect 16316 26874 16344 32166
rect 15672 26862 15804 26868
rect 15672 26846 15792 26862
rect 16224 26846 16344 26874
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15568 26580 15620 26586
rect 15568 26522 15620 26528
rect 15672 26450 15700 26726
rect 15846 26684 16154 26704
rect 15846 26682 15852 26684
rect 15908 26682 15932 26684
rect 15988 26682 16012 26684
rect 16068 26682 16092 26684
rect 16148 26682 16154 26684
rect 15908 26630 15910 26682
rect 16090 26630 16092 26682
rect 15846 26628 15852 26630
rect 15908 26628 15932 26630
rect 15988 26628 16012 26630
rect 16068 26628 16092 26630
rect 16148 26628 16154 26630
rect 15846 26608 16154 26628
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15846 25596 16154 25616
rect 15846 25594 15852 25596
rect 15908 25594 15932 25596
rect 15988 25594 16012 25596
rect 16068 25594 16092 25596
rect 16148 25594 16154 25596
rect 15908 25542 15910 25594
rect 16090 25542 16092 25594
rect 15846 25540 15852 25542
rect 15908 25540 15932 25542
rect 15988 25540 16012 25542
rect 16068 25540 16092 25542
rect 16148 25540 16154 25542
rect 15846 25520 16154 25540
rect 15846 24508 16154 24528
rect 15846 24506 15852 24508
rect 15908 24506 15932 24508
rect 15988 24506 16012 24508
rect 16068 24506 16092 24508
rect 16148 24506 16154 24508
rect 15908 24454 15910 24506
rect 16090 24454 16092 24506
rect 15846 24452 15852 24454
rect 15908 24452 15932 24454
rect 15988 24452 16012 24454
rect 16068 24452 16092 24454
rect 16148 24452 16154 24454
rect 15846 24432 16154 24452
rect 15846 23420 16154 23440
rect 15846 23418 15852 23420
rect 15908 23418 15932 23420
rect 15988 23418 16012 23420
rect 16068 23418 16092 23420
rect 16148 23418 16154 23420
rect 15908 23366 15910 23418
rect 16090 23366 16092 23418
rect 15846 23364 15852 23366
rect 15908 23364 15932 23366
rect 15988 23364 16012 23366
rect 16068 23364 16092 23366
rect 16148 23364 16154 23366
rect 15846 23344 16154 23364
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15846 22332 16154 22352
rect 15846 22330 15852 22332
rect 15908 22330 15932 22332
rect 15988 22330 16012 22332
rect 16068 22330 16092 22332
rect 16148 22330 16154 22332
rect 15908 22278 15910 22330
rect 16090 22278 16092 22330
rect 15846 22276 15852 22278
rect 15908 22276 15932 22278
rect 15988 22276 16012 22278
rect 16068 22276 16092 22278
rect 16148 22276 16154 22278
rect 15846 22256 16154 22276
rect 15846 21244 16154 21264
rect 15846 21242 15852 21244
rect 15908 21242 15932 21244
rect 15988 21242 16012 21244
rect 16068 21242 16092 21244
rect 16148 21242 16154 21244
rect 15908 21190 15910 21242
rect 16090 21190 16092 21242
rect 15846 21188 15852 21190
rect 15908 21188 15932 21190
rect 15988 21188 16012 21190
rect 16068 21188 16092 21190
rect 16148 21188 16154 21190
rect 15846 21168 16154 21188
rect 15846 20156 16154 20176
rect 15846 20154 15852 20156
rect 15908 20154 15932 20156
rect 15988 20154 16012 20156
rect 16068 20154 16092 20156
rect 16148 20154 16154 20156
rect 15908 20102 15910 20154
rect 16090 20102 16092 20154
rect 15846 20100 15852 20102
rect 15908 20100 15932 20102
rect 15988 20100 16012 20102
rect 16068 20100 16092 20102
rect 16148 20100 16154 20102
rect 15846 20080 16154 20100
rect 15846 19068 16154 19088
rect 15846 19066 15852 19068
rect 15908 19066 15932 19068
rect 15988 19066 16012 19068
rect 16068 19066 16092 19068
rect 16148 19066 16154 19068
rect 15908 19014 15910 19066
rect 16090 19014 16092 19066
rect 15846 19012 15852 19014
rect 15908 19012 15932 19014
rect 15988 19012 16012 19014
rect 16068 19012 16092 19014
rect 16148 19012 16154 19014
rect 15846 18992 16154 19012
rect 15846 17980 16154 18000
rect 15846 17978 15852 17980
rect 15908 17978 15932 17980
rect 15988 17978 16012 17980
rect 16068 17978 16092 17980
rect 16148 17978 16154 17980
rect 15908 17926 15910 17978
rect 16090 17926 16092 17978
rect 15846 17924 15852 17926
rect 15908 17924 15932 17926
rect 15988 17924 16012 17926
rect 16068 17924 16092 17926
rect 16148 17924 16154 17926
rect 15846 17904 16154 17924
rect 15846 16892 16154 16912
rect 15846 16890 15852 16892
rect 15908 16890 15932 16892
rect 15988 16890 16012 16892
rect 16068 16890 16092 16892
rect 16148 16890 16154 16892
rect 15908 16838 15910 16890
rect 16090 16838 16092 16890
rect 15846 16836 15852 16838
rect 15908 16836 15932 16838
rect 15988 16836 16012 16838
rect 16068 16836 16092 16838
rect 16148 16836 16154 16838
rect 15846 16816 16154 16836
rect 16224 16590 16252 26846
rect 16302 26752 16358 26761
rect 16302 26687 16358 26696
rect 16316 19836 16344 26687
rect 16408 25294 16436 35158
rect 16580 33040 16632 33046
rect 16580 32982 16632 32988
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16500 28150 16528 28426
rect 16488 28144 16540 28150
rect 16488 28086 16540 28092
rect 16500 27334 16528 28086
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16500 27130 16528 27270
rect 16488 27124 16540 27130
rect 16488 27066 16540 27072
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16592 25242 16620 32982
rect 16684 31822 16712 35702
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16684 31278 16712 31758
rect 16776 31754 16804 44118
rect 16960 42294 16988 45018
rect 17144 44878 17172 49710
rect 17328 47954 17356 50866
rect 17592 48612 17644 48618
rect 17592 48554 17644 48560
rect 17408 48544 17460 48550
rect 17408 48486 17460 48492
rect 17420 48074 17448 48486
rect 17408 48068 17460 48074
rect 17408 48010 17460 48016
rect 17328 47926 17448 47954
rect 17236 47666 17356 47682
rect 17236 47660 17368 47666
rect 17236 47654 17316 47660
rect 17236 46986 17264 47654
rect 17316 47602 17368 47608
rect 17314 47152 17370 47161
rect 17314 47087 17316 47096
rect 17368 47087 17370 47096
rect 17316 47058 17368 47064
rect 17224 46980 17276 46986
rect 17224 46922 17276 46928
rect 17420 45830 17448 47926
rect 17480 47660 17532 47666
rect 17532 47608 17540 47648
rect 17480 47602 17540 47608
rect 17512 47258 17540 47602
rect 17604 47530 17632 48554
rect 17696 47802 17724 51342
rect 17776 49360 17828 49366
rect 17776 49302 17828 49308
rect 17788 48754 17816 49302
rect 18524 48822 18552 52566
rect 18512 48816 18564 48822
rect 18512 48758 18564 48764
rect 17776 48748 17828 48754
rect 17776 48690 17828 48696
rect 17776 48612 17828 48618
rect 17776 48554 17828 48560
rect 17684 47796 17736 47802
rect 17684 47738 17736 47744
rect 17788 47682 17816 48554
rect 18524 48346 18552 48758
rect 18512 48340 18564 48346
rect 18512 48282 18564 48288
rect 18972 48340 19024 48346
rect 18972 48282 19024 48288
rect 18512 48136 18564 48142
rect 18512 48078 18564 48084
rect 18420 48000 18472 48006
rect 18420 47942 18472 47948
rect 17866 47832 17922 47841
rect 17866 47767 17868 47776
rect 17920 47767 17922 47776
rect 17868 47738 17920 47744
rect 17696 47654 17816 47682
rect 18328 47660 18380 47666
rect 17696 47530 17724 47654
rect 18328 47602 18380 47608
rect 17960 47592 18012 47598
rect 17788 47540 17960 47546
rect 17788 47534 18012 47540
rect 17592 47524 17644 47530
rect 17592 47466 17644 47472
rect 17684 47524 17736 47530
rect 17684 47466 17736 47472
rect 17788 47518 18000 47534
rect 17500 47252 17552 47258
rect 17500 47194 17552 47200
rect 17408 45824 17460 45830
rect 17408 45766 17460 45772
rect 17132 44872 17184 44878
rect 17132 44814 17184 44820
rect 17224 44464 17276 44470
rect 17224 44406 17276 44412
rect 17132 44328 17184 44334
rect 17132 44270 17184 44276
rect 17144 43858 17172 44270
rect 17132 43852 17184 43858
rect 17132 43794 17184 43800
rect 17040 43308 17092 43314
rect 17040 43250 17092 43256
rect 17052 42362 17080 43250
rect 17144 42770 17172 43794
rect 17132 42764 17184 42770
rect 17132 42706 17184 42712
rect 17040 42356 17092 42362
rect 17040 42298 17092 42304
rect 16948 42288 17000 42294
rect 16948 42230 17000 42236
rect 16856 42152 16908 42158
rect 16856 42094 16908 42100
rect 16868 41414 16896 42094
rect 17132 42084 17184 42090
rect 17132 42026 17184 42032
rect 16868 41386 16988 41414
rect 16960 40662 16988 41386
rect 17040 40928 17092 40934
rect 17040 40870 17092 40876
rect 16948 40656 17000 40662
rect 16948 40598 17000 40604
rect 16948 40520 17000 40526
rect 16948 40462 17000 40468
rect 16856 40384 16908 40390
rect 16856 40326 16908 40332
rect 16868 36174 16896 40326
rect 16960 39642 16988 40462
rect 17052 40118 17080 40870
rect 17040 40112 17092 40118
rect 17040 40054 17092 40060
rect 16948 39636 17000 39642
rect 16948 39578 17000 39584
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16948 34944 17000 34950
rect 16948 34886 17000 34892
rect 16960 33590 16988 34886
rect 16948 33584 17000 33590
rect 16948 33526 17000 33532
rect 17144 32910 17172 42026
rect 17236 41818 17264 44406
rect 17604 44334 17632 47466
rect 17696 44470 17724 47466
rect 17788 44538 17816 47518
rect 18144 47048 18196 47054
rect 18144 46990 18196 46996
rect 17960 46572 18012 46578
rect 17960 46514 18012 46520
rect 17972 46102 18000 46514
rect 17960 46096 18012 46102
rect 17960 46038 18012 46044
rect 17868 44804 17920 44810
rect 17868 44746 17920 44752
rect 17776 44532 17828 44538
rect 17776 44474 17828 44480
rect 17684 44464 17736 44470
rect 17684 44406 17736 44412
rect 17592 44328 17644 44334
rect 17592 44270 17644 44276
rect 17408 42152 17460 42158
rect 17408 42094 17460 42100
rect 17224 41812 17276 41818
rect 17224 41754 17276 41760
rect 17420 40730 17448 42094
rect 17604 41274 17632 44270
rect 17684 44192 17736 44198
rect 17684 44134 17736 44140
rect 17696 42226 17724 44134
rect 17776 43988 17828 43994
rect 17776 43930 17828 43936
rect 17684 42220 17736 42226
rect 17684 42162 17736 42168
rect 17788 41682 17816 43930
rect 17776 41676 17828 41682
rect 17776 41618 17828 41624
rect 17592 41268 17644 41274
rect 17644 41228 17724 41256
rect 17592 41210 17644 41216
rect 17500 41132 17552 41138
rect 17500 41074 17552 41080
rect 17512 41002 17540 41074
rect 17500 40996 17552 41002
rect 17500 40938 17552 40944
rect 17592 40928 17644 40934
rect 17592 40870 17644 40876
rect 17408 40724 17460 40730
rect 17408 40666 17460 40672
rect 17316 40656 17368 40662
rect 17316 40598 17368 40604
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 17236 39098 17264 39238
rect 17224 39092 17276 39098
rect 17224 39034 17276 39040
rect 17328 38298 17356 40598
rect 17604 39438 17632 40870
rect 17592 39432 17644 39438
rect 17592 39374 17644 39380
rect 17408 39364 17460 39370
rect 17408 39306 17460 39312
rect 17420 38894 17448 39306
rect 17408 38888 17460 38894
rect 17408 38830 17460 38836
rect 17420 38758 17448 38830
rect 17408 38752 17460 38758
rect 17408 38694 17460 38700
rect 17236 38270 17356 38298
rect 17236 37806 17264 38270
rect 17316 37868 17368 37874
rect 17316 37810 17368 37816
rect 17224 37800 17276 37806
rect 17224 37742 17276 37748
rect 17236 37466 17264 37742
rect 17224 37460 17276 37466
rect 17224 37402 17276 37408
rect 17236 36786 17264 37402
rect 17224 36780 17276 36786
rect 17224 36722 17276 36728
rect 17328 36650 17356 37810
rect 17316 36644 17368 36650
rect 17316 36586 17368 36592
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17328 34542 17356 35090
rect 17420 35018 17448 38694
rect 17696 38554 17724 41228
rect 17880 40730 17908 44746
rect 18052 44396 18104 44402
rect 18052 44338 18104 44344
rect 18064 44198 18092 44338
rect 18052 44192 18104 44198
rect 18052 44134 18104 44140
rect 18156 43450 18184 46990
rect 18340 46442 18368 47602
rect 18328 46436 18380 46442
rect 18328 46378 18380 46384
rect 18236 45892 18288 45898
rect 18236 45834 18288 45840
rect 18144 43444 18196 43450
rect 18144 43386 18196 43392
rect 18156 42650 18184 43386
rect 17972 42622 18184 42650
rect 17972 41614 18000 42622
rect 18248 42566 18276 45834
rect 18432 45558 18460 47942
rect 18524 47802 18552 48078
rect 18512 47796 18564 47802
rect 18512 47738 18564 47744
rect 18880 46572 18932 46578
rect 18880 46514 18932 46520
rect 18892 46034 18920 46514
rect 18880 46028 18932 46034
rect 18880 45970 18932 45976
rect 18420 45552 18472 45558
rect 18420 45494 18472 45500
rect 18328 44396 18380 44402
rect 18328 44338 18380 44344
rect 18236 42560 18288 42566
rect 18236 42502 18288 42508
rect 17960 41608 18012 41614
rect 17960 41550 18012 41556
rect 18236 41540 18288 41546
rect 18236 41482 18288 41488
rect 18144 41472 18196 41478
rect 18144 41414 18196 41420
rect 17868 40724 17920 40730
rect 17868 40666 17920 40672
rect 18052 40520 18104 40526
rect 18052 40462 18104 40468
rect 17960 40384 18012 40390
rect 17960 40326 18012 40332
rect 17868 39296 17920 39302
rect 17868 39238 17920 39244
rect 17880 39030 17908 39238
rect 17868 39024 17920 39030
rect 17868 38966 17920 38972
rect 17684 38548 17736 38554
rect 17684 38490 17736 38496
rect 17696 37398 17724 38490
rect 17972 38350 18000 40326
rect 18064 38554 18092 40462
rect 18052 38548 18104 38554
rect 18052 38490 18104 38496
rect 17960 38344 18012 38350
rect 17960 38286 18012 38292
rect 17684 37392 17736 37398
rect 17684 37334 17736 37340
rect 18156 35170 18184 41414
rect 18248 39914 18276 41482
rect 18340 41206 18368 44338
rect 18432 42702 18460 45494
rect 18512 45484 18564 45490
rect 18512 45426 18564 45432
rect 18420 42696 18472 42702
rect 18420 42638 18472 42644
rect 18524 42022 18552 45426
rect 18604 44396 18656 44402
rect 18604 44338 18656 44344
rect 18616 44305 18644 44338
rect 18602 44296 18658 44305
rect 18602 44231 18658 44240
rect 18788 44192 18840 44198
rect 18788 44134 18840 44140
rect 18604 42628 18656 42634
rect 18604 42570 18656 42576
rect 18512 42016 18564 42022
rect 18512 41958 18564 41964
rect 18524 41750 18552 41958
rect 18512 41744 18564 41750
rect 18512 41686 18564 41692
rect 18616 41274 18644 42570
rect 18800 42090 18828 44134
rect 18984 42566 19012 48282
rect 19076 46714 19104 56306
rect 19260 53242 19288 56782
rect 19352 56166 19380 57394
rect 19340 56160 19392 56166
rect 19340 56102 19392 56108
rect 19352 54262 19380 56102
rect 19340 54256 19392 54262
rect 19340 54198 19392 54204
rect 19444 53786 19472 62834
rect 19984 62688 20036 62694
rect 19984 62630 20036 62636
rect 19708 61872 19760 61878
rect 19708 61814 19760 61820
rect 19720 61198 19748 61814
rect 19708 61192 19760 61198
rect 19708 61134 19760 61140
rect 19708 61056 19760 61062
rect 19708 60998 19760 61004
rect 19720 60858 19748 60998
rect 19708 60852 19760 60858
rect 19708 60794 19760 60800
rect 19616 60716 19668 60722
rect 19616 60658 19668 60664
rect 19628 60518 19656 60658
rect 19616 60512 19668 60518
rect 19616 60454 19668 60460
rect 19616 60104 19668 60110
rect 19720 60092 19748 60794
rect 19800 60648 19852 60654
rect 19800 60590 19852 60596
rect 19812 60110 19840 60590
rect 19890 60208 19946 60217
rect 19890 60143 19946 60152
rect 19904 60110 19932 60143
rect 19668 60064 19748 60092
rect 19800 60104 19852 60110
rect 19616 60046 19668 60052
rect 19800 60046 19852 60052
rect 19892 60104 19944 60110
rect 19892 60046 19944 60052
rect 19524 58540 19576 58546
rect 19524 58482 19576 58488
rect 19432 53780 19484 53786
rect 19432 53722 19484 53728
rect 19340 53644 19392 53650
rect 19340 53586 19392 53592
rect 19248 53236 19300 53242
rect 19248 53178 19300 53184
rect 19156 53100 19208 53106
rect 19156 53042 19208 53048
rect 19168 51882 19196 53042
rect 19248 52964 19300 52970
rect 19248 52906 19300 52912
rect 19156 51876 19208 51882
rect 19156 51818 19208 51824
rect 19260 48142 19288 52906
rect 19352 51610 19380 53586
rect 19340 51604 19392 51610
rect 19340 51546 19392 51552
rect 19444 51074 19472 53722
rect 19536 51610 19564 58482
rect 19628 57458 19656 60046
rect 19812 57497 19840 60046
rect 19892 59628 19944 59634
rect 19892 59570 19944 59576
rect 19798 57488 19854 57497
rect 19616 57452 19668 57458
rect 19904 57458 19932 59570
rect 19668 57412 19748 57440
rect 19798 57423 19800 57432
rect 19616 57394 19668 57400
rect 19616 55684 19668 55690
rect 19616 55626 19668 55632
rect 19524 51604 19576 51610
rect 19524 51546 19576 51552
rect 19352 51046 19472 51074
rect 19248 48136 19300 48142
rect 19248 48078 19300 48084
rect 19156 47456 19208 47462
rect 19156 47398 19208 47404
rect 19168 47161 19196 47398
rect 19260 47190 19288 48078
rect 19248 47184 19300 47190
rect 19154 47152 19210 47161
rect 19248 47126 19300 47132
rect 19154 47087 19210 47096
rect 19352 47054 19380 51046
rect 19432 50992 19484 50998
rect 19432 50934 19484 50940
rect 19444 48210 19472 50934
rect 19524 49836 19576 49842
rect 19524 49778 19576 49784
rect 19536 48618 19564 49778
rect 19524 48612 19576 48618
rect 19524 48554 19576 48560
rect 19524 48272 19576 48278
rect 19524 48214 19576 48220
rect 19432 48204 19484 48210
rect 19432 48146 19484 48152
rect 19432 48000 19484 48006
rect 19432 47942 19484 47948
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 19064 46708 19116 46714
rect 19064 46650 19116 46656
rect 19444 46646 19472 47942
rect 19432 46640 19484 46646
rect 19432 46582 19484 46588
rect 19536 45506 19564 48214
rect 19628 47546 19656 55626
rect 19720 55214 19748 57412
rect 19852 57423 19854 57432
rect 19892 57452 19944 57458
rect 19800 57394 19852 57400
rect 19892 57394 19944 57400
rect 19812 56778 19840 57394
rect 19800 56772 19852 56778
rect 19800 56714 19852 56720
rect 19800 55276 19852 55282
rect 19800 55218 19852 55224
rect 19708 55208 19760 55214
rect 19708 55150 19760 55156
rect 19812 55162 19840 55218
rect 19812 55134 19932 55162
rect 19800 55072 19852 55078
rect 19800 55014 19852 55020
rect 19812 54194 19840 55014
rect 19904 54330 19932 55134
rect 19892 54324 19944 54330
rect 19892 54266 19944 54272
rect 19800 54188 19852 54194
rect 19800 54130 19852 54136
rect 19708 54120 19760 54126
rect 19708 54062 19760 54068
rect 19720 53242 19748 54062
rect 19800 53644 19852 53650
rect 19800 53586 19852 53592
rect 19708 53236 19760 53242
rect 19708 53178 19760 53184
rect 19812 52902 19840 53586
rect 19996 53582 20024 62630
rect 20168 61328 20220 61334
rect 20168 61270 20220 61276
rect 20180 59106 20208 61270
rect 20260 61192 20312 61198
rect 20260 61134 20312 61140
rect 20272 59226 20300 61134
rect 20548 60178 20576 63838
rect 20732 63442 20760 63990
rect 20720 63436 20772 63442
rect 20720 63378 20772 63384
rect 21272 63232 21324 63238
rect 21272 63174 21324 63180
rect 20811 63132 21119 63152
rect 20811 63130 20817 63132
rect 20873 63130 20897 63132
rect 20953 63130 20977 63132
rect 21033 63130 21057 63132
rect 21113 63130 21119 63132
rect 20873 63078 20875 63130
rect 21055 63078 21057 63130
rect 20811 63076 20817 63078
rect 20873 63076 20897 63078
rect 20953 63076 20977 63078
rect 21033 63076 21057 63078
rect 21113 63076 21119 63078
rect 20811 63056 21119 63076
rect 21088 62688 21140 62694
rect 21088 62630 21140 62636
rect 21100 62354 21128 62630
rect 21088 62348 21140 62354
rect 21088 62290 21140 62296
rect 20811 62044 21119 62064
rect 20811 62042 20817 62044
rect 20873 62042 20897 62044
rect 20953 62042 20977 62044
rect 21033 62042 21057 62044
rect 21113 62042 21119 62044
rect 20873 61990 20875 62042
rect 21055 61990 21057 62042
rect 20811 61988 20817 61990
rect 20873 61988 20897 61990
rect 20953 61988 20977 61990
rect 21033 61988 21057 61990
rect 21113 61988 21119 61990
rect 20811 61968 21119 61988
rect 21180 61872 21232 61878
rect 21180 61814 21232 61820
rect 20811 60956 21119 60976
rect 20811 60954 20817 60956
rect 20873 60954 20897 60956
rect 20953 60954 20977 60956
rect 21033 60954 21057 60956
rect 21113 60954 21119 60956
rect 20873 60902 20875 60954
rect 21055 60902 21057 60954
rect 20811 60900 20817 60902
rect 20873 60900 20897 60902
rect 20953 60900 20977 60902
rect 21033 60900 21057 60902
rect 21113 60900 21119 60902
rect 20811 60880 21119 60900
rect 20810 60752 20866 60761
rect 21192 60722 21220 61814
rect 20810 60687 20812 60696
rect 20864 60687 20866 60696
rect 21180 60716 21232 60722
rect 20812 60658 20864 60664
rect 21180 60658 21232 60664
rect 20628 60512 20680 60518
rect 20628 60454 20680 60460
rect 20352 60172 20404 60178
rect 20352 60114 20404 60120
rect 20536 60172 20588 60178
rect 20536 60114 20588 60120
rect 20260 59220 20312 59226
rect 20260 59162 20312 59168
rect 20180 59078 20300 59106
rect 20168 58948 20220 58954
rect 20168 58890 20220 58896
rect 20076 58540 20128 58546
rect 20076 58482 20128 58488
rect 19984 53576 20036 53582
rect 19984 53518 20036 53524
rect 19800 52896 19852 52902
rect 19800 52838 19852 52844
rect 20088 52714 20116 58482
rect 20180 56166 20208 58890
rect 20272 57526 20300 59078
rect 20364 58546 20392 60114
rect 20640 60042 20668 60454
rect 20536 60036 20588 60042
rect 20536 59978 20588 59984
rect 20628 60036 20680 60042
rect 20628 59978 20680 59984
rect 20548 59498 20576 59978
rect 20811 59868 21119 59888
rect 20811 59866 20817 59868
rect 20873 59866 20897 59868
rect 20953 59866 20977 59868
rect 21033 59866 21057 59868
rect 21113 59866 21119 59868
rect 20873 59814 20875 59866
rect 21055 59814 21057 59866
rect 20811 59812 20817 59814
rect 20873 59812 20897 59814
rect 20953 59812 20977 59814
rect 21033 59812 21057 59814
rect 21113 59812 21119 59814
rect 20811 59792 21119 59812
rect 20536 59492 20588 59498
rect 20536 59434 20588 59440
rect 20536 59220 20588 59226
rect 20536 59162 20588 59168
rect 20548 59022 20576 59162
rect 20536 59016 20588 59022
rect 20536 58958 20588 58964
rect 20352 58540 20404 58546
rect 20352 58482 20404 58488
rect 20444 57792 20496 57798
rect 20444 57734 20496 57740
rect 20260 57520 20312 57526
rect 20260 57462 20312 57468
rect 20352 57248 20404 57254
rect 20352 57190 20404 57196
rect 20364 56846 20392 57190
rect 20352 56840 20404 56846
rect 20352 56782 20404 56788
rect 20456 56778 20484 57734
rect 20548 57594 20576 58958
rect 20811 58780 21119 58800
rect 20811 58778 20817 58780
rect 20873 58778 20897 58780
rect 20953 58778 20977 58780
rect 21033 58778 21057 58780
rect 21113 58778 21119 58780
rect 20873 58726 20875 58778
rect 21055 58726 21057 58778
rect 20811 58724 20817 58726
rect 20873 58724 20897 58726
rect 20953 58724 20977 58726
rect 21033 58724 21057 58726
rect 21113 58724 21119 58726
rect 20811 58704 21119 58724
rect 21192 58614 21220 60658
rect 21180 58608 21232 58614
rect 21180 58550 21232 58556
rect 21180 58472 21232 58478
rect 21180 58414 21232 58420
rect 20811 57692 21119 57712
rect 20811 57690 20817 57692
rect 20873 57690 20897 57692
rect 20953 57690 20977 57692
rect 21033 57690 21057 57692
rect 21113 57690 21119 57692
rect 20873 57638 20875 57690
rect 21055 57638 21057 57690
rect 20811 57636 20817 57638
rect 20873 57636 20897 57638
rect 20953 57636 20977 57638
rect 21033 57636 21057 57638
rect 21113 57636 21119 57638
rect 20811 57616 21119 57636
rect 20536 57588 20588 57594
rect 20536 57530 20588 57536
rect 20260 56772 20312 56778
rect 20260 56714 20312 56720
rect 20444 56772 20496 56778
rect 20444 56714 20496 56720
rect 20168 56160 20220 56166
rect 20168 56102 20220 56108
rect 20180 53174 20208 56102
rect 20272 55214 20300 56714
rect 20260 55208 20312 55214
rect 20260 55150 20312 55156
rect 20168 53168 20220 53174
rect 20168 53110 20220 53116
rect 19720 52686 20116 52714
rect 19720 51066 19748 52686
rect 19892 52420 19944 52426
rect 19892 52362 19944 52368
rect 19800 52352 19852 52358
rect 19800 52294 19852 52300
rect 19812 52154 19840 52294
rect 19800 52148 19852 52154
rect 19800 52090 19852 52096
rect 19812 51338 19840 52090
rect 19904 51474 19932 52362
rect 19892 51468 19944 51474
rect 19892 51410 19944 51416
rect 19800 51332 19852 51338
rect 19800 51274 19852 51280
rect 19812 51074 19840 51274
rect 19708 51060 19760 51066
rect 19812 51046 19932 51074
rect 19708 51002 19760 51008
rect 19708 50312 19760 50318
rect 19708 50254 19760 50260
rect 19720 49434 19748 50254
rect 19708 49428 19760 49434
rect 19708 49370 19760 49376
rect 19800 49292 19852 49298
rect 19800 49234 19852 49240
rect 19812 48822 19840 49234
rect 19800 48816 19852 48822
rect 19800 48758 19852 48764
rect 19800 48204 19852 48210
rect 19800 48146 19852 48152
rect 19628 47518 19748 47546
rect 19812 47530 19840 48146
rect 19616 47184 19668 47190
rect 19616 47126 19668 47132
rect 19260 45478 19564 45506
rect 19260 44334 19288 45478
rect 19524 45280 19576 45286
rect 19524 45222 19576 45228
rect 19432 45008 19484 45014
rect 19432 44950 19484 44956
rect 19340 44872 19392 44878
rect 19340 44814 19392 44820
rect 19248 44328 19300 44334
rect 19248 44270 19300 44276
rect 19156 43920 19208 43926
rect 19156 43862 19208 43868
rect 18972 42560 19024 42566
rect 18972 42502 19024 42508
rect 18880 42152 18932 42158
rect 18880 42094 18932 42100
rect 18788 42084 18840 42090
rect 18788 42026 18840 42032
rect 18604 41268 18656 41274
rect 18604 41210 18656 41216
rect 18328 41200 18380 41206
rect 18328 41142 18380 41148
rect 18236 39908 18288 39914
rect 18236 39850 18288 39856
rect 18248 37942 18276 39850
rect 18236 37936 18288 37942
rect 18236 37878 18288 37884
rect 18340 37670 18368 41142
rect 18696 40996 18748 41002
rect 18696 40938 18748 40944
rect 18708 39642 18736 40938
rect 18696 39636 18748 39642
rect 18696 39578 18748 39584
rect 18696 39364 18748 39370
rect 18696 39306 18748 39312
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18432 38962 18460 39238
rect 18512 39092 18564 39098
rect 18512 39034 18564 39040
rect 18420 38956 18472 38962
rect 18420 38898 18472 38904
rect 18524 38010 18552 39034
rect 18512 38004 18564 38010
rect 18512 37946 18564 37952
rect 18328 37664 18380 37670
rect 18328 37606 18380 37612
rect 18234 37360 18290 37369
rect 18234 37295 18236 37304
rect 18288 37295 18290 37304
rect 18236 37266 18288 37272
rect 18064 35142 18184 35170
rect 17408 35012 17460 35018
rect 17408 34954 17460 34960
rect 17420 34542 17448 34954
rect 17960 34944 18012 34950
rect 17960 34886 18012 34892
rect 17972 34746 18000 34886
rect 17960 34740 18012 34746
rect 17960 34682 18012 34688
rect 17316 34536 17368 34542
rect 17316 34478 17368 34484
rect 17408 34536 17460 34542
rect 17408 34478 17460 34484
rect 17224 34400 17276 34406
rect 17224 34342 17276 34348
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 17040 32836 17092 32842
rect 17040 32778 17092 32784
rect 16776 31726 16896 31754
rect 16776 31686 16804 31726
rect 16764 31680 16816 31686
rect 16764 31622 16816 31628
rect 16672 31272 16724 31278
rect 16672 31214 16724 31220
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16684 28762 16712 29038
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 16592 25214 16712 25242
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24206 16620 25094
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16684 24018 16712 25214
rect 16592 23990 16712 24018
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16500 20058 16528 20402
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16488 19848 16540 19854
rect 16316 19808 16488 19836
rect 16488 19790 16540 19796
rect 16500 16658 16528 19790
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 15846 15804 16154 15824
rect 15846 15802 15852 15804
rect 15908 15802 15932 15804
rect 15988 15802 16012 15804
rect 16068 15802 16092 15804
rect 16148 15802 16154 15804
rect 15908 15750 15910 15802
rect 16090 15750 16092 15802
rect 15846 15748 15852 15750
rect 15908 15748 15932 15750
rect 15988 15748 16012 15750
rect 16068 15748 16092 15750
rect 16148 15748 16154 15750
rect 15846 15728 16154 15748
rect 16592 15502 16620 23990
rect 16776 23882 16804 31078
rect 16868 29306 16896 31726
rect 16948 31204 17000 31210
rect 16948 31146 17000 31152
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16960 29238 16988 31146
rect 17052 29850 17080 32778
rect 17144 32502 17172 32846
rect 17132 32496 17184 32502
rect 17132 32438 17184 32444
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 16948 29232 17000 29238
rect 16948 29174 17000 29180
rect 17052 28558 17080 29786
rect 17040 28552 17092 28558
rect 17040 28494 17092 28500
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 27402 16988 28358
rect 16948 27396 17000 27402
rect 16948 27338 17000 27344
rect 16856 25424 16908 25430
rect 16856 25366 16908 25372
rect 16684 23854 16804 23882
rect 16684 21554 16712 23854
rect 16868 22094 16896 25366
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16960 24138 16988 24550
rect 16948 24132 17000 24138
rect 16948 24074 17000 24080
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17144 22778 17172 23054
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 16776 22066 16896 22094
rect 17236 22094 17264 34342
rect 17328 34066 17356 34478
rect 17316 34060 17368 34066
rect 17316 34002 17368 34008
rect 17420 33862 17448 34478
rect 17500 34400 17552 34406
rect 17500 34342 17552 34348
rect 17512 33998 17540 34342
rect 17868 34128 17920 34134
rect 17868 34070 17920 34076
rect 17500 33992 17552 33998
rect 17500 33934 17552 33940
rect 17408 33856 17460 33862
rect 17408 33798 17460 33804
rect 17316 33652 17368 33658
rect 17316 33594 17368 33600
rect 17328 31482 17356 33594
rect 17500 33516 17552 33522
rect 17500 33458 17552 33464
rect 17408 33448 17460 33454
rect 17408 33390 17460 33396
rect 17420 32978 17448 33390
rect 17408 32972 17460 32978
rect 17408 32914 17460 32920
rect 17420 32502 17448 32914
rect 17408 32496 17460 32502
rect 17408 32438 17460 32444
rect 17512 31754 17540 33458
rect 17684 31816 17736 31822
rect 17684 31758 17736 31764
rect 17512 31726 17632 31754
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17604 30598 17632 31726
rect 17696 30954 17724 31758
rect 17880 31754 17908 34070
rect 18064 33930 18092 35142
rect 18340 34762 18368 37606
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 18432 36650 18460 37198
rect 18420 36644 18472 36650
rect 18420 36586 18472 36592
rect 18524 35034 18552 37946
rect 18708 37505 18736 39306
rect 18892 38298 18920 42094
rect 18800 38270 18920 38298
rect 18694 37496 18750 37505
rect 18694 37431 18750 37440
rect 18432 35006 18552 35034
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 18432 34950 18460 35006
rect 18420 34944 18472 34950
rect 18420 34886 18472 34892
rect 18340 34734 18552 34762
rect 18328 34536 18380 34542
rect 18328 34478 18380 34484
rect 18052 33924 18104 33930
rect 18052 33866 18104 33872
rect 18064 32774 18092 33866
rect 18340 33454 18368 34478
rect 18328 33448 18380 33454
rect 18328 33390 18380 33396
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 18064 32570 18092 32710
rect 18052 32564 18104 32570
rect 18052 32506 18104 32512
rect 18328 32360 18380 32366
rect 18328 32302 18380 32308
rect 18144 31884 18196 31890
rect 18144 31826 18196 31832
rect 17880 31726 18092 31754
rect 17696 30926 17816 30954
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17316 28960 17368 28966
rect 17316 28902 17368 28908
rect 17328 28694 17356 28902
rect 17316 28688 17368 28694
rect 17316 28630 17368 28636
rect 17604 28626 17632 30534
rect 17788 30054 17816 30926
rect 17960 30864 18012 30870
rect 17960 30806 18012 30812
rect 17972 30326 18000 30806
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 18064 30138 18092 31726
rect 18156 31142 18184 31826
rect 18236 31816 18288 31822
rect 18340 31770 18368 32302
rect 18420 32224 18472 32230
rect 18420 32166 18472 32172
rect 18288 31764 18368 31770
rect 18236 31758 18368 31764
rect 18248 31742 18368 31758
rect 18340 31346 18368 31742
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18144 31136 18196 31142
rect 18144 31078 18196 31084
rect 17972 30110 18092 30138
rect 17776 30048 17828 30054
rect 17776 29990 17828 29996
rect 17592 28620 17644 28626
rect 17592 28562 17644 28568
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17604 26926 17632 27338
rect 17592 26920 17644 26926
rect 17592 26862 17644 26868
rect 17868 25696 17920 25702
rect 17868 25638 17920 25644
rect 17880 25226 17908 25638
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17512 23866 17540 24754
rect 17696 24410 17724 25162
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17684 24404 17736 24410
rect 17684 24346 17736 24352
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17696 23730 17724 24346
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17880 23594 17908 24686
rect 17868 23588 17920 23594
rect 17868 23530 17920 23536
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 17236 22066 17356 22094
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16684 20466 16712 21286
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16684 19514 16712 19790
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15706 16712 15846
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 15846 14716 16154 14736
rect 15846 14714 15852 14716
rect 15908 14714 15932 14716
rect 15988 14714 16012 14716
rect 16068 14714 16092 14716
rect 16148 14714 16154 14716
rect 15908 14662 15910 14714
rect 16090 14662 16092 14714
rect 15846 14660 15852 14662
rect 15908 14660 15932 14662
rect 15988 14660 16012 14662
rect 16068 14660 16092 14662
rect 16148 14660 16154 14662
rect 15846 14640 16154 14660
rect 15846 13628 16154 13648
rect 15846 13626 15852 13628
rect 15908 13626 15932 13628
rect 15988 13626 16012 13628
rect 16068 13626 16092 13628
rect 16148 13626 16154 13628
rect 15908 13574 15910 13626
rect 16090 13574 16092 13626
rect 15846 13572 15852 13574
rect 15908 13572 15932 13574
rect 15988 13572 16012 13574
rect 16068 13572 16092 13574
rect 16148 13572 16154 13574
rect 15846 13552 16154 13572
rect 15846 12540 16154 12560
rect 15846 12538 15852 12540
rect 15908 12538 15932 12540
rect 15988 12538 16012 12540
rect 16068 12538 16092 12540
rect 16148 12538 16154 12540
rect 15908 12486 15910 12538
rect 16090 12486 16092 12538
rect 15846 12484 15852 12486
rect 15908 12484 15932 12486
rect 15988 12484 16012 12486
rect 16068 12484 16092 12486
rect 16148 12484 16154 12486
rect 15846 12464 16154 12484
rect 15846 11452 16154 11472
rect 15846 11450 15852 11452
rect 15908 11450 15932 11452
rect 15988 11450 16012 11452
rect 16068 11450 16092 11452
rect 16148 11450 16154 11452
rect 15908 11398 15910 11450
rect 16090 11398 16092 11450
rect 15846 11396 15852 11398
rect 15908 11396 15932 11398
rect 15988 11396 16012 11398
rect 16068 11396 16092 11398
rect 16148 11396 16154 11398
rect 15846 11376 16154 11396
rect 15846 10364 16154 10384
rect 15846 10362 15852 10364
rect 15908 10362 15932 10364
rect 15988 10362 16012 10364
rect 16068 10362 16092 10364
rect 16148 10362 16154 10364
rect 15908 10310 15910 10362
rect 16090 10310 16092 10362
rect 15846 10308 15852 10310
rect 15908 10308 15932 10310
rect 15988 10308 16012 10310
rect 16068 10308 16092 10310
rect 16148 10308 16154 10310
rect 15846 10288 16154 10308
rect 15846 9276 16154 9296
rect 15846 9274 15852 9276
rect 15908 9274 15932 9276
rect 15988 9274 16012 9276
rect 16068 9274 16092 9276
rect 16148 9274 16154 9276
rect 15908 9222 15910 9274
rect 16090 9222 16092 9274
rect 15846 9220 15852 9222
rect 15908 9220 15932 9222
rect 15988 9220 16012 9222
rect 16068 9220 16092 9222
rect 16148 9220 16154 9222
rect 15846 9200 16154 9220
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 15846 8188 16154 8208
rect 15846 8186 15852 8188
rect 15908 8186 15932 8188
rect 15988 8186 16012 8188
rect 16068 8186 16092 8188
rect 16148 8186 16154 8188
rect 15908 8134 15910 8186
rect 16090 8134 16092 8186
rect 15846 8132 15852 8134
rect 15908 8132 15932 8134
rect 15988 8132 16012 8134
rect 16068 8132 16092 8134
rect 16148 8132 16154 8134
rect 15846 8112 16154 8132
rect 10880 7644 11188 7664
rect 10880 7642 10886 7644
rect 10942 7642 10966 7644
rect 11022 7642 11046 7644
rect 11102 7642 11126 7644
rect 11182 7642 11188 7644
rect 10942 7590 10944 7642
rect 11124 7590 11126 7642
rect 10880 7588 10886 7590
rect 10942 7588 10966 7590
rect 11022 7588 11046 7590
rect 11102 7588 11126 7590
rect 11182 7588 11188 7590
rect 10880 7568 11188 7588
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 5915 7100 6223 7120
rect 5915 7098 5921 7100
rect 5977 7098 6001 7100
rect 6057 7098 6081 7100
rect 6137 7098 6161 7100
rect 6217 7098 6223 7100
rect 5977 7046 5979 7098
rect 6159 7046 6161 7098
rect 5915 7044 5921 7046
rect 5977 7044 6001 7046
rect 6057 7044 6081 7046
rect 6137 7044 6161 7046
rect 6217 7044 6223 7046
rect 5915 7024 6223 7044
rect 15846 7100 16154 7120
rect 15846 7098 15852 7100
rect 15908 7098 15932 7100
rect 15988 7098 16012 7100
rect 16068 7098 16092 7100
rect 16148 7098 16154 7100
rect 15908 7046 15910 7098
rect 16090 7046 16092 7098
rect 15846 7044 15852 7046
rect 15908 7044 15932 7046
rect 15988 7044 16012 7046
rect 16068 7044 16092 7046
rect 16148 7044 16154 7046
rect 15846 7024 16154 7044
rect 16776 6914 16804 22066
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 16854 16824 16910 16833
rect 17236 16794 17264 17138
rect 16854 16759 16910 16768
rect 17224 16788 17276 16794
rect 16868 16658 16896 16759
rect 17224 16730 17276 16736
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16868 16114 16896 16390
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16960 15706 16988 16118
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 14618 17264 14826
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17328 12238 17356 22066
rect 17880 21690 17908 22578
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17788 19854 17816 20878
rect 17880 20398 17908 21626
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16182 17724 16934
rect 17788 16182 17816 19790
rect 17880 19446 17908 20334
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17972 16998 18000 30110
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 18340 27878 18368 28494
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 18064 25974 18092 26522
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 18340 25362 18368 27814
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18064 24818 18092 25094
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18156 23866 18184 24550
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18156 22778 18184 23802
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 18432 21554 18460 32166
rect 18524 31754 18552 34734
rect 18616 32366 18644 35022
rect 18708 34678 18736 37431
rect 18800 35086 18828 38270
rect 18880 38208 18932 38214
rect 18880 38150 18932 38156
rect 18788 35080 18840 35086
rect 18788 35022 18840 35028
rect 18696 34672 18748 34678
rect 18696 34614 18748 34620
rect 18696 32564 18748 32570
rect 18696 32506 18748 32512
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18708 31754 18736 32506
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18800 31890 18828 32370
rect 18788 31884 18840 31890
rect 18788 31826 18840 31832
rect 18524 31726 18644 31754
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18524 30598 18552 31214
rect 18512 30592 18564 30598
rect 18512 30534 18564 30540
rect 18512 25832 18564 25838
rect 18512 25774 18564 25780
rect 18524 25294 18552 25774
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18616 24886 18644 31726
rect 18696 31748 18748 31754
rect 18696 31690 18748 31696
rect 18788 31136 18840 31142
rect 18788 31078 18840 31084
rect 18696 30728 18748 30734
rect 18696 30670 18748 30676
rect 18708 30394 18736 30670
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 18708 29850 18736 30194
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18800 29646 18828 31078
rect 18788 29640 18840 29646
rect 18788 29582 18840 29588
rect 18892 27062 18920 38150
rect 18970 37360 19026 37369
rect 18970 37295 18972 37304
rect 19024 37295 19026 37304
rect 18972 37266 19024 37272
rect 18972 36780 19024 36786
rect 18972 36722 19024 36728
rect 18984 33114 19012 36722
rect 19064 34944 19116 34950
rect 19064 34886 19116 34892
rect 19076 34746 19104 34886
rect 19064 34740 19116 34746
rect 19064 34682 19116 34688
rect 18972 33108 19024 33114
rect 18972 33050 19024 33056
rect 19076 32842 19104 34682
rect 19064 32836 19116 32842
rect 19064 32778 19116 32784
rect 19076 32570 19104 32778
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18972 31952 19024 31958
rect 18972 31894 19024 31900
rect 18984 30802 19012 31894
rect 19064 31136 19116 31142
rect 19064 31078 19116 31084
rect 18972 30796 19024 30802
rect 18972 30738 19024 30744
rect 19076 30734 19104 31078
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 18972 30048 19024 30054
rect 18972 29990 19024 29996
rect 18880 27056 18932 27062
rect 18880 26998 18932 27004
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18984 24274 19012 29990
rect 19076 29073 19104 30194
rect 19062 29064 19118 29073
rect 19062 28999 19118 29008
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18524 23730 18552 24142
rect 19168 23730 19196 43862
rect 19248 43716 19300 43722
rect 19248 43658 19300 43664
rect 19260 42362 19288 43658
rect 19248 42356 19300 42362
rect 19248 42298 19300 42304
rect 19352 41682 19380 44814
rect 19340 41676 19392 41682
rect 19340 41618 19392 41624
rect 19340 41132 19392 41138
rect 19340 41074 19392 41080
rect 19352 40730 19380 41074
rect 19340 40724 19392 40730
rect 19340 40666 19392 40672
rect 19340 38752 19392 38758
rect 19340 38694 19392 38700
rect 19352 38350 19380 38694
rect 19340 38344 19392 38350
rect 19340 38286 19392 38292
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 19260 36378 19288 37198
rect 19340 36576 19392 36582
rect 19340 36518 19392 36524
rect 19248 36372 19300 36378
rect 19248 36314 19300 36320
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19260 35290 19288 36110
rect 19248 35284 19300 35290
rect 19248 35226 19300 35232
rect 19352 25906 19380 36518
rect 19444 33946 19472 44950
rect 19536 44470 19564 45222
rect 19524 44464 19576 44470
rect 19524 44406 19576 44412
rect 19524 44328 19576 44334
rect 19524 44270 19576 44276
rect 19536 42022 19564 44270
rect 19628 43382 19656 47126
rect 19720 43994 19748 47518
rect 19800 47524 19852 47530
rect 19800 47466 19852 47472
rect 19904 46170 19932 51046
rect 20168 50720 20220 50726
rect 20168 50662 20220 50668
rect 19984 50312 20036 50318
rect 19984 50254 20036 50260
rect 19996 49978 20024 50254
rect 19984 49972 20036 49978
rect 19984 49914 20036 49920
rect 20076 49088 20128 49094
rect 20180 49076 20208 50662
rect 20128 49048 20208 49076
rect 20076 49030 20128 49036
rect 20180 48822 20208 49048
rect 20168 48816 20220 48822
rect 20168 48758 20220 48764
rect 19984 47660 20036 47666
rect 19984 47602 20036 47608
rect 19892 46164 19944 46170
rect 19892 46106 19944 46112
rect 19892 45892 19944 45898
rect 19892 45834 19944 45840
rect 19800 44940 19852 44946
rect 19800 44882 19852 44888
rect 19708 43988 19760 43994
rect 19708 43930 19760 43936
rect 19812 43858 19840 44882
rect 19904 44538 19932 45834
rect 19996 45354 20024 47602
rect 20076 46912 20128 46918
rect 20076 46854 20128 46860
rect 19984 45348 20036 45354
rect 19984 45290 20036 45296
rect 19984 44804 20036 44810
rect 19984 44746 20036 44752
rect 19892 44532 19944 44538
rect 19892 44474 19944 44480
rect 19892 43920 19944 43926
rect 19892 43862 19944 43868
rect 19800 43852 19852 43858
rect 19800 43794 19852 43800
rect 19708 43444 19760 43450
rect 19708 43386 19760 43392
rect 19616 43376 19668 43382
rect 19616 43318 19668 43324
rect 19720 43194 19748 43386
rect 19628 43166 19748 43194
rect 19524 42016 19576 42022
rect 19524 41958 19576 41964
rect 19524 41472 19576 41478
rect 19524 41414 19576 41420
rect 19536 39030 19564 41414
rect 19628 41206 19656 43166
rect 19904 42650 19932 43862
rect 19996 43790 20024 44746
rect 19984 43784 20036 43790
rect 19984 43726 20036 43732
rect 20088 42702 20116 46854
rect 20180 43654 20208 48758
rect 20168 43648 20220 43654
rect 20168 43590 20220 43596
rect 19812 42622 19932 42650
rect 20076 42696 20128 42702
rect 20076 42638 20128 42644
rect 19708 41540 19760 41546
rect 19708 41482 19760 41488
rect 19720 41206 19748 41482
rect 19616 41200 19668 41206
rect 19616 41142 19668 41148
rect 19708 41200 19760 41206
rect 19708 41142 19760 41148
rect 19616 40384 19668 40390
rect 19616 40326 19668 40332
rect 19628 39930 19656 40326
rect 19720 40118 19748 41142
rect 19708 40112 19760 40118
rect 19708 40054 19760 40060
rect 19628 39902 19748 39930
rect 19616 39840 19668 39846
rect 19616 39782 19668 39788
rect 19524 39024 19576 39030
rect 19524 38966 19576 38972
rect 19628 37874 19656 39782
rect 19616 37868 19668 37874
rect 19616 37810 19668 37816
rect 19524 35692 19576 35698
rect 19720 35680 19748 39902
rect 19812 36582 19840 42622
rect 20076 42220 20128 42226
rect 20076 42162 20128 42168
rect 19892 41608 19944 41614
rect 19892 41550 19944 41556
rect 19904 41002 19932 41550
rect 20088 41546 20116 42162
rect 20272 42106 20300 55150
rect 20444 54732 20496 54738
rect 20444 54674 20496 54680
rect 20456 52578 20484 54674
rect 20548 52698 20576 57530
rect 21088 57520 21140 57526
rect 20810 57488 20866 57497
rect 20628 57452 20680 57458
rect 21088 57462 21140 57468
rect 20810 57423 20812 57432
rect 20628 57394 20680 57400
rect 20864 57423 20866 57432
rect 20812 57394 20864 57400
rect 20640 56710 20668 57394
rect 20720 57316 20772 57322
rect 20720 57258 20772 57264
rect 20628 56704 20680 56710
rect 20628 56646 20680 56652
rect 20640 55214 20668 56646
rect 20732 55418 20760 57258
rect 21100 57050 21128 57462
rect 21088 57044 21140 57050
rect 21088 56986 21140 56992
rect 20811 56604 21119 56624
rect 20811 56602 20817 56604
rect 20873 56602 20897 56604
rect 20953 56602 20977 56604
rect 21033 56602 21057 56604
rect 21113 56602 21119 56604
rect 20873 56550 20875 56602
rect 21055 56550 21057 56602
rect 20811 56548 20817 56550
rect 20873 56548 20897 56550
rect 20953 56548 20977 56550
rect 21033 56548 21057 56550
rect 21113 56548 21119 56550
rect 20811 56528 21119 56548
rect 21192 55962 21220 58414
rect 21284 57322 21312 63174
rect 21376 59226 21404 66226
rect 22204 66212 22232 69226
rect 22296 69018 22324 69838
rect 22388 69494 22416 70366
rect 22376 69488 22428 69494
rect 22376 69430 22428 69436
rect 22480 69426 22508 71402
rect 22468 69420 22520 69426
rect 22468 69362 22520 69368
rect 22284 69012 22336 69018
rect 22284 68954 22336 68960
rect 22468 68196 22520 68202
rect 22468 68138 22520 68144
rect 22376 66224 22428 66230
rect 22204 66184 22376 66212
rect 21916 66156 21968 66162
rect 21916 66098 21968 66104
rect 21824 65952 21876 65958
rect 21824 65894 21876 65900
rect 21836 65142 21864 65894
rect 21928 65210 21956 66098
rect 21916 65204 21968 65210
rect 21916 65146 21968 65152
rect 21824 65136 21876 65142
rect 21824 65078 21876 65084
rect 21548 64864 21600 64870
rect 21548 64806 21600 64812
rect 21560 60722 21588 64806
rect 21640 64592 21692 64598
rect 21640 64534 21692 64540
rect 21652 64462 21680 64534
rect 21640 64456 21692 64462
rect 21640 64398 21692 64404
rect 21916 64388 21968 64394
rect 22204 64376 22232 66184
rect 22376 66166 22428 66172
rect 22376 66088 22428 66094
rect 22376 66030 22428 66036
rect 22388 64598 22416 66030
rect 22376 64592 22428 64598
rect 22376 64534 22428 64540
rect 21968 64348 22232 64376
rect 21916 64330 21968 64336
rect 21824 62212 21876 62218
rect 21824 62154 21876 62160
rect 21836 61946 21864 62154
rect 21824 61940 21876 61946
rect 21824 61882 21876 61888
rect 21928 61724 21956 64330
rect 22100 62348 22152 62354
rect 22100 62290 22152 62296
rect 22112 61810 22140 62290
rect 22388 61878 22416 64534
rect 22376 61872 22428 61878
rect 22376 61814 22428 61820
rect 22480 61810 22508 68138
rect 22560 66836 22612 66842
rect 22560 66778 22612 66784
rect 22572 66638 22600 66778
rect 22560 66632 22612 66638
rect 22560 66574 22612 66580
rect 22558 66192 22614 66201
rect 22558 66127 22560 66136
rect 22612 66127 22614 66136
rect 22560 66098 22612 66104
rect 22664 66065 22692 74054
rect 22848 73574 22876 74598
rect 22836 73568 22888 73574
rect 22836 73510 22888 73516
rect 22848 66706 22876 73510
rect 24216 70100 24268 70106
rect 24216 70042 24268 70048
rect 23572 67244 23624 67250
rect 23572 67186 23624 67192
rect 23584 66842 23612 67186
rect 23940 67040 23992 67046
rect 23940 66982 23992 66988
rect 23572 66836 23624 66842
rect 23572 66778 23624 66784
rect 23296 66768 23348 66774
rect 23296 66710 23348 66716
rect 22836 66700 22888 66706
rect 22836 66642 22888 66648
rect 23020 66224 23072 66230
rect 23020 66166 23072 66172
rect 22650 66056 22706 66065
rect 22650 65991 22706 66000
rect 22744 65408 22796 65414
rect 22744 65350 22796 65356
rect 22756 64462 22784 65350
rect 22744 64456 22796 64462
rect 22744 64398 22796 64404
rect 22928 63980 22980 63986
rect 22928 63922 22980 63928
rect 22100 61804 22152 61810
rect 22100 61746 22152 61752
rect 22468 61804 22520 61810
rect 22468 61746 22520 61752
rect 22008 61736 22060 61742
rect 21928 61696 22008 61724
rect 22008 61678 22060 61684
rect 22020 60790 22048 61678
rect 22836 61600 22888 61606
rect 22836 61542 22888 61548
rect 22376 61192 22428 61198
rect 22376 61134 22428 61140
rect 22008 60784 22060 60790
rect 22388 60761 22416 61134
rect 22652 60784 22704 60790
rect 22008 60726 22060 60732
rect 22374 60752 22430 60761
rect 21548 60716 21600 60722
rect 22652 60726 22704 60732
rect 22374 60687 22430 60696
rect 21548 60658 21600 60664
rect 22100 60512 22152 60518
rect 22100 60454 22152 60460
rect 21732 60308 21784 60314
rect 21732 60250 21784 60256
rect 21456 60036 21508 60042
rect 21456 59978 21508 59984
rect 21364 59220 21416 59226
rect 21364 59162 21416 59168
rect 21272 57316 21324 57322
rect 21272 57258 21324 57264
rect 21376 56982 21404 59162
rect 21364 56976 21416 56982
rect 21364 56918 21416 56924
rect 21272 56840 21324 56846
rect 21272 56782 21324 56788
rect 21284 55962 21312 56782
rect 21180 55956 21232 55962
rect 21180 55898 21232 55904
rect 21272 55956 21324 55962
rect 21272 55898 21324 55904
rect 20811 55516 21119 55536
rect 20811 55514 20817 55516
rect 20873 55514 20897 55516
rect 20953 55514 20977 55516
rect 21033 55514 21057 55516
rect 21113 55514 21119 55516
rect 20873 55462 20875 55514
rect 21055 55462 21057 55514
rect 20811 55460 20817 55462
rect 20873 55460 20897 55462
rect 20953 55460 20977 55462
rect 21033 55460 21057 55462
rect 21113 55460 21119 55462
rect 20811 55440 21119 55460
rect 20720 55412 20772 55418
rect 20720 55354 20772 55360
rect 20628 55208 20680 55214
rect 20628 55150 20680 55156
rect 20811 54428 21119 54448
rect 20811 54426 20817 54428
rect 20873 54426 20897 54428
rect 20953 54426 20977 54428
rect 21033 54426 21057 54428
rect 21113 54426 21119 54428
rect 20873 54374 20875 54426
rect 21055 54374 21057 54426
rect 20811 54372 20817 54374
rect 20873 54372 20897 54374
rect 20953 54372 20977 54374
rect 21033 54372 21057 54374
rect 21113 54372 21119 54374
rect 20811 54352 21119 54372
rect 21192 53514 21220 55898
rect 21272 55276 21324 55282
rect 21272 55218 21324 55224
rect 21180 53508 21232 53514
rect 21180 53450 21232 53456
rect 21284 53446 21312 55218
rect 21272 53440 21324 53446
rect 21272 53382 21324 53388
rect 20811 53340 21119 53360
rect 20811 53338 20817 53340
rect 20873 53338 20897 53340
rect 20953 53338 20977 53340
rect 21033 53338 21057 53340
rect 21113 53338 21119 53340
rect 20873 53286 20875 53338
rect 21055 53286 21057 53338
rect 20811 53284 20817 53286
rect 20873 53284 20897 53286
rect 20953 53284 20977 53286
rect 21033 53284 21057 53286
rect 21113 53284 21119 53286
rect 20811 53264 21119 53284
rect 20720 53168 20772 53174
rect 20720 53110 20772 53116
rect 20628 52896 20680 52902
rect 20628 52838 20680 52844
rect 20536 52692 20588 52698
rect 20536 52634 20588 52640
rect 20456 52550 20576 52578
rect 20640 52562 20668 52838
rect 20444 52352 20496 52358
rect 20444 52294 20496 52300
rect 20352 51060 20404 51066
rect 20352 51002 20404 51008
rect 20364 49842 20392 51002
rect 20352 49836 20404 49842
rect 20352 49778 20404 49784
rect 20352 49156 20404 49162
rect 20352 49098 20404 49104
rect 20364 48686 20392 49098
rect 20352 48680 20404 48686
rect 20352 48622 20404 48628
rect 20352 48136 20404 48142
rect 20350 48104 20352 48113
rect 20404 48104 20406 48113
rect 20350 48039 20406 48048
rect 20352 48000 20404 48006
rect 20352 47942 20404 47948
rect 20364 45626 20392 47942
rect 20352 45620 20404 45626
rect 20352 45562 20404 45568
rect 20272 42078 20392 42106
rect 20260 42016 20312 42022
rect 20260 41958 20312 41964
rect 20168 41676 20220 41682
rect 20168 41618 20220 41624
rect 20076 41540 20128 41546
rect 20076 41482 20128 41488
rect 19984 41268 20036 41274
rect 19984 41210 20036 41216
rect 19892 40996 19944 41002
rect 19892 40938 19944 40944
rect 19890 40624 19946 40633
rect 19890 40559 19892 40568
rect 19944 40559 19946 40568
rect 19892 40530 19944 40536
rect 19996 40186 20024 41210
rect 19984 40180 20036 40186
rect 19984 40122 20036 40128
rect 20088 40066 20116 41482
rect 20180 41070 20208 41618
rect 20168 41064 20220 41070
rect 20168 41006 20220 41012
rect 19996 40038 20116 40066
rect 19996 38350 20024 40038
rect 20168 39296 20220 39302
rect 20168 39238 20220 39244
rect 20180 38962 20208 39238
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 20168 38956 20220 38962
rect 20168 38898 20220 38904
rect 19984 38344 20036 38350
rect 19984 38286 20036 38292
rect 19890 37360 19946 37369
rect 19890 37295 19946 37304
rect 19904 37194 19932 37295
rect 19892 37188 19944 37194
rect 19892 37130 19944 37136
rect 19892 36644 19944 36650
rect 19892 36586 19944 36592
rect 19800 36576 19852 36582
rect 19800 36518 19852 36524
rect 19524 35634 19576 35640
rect 19628 35652 19748 35680
rect 19536 34134 19564 35634
rect 19628 34898 19656 35652
rect 19708 35556 19760 35562
rect 19708 35498 19760 35504
rect 19720 35290 19748 35498
rect 19800 35488 19852 35494
rect 19800 35430 19852 35436
rect 19708 35284 19760 35290
rect 19708 35226 19760 35232
rect 19720 35057 19748 35226
rect 19706 35048 19762 35057
rect 19812 35018 19840 35430
rect 19706 34983 19762 34992
rect 19800 35012 19852 35018
rect 19800 34954 19852 34960
rect 19628 34870 19840 34898
rect 19706 34640 19762 34649
rect 19616 34604 19668 34610
rect 19706 34575 19762 34584
rect 19616 34546 19668 34552
rect 19628 34202 19656 34546
rect 19616 34196 19668 34202
rect 19616 34138 19668 34144
rect 19524 34128 19576 34134
rect 19524 34070 19576 34076
rect 19444 33918 19656 33946
rect 19432 33856 19484 33862
rect 19432 33798 19484 33804
rect 19444 33522 19472 33798
rect 19524 33584 19576 33590
rect 19524 33526 19576 33532
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19444 32910 19472 33458
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 19536 31414 19564 33526
rect 19524 31408 19576 31414
rect 19524 31350 19576 31356
rect 19628 30734 19656 33918
rect 19720 32978 19748 34575
rect 19708 32972 19760 32978
rect 19708 32914 19760 32920
rect 19616 30728 19668 30734
rect 19616 30670 19668 30676
rect 19524 30592 19576 30598
rect 19524 30534 19576 30540
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 19444 27878 19472 30262
rect 19536 29170 19564 30534
rect 19812 30326 19840 34870
rect 19904 34542 19932 36586
rect 19892 34536 19944 34542
rect 19892 34478 19944 34484
rect 19892 34128 19944 34134
rect 19892 34070 19944 34076
rect 19904 33590 19932 34070
rect 19996 33998 20024 38286
rect 20088 36582 20116 38898
rect 20168 37664 20220 37670
rect 20168 37606 20220 37612
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 20088 34678 20116 36518
rect 20076 34672 20128 34678
rect 20076 34614 20128 34620
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 19892 33584 19944 33590
rect 19892 33526 19944 33532
rect 19892 32428 19944 32434
rect 19892 32370 19944 32376
rect 19904 32026 19932 32370
rect 19892 32020 19944 32026
rect 19892 31962 19944 31968
rect 19996 31890 20024 33934
rect 20180 32502 20208 37606
rect 20272 34762 20300 41958
rect 20364 36242 20392 42078
rect 20456 41414 20484 52294
rect 20548 50425 20576 52550
rect 20628 52556 20680 52562
rect 20628 52498 20680 52504
rect 20640 51406 20668 52498
rect 20732 52494 20760 53110
rect 20720 52488 20772 52494
rect 20720 52430 20772 52436
rect 20732 52018 20760 52430
rect 20811 52252 21119 52272
rect 20811 52250 20817 52252
rect 20873 52250 20897 52252
rect 20953 52250 20977 52252
rect 21033 52250 21057 52252
rect 21113 52250 21119 52252
rect 20873 52198 20875 52250
rect 21055 52198 21057 52250
rect 20811 52196 20817 52198
rect 20873 52196 20897 52198
rect 20953 52196 20977 52198
rect 21033 52196 21057 52198
rect 21113 52196 21119 52198
rect 20811 52176 21119 52196
rect 20720 52012 20772 52018
rect 20720 51954 20772 51960
rect 20628 51400 20680 51406
rect 20628 51342 20680 51348
rect 20628 51264 20680 51270
rect 20628 51206 20680 51212
rect 20534 50416 20590 50425
rect 20534 50351 20590 50360
rect 20640 49366 20668 51206
rect 20811 51164 21119 51184
rect 20811 51162 20817 51164
rect 20873 51162 20897 51164
rect 20953 51162 20977 51164
rect 21033 51162 21057 51164
rect 21113 51162 21119 51164
rect 20873 51110 20875 51162
rect 21055 51110 21057 51162
rect 20811 51108 20817 51110
rect 20873 51108 20897 51110
rect 20953 51108 20977 51110
rect 21033 51108 21057 51110
rect 21113 51108 21119 51110
rect 20811 51088 21119 51108
rect 21284 50998 21312 53382
rect 21364 51264 21416 51270
rect 21364 51206 21416 51212
rect 21272 50992 21324 50998
rect 21086 50960 21142 50969
rect 21272 50934 21324 50940
rect 21086 50895 21142 50904
rect 21100 50318 21128 50895
rect 21088 50312 21140 50318
rect 21088 50254 21140 50260
rect 20811 50076 21119 50096
rect 20811 50074 20817 50076
rect 20873 50074 20897 50076
rect 20953 50074 20977 50076
rect 21033 50074 21057 50076
rect 21113 50074 21119 50076
rect 20873 50022 20875 50074
rect 21055 50022 21057 50074
rect 20811 50020 20817 50022
rect 20873 50020 20897 50022
rect 20953 50020 20977 50022
rect 21033 50020 21057 50022
rect 21113 50020 21119 50022
rect 20811 50000 21119 50020
rect 20628 49360 20680 49366
rect 20628 49302 20680 49308
rect 21272 49156 21324 49162
rect 21272 49098 21324 49104
rect 20720 49088 20772 49094
rect 20720 49030 20772 49036
rect 20732 48822 20760 49030
rect 20811 48988 21119 49008
rect 20811 48986 20817 48988
rect 20873 48986 20897 48988
rect 20953 48986 20977 48988
rect 21033 48986 21057 48988
rect 21113 48986 21119 48988
rect 20873 48934 20875 48986
rect 21055 48934 21057 48986
rect 20811 48932 20817 48934
rect 20873 48932 20897 48934
rect 20953 48932 20977 48934
rect 21033 48932 21057 48934
rect 21113 48932 21119 48934
rect 20811 48912 21119 48932
rect 20720 48816 20772 48822
rect 20720 48758 20772 48764
rect 20628 48544 20680 48550
rect 20628 48486 20680 48492
rect 20536 48000 20588 48006
rect 20536 47942 20588 47948
rect 20548 47258 20576 47942
rect 20536 47252 20588 47258
rect 20536 47194 20588 47200
rect 20536 46980 20588 46986
rect 20536 46922 20588 46928
rect 20548 43450 20576 46922
rect 20640 44810 20668 48486
rect 20732 48142 20760 48758
rect 20720 48136 20772 48142
rect 20720 48078 20772 48084
rect 20811 47900 21119 47920
rect 20811 47898 20817 47900
rect 20873 47898 20897 47900
rect 20953 47898 20977 47900
rect 21033 47898 21057 47900
rect 21113 47898 21119 47900
rect 20873 47846 20875 47898
rect 21055 47846 21057 47898
rect 20811 47844 20817 47846
rect 20873 47844 20897 47846
rect 20953 47844 20977 47846
rect 21033 47844 21057 47846
rect 21113 47844 21119 47846
rect 20811 47824 21119 47844
rect 20720 47456 20772 47462
rect 20720 47398 20772 47404
rect 20732 46034 20760 47398
rect 21180 46980 21232 46986
rect 21180 46922 21232 46928
rect 20811 46812 21119 46832
rect 20811 46810 20817 46812
rect 20873 46810 20897 46812
rect 20953 46810 20977 46812
rect 21033 46810 21057 46812
rect 21113 46810 21119 46812
rect 20873 46758 20875 46810
rect 21055 46758 21057 46810
rect 20811 46756 20817 46758
rect 20873 46756 20897 46758
rect 20953 46756 20977 46758
rect 21033 46756 21057 46758
rect 21113 46756 21119 46758
rect 20811 46736 21119 46756
rect 20720 46028 20772 46034
rect 20720 45970 20772 45976
rect 20811 45724 21119 45744
rect 20811 45722 20817 45724
rect 20873 45722 20897 45724
rect 20953 45722 20977 45724
rect 21033 45722 21057 45724
rect 21113 45722 21119 45724
rect 20873 45670 20875 45722
rect 21055 45670 21057 45722
rect 20811 45668 20817 45670
rect 20873 45668 20897 45670
rect 20953 45668 20977 45670
rect 21033 45668 21057 45670
rect 21113 45668 21119 45670
rect 20811 45648 21119 45668
rect 21192 45558 21220 46922
rect 21284 46646 21312 49098
rect 21272 46640 21324 46646
rect 21272 46582 21324 46588
rect 21180 45552 21232 45558
rect 21180 45494 21232 45500
rect 20720 45484 20772 45490
rect 20720 45426 20772 45432
rect 20628 44804 20680 44810
rect 20628 44746 20680 44752
rect 20628 44532 20680 44538
rect 20628 44474 20680 44480
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 20640 43246 20668 44474
rect 20628 43240 20680 43246
rect 20628 43182 20680 43188
rect 20628 42220 20680 42226
rect 20628 42162 20680 42168
rect 20640 41818 20668 42162
rect 20628 41812 20680 41818
rect 20628 41754 20680 41760
rect 20732 41614 20760 45426
rect 20904 45416 20956 45422
rect 20904 45358 20956 45364
rect 20996 45416 21048 45422
rect 20996 45358 21048 45364
rect 20916 45014 20944 45358
rect 20904 45008 20956 45014
rect 20904 44950 20956 44956
rect 21008 44946 21036 45358
rect 20996 44940 21048 44946
rect 20996 44882 21048 44888
rect 21192 44742 21220 45494
rect 21180 44736 21232 44742
rect 21180 44678 21232 44684
rect 20811 44636 21119 44656
rect 20811 44634 20817 44636
rect 20873 44634 20897 44636
rect 20953 44634 20977 44636
rect 21033 44634 21057 44636
rect 21113 44634 21119 44636
rect 20873 44582 20875 44634
rect 21055 44582 21057 44634
rect 20811 44580 20817 44582
rect 20873 44580 20897 44582
rect 20953 44580 20977 44582
rect 21033 44580 21057 44582
rect 21113 44580 21119 44582
rect 20811 44560 21119 44580
rect 21284 44470 21312 46582
rect 21272 44464 21324 44470
rect 21272 44406 21324 44412
rect 20996 44192 21048 44198
rect 20996 44134 21048 44140
rect 21008 43858 21036 44134
rect 20996 43852 21048 43858
rect 20996 43794 21048 43800
rect 20811 43548 21119 43568
rect 20811 43546 20817 43548
rect 20873 43546 20897 43548
rect 20953 43546 20977 43548
rect 21033 43546 21057 43548
rect 21113 43546 21119 43548
rect 20873 43494 20875 43546
rect 21055 43494 21057 43546
rect 20811 43492 20817 43494
rect 20873 43492 20897 43494
rect 20953 43492 20977 43494
rect 21033 43492 21057 43494
rect 21113 43492 21119 43494
rect 20811 43472 21119 43492
rect 21376 43110 21404 51206
rect 21468 50522 21496 59978
rect 21744 59430 21772 60250
rect 21916 60036 21968 60042
rect 21916 59978 21968 59984
rect 21732 59424 21784 59430
rect 21732 59366 21784 59372
rect 21824 59152 21876 59158
rect 21824 59094 21876 59100
rect 21640 58608 21692 58614
rect 21640 58550 21692 58556
rect 21548 58064 21600 58070
rect 21548 58006 21600 58012
rect 21560 57254 21588 58006
rect 21548 57248 21600 57254
rect 21548 57190 21600 57196
rect 21548 57044 21600 57050
rect 21548 56986 21600 56992
rect 21560 56846 21588 56986
rect 21548 56840 21600 56846
rect 21548 56782 21600 56788
rect 21548 56160 21600 56166
rect 21548 56102 21600 56108
rect 21560 51097 21588 56102
rect 21546 51088 21602 51097
rect 21546 51023 21602 51032
rect 21546 50960 21602 50969
rect 21546 50895 21602 50904
rect 21456 50516 21508 50522
rect 21456 50458 21508 50464
rect 21560 50182 21588 50895
rect 21652 50454 21680 58550
rect 21732 57384 21784 57390
rect 21732 57326 21784 57332
rect 21744 52630 21772 57326
rect 21836 56846 21864 59094
rect 21824 56840 21876 56846
rect 21824 56782 21876 56788
rect 21824 56704 21876 56710
rect 21824 56646 21876 56652
rect 21836 55894 21864 56646
rect 21824 55888 21876 55894
rect 21824 55830 21876 55836
rect 21928 55706 21956 59978
rect 22112 56794 22140 60454
rect 22388 60314 22416 60687
rect 22376 60308 22428 60314
rect 22376 60250 22428 60256
rect 22560 56976 22612 56982
rect 22560 56918 22612 56924
rect 22020 56766 22140 56794
rect 22020 56250 22048 56766
rect 22100 56704 22152 56710
rect 22100 56646 22152 56652
rect 22468 56704 22520 56710
rect 22468 56646 22520 56652
rect 22112 56370 22140 56646
rect 22480 56506 22508 56646
rect 22468 56500 22520 56506
rect 22468 56442 22520 56448
rect 22100 56364 22152 56370
rect 22100 56306 22152 56312
rect 22020 56222 22140 56250
rect 21836 55678 21956 55706
rect 21836 54874 21864 55678
rect 21916 55616 21968 55622
rect 21916 55558 21968 55564
rect 21824 54868 21876 54874
rect 21824 54810 21876 54816
rect 21928 53122 21956 55558
rect 22112 55434 22140 56222
rect 22468 55752 22520 55758
rect 22468 55694 22520 55700
rect 22112 55406 22232 55434
rect 22100 54596 22152 54602
rect 22100 54538 22152 54544
rect 22112 53242 22140 54538
rect 22204 53718 22232 55406
rect 22480 54890 22508 55694
rect 22572 55622 22600 56918
rect 22560 55616 22612 55622
rect 22560 55558 22612 55564
rect 22480 54862 22600 54890
rect 22284 54528 22336 54534
rect 22284 54470 22336 54476
rect 22192 53712 22244 53718
rect 22192 53654 22244 53660
rect 22100 53236 22152 53242
rect 22100 53178 22152 53184
rect 21824 53100 21876 53106
rect 21928 53094 22048 53122
rect 21824 53042 21876 53048
rect 21732 52624 21784 52630
rect 21732 52566 21784 52572
rect 21732 51944 21784 51950
rect 21732 51886 21784 51892
rect 21744 50522 21772 51886
rect 21732 50516 21784 50522
rect 21732 50458 21784 50464
rect 21640 50448 21692 50454
rect 21640 50390 21692 50396
rect 21640 50312 21692 50318
rect 21640 50254 21692 50260
rect 21548 50176 21600 50182
rect 21548 50118 21600 50124
rect 21548 49632 21600 49638
rect 21548 49574 21600 49580
rect 21560 48822 21588 49574
rect 21548 48816 21600 48822
rect 21548 48758 21600 48764
rect 21652 48498 21680 50254
rect 21744 49230 21772 50458
rect 21732 49224 21784 49230
rect 21732 49166 21784 49172
rect 21730 48648 21786 48657
rect 21730 48583 21786 48592
rect 21560 48470 21680 48498
rect 21456 46368 21508 46374
rect 21456 46310 21508 46316
rect 21364 43104 21416 43110
rect 21364 43046 21416 43052
rect 20811 42460 21119 42480
rect 20811 42458 20817 42460
rect 20873 42458 20897 42460
rect 20953 42458 20977 42460
rect 21033 42458 21057 42460
rect 21113 42458 21119 42460
rect 20873 42406 20875 42458
rect 21055 42406 21057 42458
rect 20811 42404 20817 42406
rect 20873 42404 20897 42406
rect 20953 42404 20977 42406
rect 21033 42404 21057 42406
rect 21113 42404 21119 42406
rect 20811 42384 21119 42404
rect 21364 42356 21416 42362
rect 21364 42298 21416 42304
rect 20720 41608 20772 41614
rect 20720 41550 20772 41556
rect 20720 41472 20772 41478
rect 20720 41414 20772 41420
rect 20456 41386 20576 41414
rect 20444 41064 20496 41070
rect 20444 41006 20496 41012
rect 20456 40118 20484 41006
rect 20444 40112 20496 40118
rect 20444 40054 20496 40060
rect 20352 36236 20404 36242
rect 20352 36178 20404 36184
rect 20352 36032 20404 36038
rect 20352 35974 20404 35980
rect 20364 35698 20392 35974
rect 20548 35834 20576 41386
rect 20732 39506 20760 41414
rect 20811 41372 21119 41392
rect 20811 41370 20817 41372
rect 20873 41370 20897 41372
rect 20953 41370 20977 41372
rect 21033 41370 21057 41372
rect 21113 41370 21119 41372
rect 20873 41318 20875 41370
rect 21055 41318 21057 41370
rect 20811 41316 20817 41318
rect 20873 41316 20897 41318
rect 20953 41316 20977 41318
rect 21033 41316 21057 41318
rect 21113 41316 21119 41318
rect 20811 41296 21119 41316
rect 21376 41256 21404 42298
rect 21468 42022 21496 46310
rect 21456 42016 21508 42022
rect 21456 41958 21508 41964
rect 21376 41228 21496 41256
rect 21364 41132 21416 41138
rect 21364 41074 21416 41080
rect 21180 40996 21232 41002
rect 21180 40938 21232 40944
rect 20811 40284 21119 40304
rect 20811 40282 20817 40284
rect 20873 40282 20897 40284
rect 20953 40282 20977 40284
rect 21033 40282 21057 40284
rect 21113 40282 21119 40284
rect 20873 40230 20875 40282
rect 21055 40230 21057 40282
rect 20811 40228 20817 40230
rect 20873 40228 20897 40230
rect 20953 40228 20977 40230
rect 21033 40228 21057 40230
rect 21113 40228 21119 40230
rect 20811 40208 21119 40228
rect 21192 40050 21220 40938
rect 21272 40928 21324 40934
rect 21270 40896 21272 40905
rect 21324 40896 21326 40905
rect 21270 40831 21326 40840
rect 21180 40044 21232 40050
rect 21180 39986 21232 39992
rect 20720 39500 20772 39506
rect 20720 39442 20772 39448
rect 20811 39196 21119 39216
rect 20811 39194 20817 39196
rect 20873 39194 20897 39196
rect 20953 39194 20977 39196
rect 21033 39194 21057 39196
rect 21113 39194 21119 39196
rect 20873 39142 20875 39194
rect 21055 39142 21057 39194
rect 20811 39140 20817 39142
rect 20873 39140 20897 39142
rect 20953 39140 20977 39142
rect 21033 39140 21057 39142
rect 21113 39140 21119 39142
rect 20811 39120 21119 39140
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 20824 38554 20852 38966
rect 21088 38820 21140 38826
rect 21088 38762 21140 38768
rect 21100 38554 21128 38762
rect 20812 38548 20864 38554
rect 20812 38490 20864 38496
rect 21088 38548 21140 38554
rect 21088 38490 21140 38496
rect 20811 38108 21119 38128
rect 20811 38106 20817 38108
rect 20873 38106 20897 38108
rect 20953 38106 20977 38108
rect 21033 38106 21057 38108
rect 21113 38106 21119 38108
rect 20873 38054 20875 38106
rect 21055 38054 21057 38106
rect 20811 38052 20817 38054
rect 20873 38052 20897 38054
rect 20953 38052 20977 38054
rect 21033 38052 21057 38054
rect 21113 38052 21119 38054
rect 20811 38032 21119 38052
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 20811 37020 21119 37040
rect 20811 37018 20817 37020
rect 20873 37018 20897 37020
rect 20953 37018 20977 37020
rect 21033 37018 21057 37020
rect 21113 37018 21119 37020
rect 20873 36966 20875 37018
rect 21055 36966 21057 37018
rect 20811 36964 20817 36966
rect 20873 36964 20897 36966
rect 20953 36964 20977 36966
rect 21033 36964 21057 36966
rect 21113 36964 21119 36966
rect 20811 36944 21119 36964
rect 21180 36780 21232 36786
rect 21180 36722 21232 36728
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20536 35828 20588 35834
rect 20536 35770 20588 35776
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20272 34734 20392 34762
rect 20456 34746 20484 35022
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20272 33114 20300 34546
rect 20260 33108 20312 33114
rect 20260 33050 20312 33056
rect 20168 32496 20220 32502
rect 20168 32438 20220 32444
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 19892 30388 19944 30394
rect 19892 30330 19944 30336
rect 19800 30320 19852 30326
rect 19720 30280 19800 30308
rect 19616 29232 19668 29238
rect 19614 29200 19616 29209
rect 19668 29200 19670 29209
rect 19524 29164 19576 29170
rect 19614 29135 19670 29144
rect 19524 29106 19576 29112
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 19628 28490 19656 28698
rect 19720 28558 19748 30280
rect 19800 30262 19852 30268
rect 19800 30048 19852 30054
rect 19800 29990 19852 29996
rect 19812 29646 19840 29990
rect 19904 29850 19932 30330
rect 19892 29844 19944 29850
rect 19892 29786 19944 29792
rect 19800 29640 19852 29646
rect 19800 29582 19852 29588
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19996 29238 20024 29446
rect 19984 29232 20036 29238
rect 19984 29174 20036 29180
rect 20364 28762 20392 34734
rect 20444 34740 20496 34746
rect 20444 34682 20496 34688
rect 20444 34536 20496 34542
rect 20444 34478 20496 34484
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20456 28642 20484 34478
rect 20640 33402 20668 36178
rect 21192 36174 21220 36722
rect 21180 36168 21232 36174
rect 21180 36110 21232 36116
rect 20811 35932 21119 35952
rect 20811 35930 20817 35932
rect 20873 35930 20897 35932
rect 20953 35930 20977 35932
rect 21033 35930 21057 35932
rect 21113 35930 21119 35932
rect 20873 35878 20875 35930
rect 21055 35878 21057 35930
rect 20811 35876 20817 35878
rect 20873 35876 20897 35878
rect 20953 35876 20977 35878
rect 21033 35876 21057 35878
rect 21113 35876 21119 35878
rect 20811 35856 21119 35876
rect 20812 35624 20864 35630
rect 20812 35566 20864 35572
rect 20824 35290 20852 35566
rect 20812 35284 20864 35290
rect 20812 35226 20864 35232
rect 21192 35086 21220 36110
rect 21284 35698 21312 37198
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 21180 35080 21232 35086
rect 21180 35022 21232 35028
rect 20811 34844 21119 34864
rect 20811 34842 20817 34844
rect 20873 34842 20897 34844
rect 20953 34842 20977 34844
rect 21033 34842 21057 34844
rect 21113 34842 21119 34844
rect 20873 34790 20875 34842
rect 21055 34790 21057 34842
rect 20811 34788 20817 34790
rect 20873 34788 20897 34790
rect 20953 34788 20977 34790
rect 21033 34788 21057 34790
rect 21113 34788 21119 34790
rect 20811 34768 21119 34788
rect 20811 33756 21119 33776
rect 20811 33754 20817 33756
rect 20873 33754 20897 33756
rect 20953 33754 20977 33756
rect 21033 33754 21057 33756
rect 21113 33754 21119 33756
rect 20873 33702 20875 33754
rect 21055 33702 21057 33754
rect 20811 33700 20817 33702
rect 20873 33700 20897 33702
rect 20953 33700 20977 33702
rect 21033 33700 21057 33702
rect 21113 33700 21119 33702
rect 20811 33680 21119 33700
rect 20548 33374 20668 33402
rect 20548 33046 20576 33374
rect 20628 33312 20680 33318
rect 20628 33254 20680 33260
rect 20536 33040 20588 33046
rect 20536 32982 20588 32988
rect 20536 32904 20588 32910
rect 20536 32846 20588 32852
rect 20548 32570 20576 32846
rect 20536 32564 20588 32570
rect 20536 32506 20588 32512
rect 20640 30666 20668 33254
rect 21284 32910 21312 35634
rect 21376 35562 21404 41074
rect 21468 40118 21496 41228
rect 21560 41018 21588 48470
rect 21744 48362 21772 48583
rect 21652 48334 21772 48362
rect 21652 41138 21680 48334
rect 21732 48136 21784 48142
rect 21732 48078 21784 48084
rect 21640 41132 21692 41138
rect 21640 41074 21692 41080
rect 21560 40990 21680 41018
rect 21744 41002 21772 48078
rect 21836 41818 21864 53042
rect 21916 52964 21968 52970
rect 21916 52906 21968 52912
rect 21928 52562 21956 52906
rect 21916 52556 21968 52562
rect 21916 52498 21968 52504
rect 22020 50969 22048 53094
rect 22100 53100 22152 53106
rect 22100 53042 22152 53048
rect 22112 50998 22140 53042
rect 22192 52420 22244 52426
rect 22192 52362 22244 52368
rect 22204 51610 22232 52362
rect 22192 51604 22244 51610
rect 22192 51546 22244 51552
rect 22100 50992 22152 50998
rect 22006 50960 22062 50969
rect 22100 50934 22152 50940
rect 22296 50930 22324 54470
rect 22376 53576 22428 53582
rect 22376 53518 22428 53524
rect 22388 53106 22416 53518
rect 22572 53514 22600 54862
rect 22664 54806 22692 60726
rect 22848 60722 22876 61542
rect 22836 60716 22888 60722
rect 22836 60658 22888 60664
rect 22744 56704 22796 56710
rect 22744 56646 22796 56652
rect 22756 56438 22784 56646
rect 22744 56432 22796 56438
rect 22744 56374 22796 56380
rect 22744 55616 22796 55622
rect 22744 55558 22796 55564
rect 22652 54800 22704 54806
rect 22652 54742 22704 54748
rect 22560 53508 22612 53514
rect 22560 53450 22612 53456
rect 22468 53440 22520 53446
rect 22468 53382 22520 53388
rect 22376 53100 22428 53106
rect 22376 53042 22428 53048
rect 22480 52154 22508 53382
rect 22468 52148 22520 52154
rect 22468 52090 22520 52096
rect 22560 51944 22612 51950
rect 22560 51886 22612 51892
rect 22468 51400 22520 51406
rect 22468 51342 22520 51348
rect 22480 51066 22508 51342
rect 22376 51060 22428 51066
rect 22376 51002 22428 51008
rect 22468 51060 22520 51066
rect 22468 51002 22520 51008
rect 22006 50895 22062 50904
rect 22284 50924 22336 50930
rect 22284 50866 22336 50872
rect 22192 50856 22244 50862
rect 22192 50798 22244 50804
rect 21916 50788 21968 50794
rect 21916 50730 21968 50736
rect 22008 50788 22060 50794
rect 22008 50730 22060 50736
rect 21928 49609 21956 50730
rect 22020 49706 22048 50730
rect 22100 50720 22152 50726
rect 22100 50662 22152 50668
rect 22008 49700 22060 49706
rect 22008 49642 22060 49648
rect 21914 49600 21970 49609
rect 21914 49535 21970 49544
rect 22112 48754 22140 50662
rect 22204 49212 22232 50798
rect 22388 50522 22416 51002
rect 22376 50516 22428 50522
rect 22376 50458 22428 50464
rect 22468 50312 22520 50318
rect 22468 50254 22520 50260
rect 22376 49836 22428 49842
rect 22376 49778 22428 49784
rect 22388 49434 22416 49778
rect 22376 49428 22428 49434
rect 22376 49370 22428 49376
rect 22284 49224 22336 49230
rect 22204 49184 22284 49212
rect 22100 48748 22152 48754
rect 22100 48690 22152 48696
rect 22100 48544 22152 48550
rect 22100 48486 22152 48492
rect 21916 46028 21968 46034
rect 21916 45970 21968 45976
rect 21928 45554 21956 45970
rect 22112 45558 22140 48486
rect 22204 46481 22232 49184
rect 22284 49166 22336 49172
rect 22480 49162 22508 50254
rect 22468 49156 22520 49162
rect 22468 49098 22520 49104
rect 22376 48816 22428 48822
rect 22376 48758 22428 48764
rect 22388 48124 22416 48758
rect 22480 48278 22508 49098
rect 22468 48272 22520 48278
rect 22468 48214 22520 48220
rect 22388 48096 22508 48124
rect 22284 47048 22336 47054
rect 22284 46990 22336 46996
rect 22190 46472 22246 46481
rect 22190 46407 22246 46416
rect 22192 46368 22244 46374
rect 22192 46310 22244 46316
rect 22204 45966 22232 46310
rect 22296 46170 22324 46990
rect 22376 46912 22428 46918
rect 22376 46854 22428 46860
rect 22388 46578 22416 46854
rect 22376 46572 22428 46578
rect 22376 46514 22428 46520
rect 22480 46510 22508 48096
rect 22572 47190 22600 51886
rect 22652 51400 22704 51406
rect 22652 51342 22704 51348
rect 22664 50289 22692 51342
rect 22756 50726 22784 55558
rect 22834 55312 22890 55321
rect 22834 55247 22890 55256
rect 22848 54262 22876 55247
rect 22836 54256 22888 54262
rect 22836 54198 22888 54204
rect 22940 52018 22968 63922
rect 23032 59566 23060 66166
rect 23308 66162 23336 66710
rect 23584 66638 23612 66778
rect 23572 66632 23624 66638
rect 23572 66574 23624 66580
rect 23388 66496 23440 66502
rect 23388 66438 23440 66444
rect 23296 66156 23348 66162
rect 23296 66098 23348 66104
rect 23204 65204 23256 65210
rect 23204 65146 23256 65152
rect 23216 63986 23244 65146
rect 23400 64870 23428 66438
rect 23584 66162 23612 66574
rect 23664 66496 23716 66502
rect 23664 66438 23716 66444
rect 23572 66156 23624 66162
rect 23572 66098 23624 66104
rect 23480 65952 23532 65958
rect 23480 65894 23532 65900
rect 23492 65006 23520 65894
rect 23480 65000 23532 65006
rect 23480 64942 23532 64948
rect 23388 64864 23440 64870
rect 23388 64806 23440 64812
rect 23480 64456 23532 64462
rect 23480 64398 23532 64404
rect 23492 63986 23520 64398
rect 23204 63980 23256 63986
rect 23204 63922 23256 63928
rect 23480 63980 23532 63986
rect 23480 63922 23532 63928
rect 23388 63572 23440 63578
rect 23388 63514 23440 63520
rect 23112 60716 23164 60722
rect 23112 60658 23164 60664
rect 23124 60058 23152 60658
rect 23204 60104 23256 60110
rect 23124 60052 23204 60058
rect 23124 60046 23256 60052
rect 23124 60030 23244 60046
rect 23124 59634 23152 60030
rect 23296 59968 23348 59974
rect 23296 59910 23348 59916
rect 23112 59628 23164 59634
rect 23112 59570 23164 59576
rect 23020 59560 23072 59566
rect 23020 59502 23072 59508
rect 23020 57996 23072 58002
rect 23020 57938 23072 57944
rect 23032 57338 23060 57938
rect 23124 57458 23152 59570
rect 23204 59424 23256 59430
rect 23204 59366 23256 59372
rect 23112 57452 23164 57458
rect 23112 57394 23164 57400
rect 23032 57310 23152 57338
rect 23020 57248 23072 57254
rect 23020 57190 23072 57196
rect 23032 56846 23060 57190
rect 23020 56840 23072 56846
rect 23020 56782 23072 56788
rect 23020 56500 23072 56506
rect 23020 56442 23072 56448
rect 23032 52358 23060 56442
rect 23124 55758 23152 57310
rect 23112 55752 23164 55758
rect 23112 55694 23164 55700
rect 23112 55412 23164 55418
rect 23112 55354 23164 55360
rect 23124 53650 23152 55354
rect 23216 55321 23244 59366
rect 23308 56545 23336 59910
rect 23400 59226 23428 63514
rect 23492 62286 23520 63922
rect 23584 63510 23612 66098
rect 23676 63578 23704 66438
rect 23756 65000 23808 65006
rect 23756 64942 23808 64948
rect 23664 63572 23716 63578
rect 23664 63514 23716 63520
rect 23572 63504 23624 63510
rect 23572 63446 23624 63452
rect 23664 63436 23716 63442
rect 23664 63378 23716 63384
rect 23480 62280 23532 62286
rect 23480 62222 23532 62228
rect 23492 61606 23520 62222
rect 23480 61600 23532 61606
rect 23480 61542 23532 61548
rect 23492 61198 23520 61542
rect 23480 61192 23532 61198
rect 23480 61134 23532 61140
rect 23480 61056 23532 61062
rect 23480 60998 23532 61004
rect 23492 60246 23520 60998
rect 23572 60512 23624 60518
rect 23572 60454 23624 60460
rect 23480 60240 23532 60246
rect 23480 60182 23532 60188
rect 23480 59560 23532 59566
rect 23480 59502 23532 59508
rect 23388 59220 23440 59226
rect 23388 59162 23440 59168
rect 23492 57089 23520 59502
rect 23478 57080 23534 57089
rect 23478 57015 23534 57024
rect 23480 56976 23532 56982
rect 23480 56918 23532 56924
rect 23388 56772 23440 56778
rect 23388 56714 23440 56720
rect 23294 56536 23350 56545
rect 23294 56471 23350 56480
rect 23296 56364 23348 56370
rect 23296 56306 23348 56312
rect 23202 55312 23258 55321
rect 23308 55282 23336 56306
rect 23202 55247 23258 55256
rect 23296 55276 23348 55282
rect 23296 55218 23348 55224
rect 23204 55208 23256 55214
rect 23202 55176 23204 55185
rect 23256 55176 23258 55185
rect 23202 55111 23258 55120
rect 23204 55072 23256 55078
rect 23204 55014 23256 55020
rect 23112 53644 23164 53650
rect 23112 53586 23164 53592
rect 23112 53508 23164 53514
rect 23112 53450 23164 53456
rect 23020 52352 23072 52358
rect 23020 52294 23072 52300
rect 23020 52148 23072 52154
rect 23020 52090 23072 52096
rect 22928 52012 22980 52018
rect 22928 51954 22980 51960
rect 22836 51400 22888 51406
rect 22836 51342 22888 51348
rect 22744 50720 22796 50726
rect 22744 50662 22796 50668
rect 22650 50280 22706 50289
rect 22650 50215 22706 50224
rect 22652 50176 22704 50182
rect 22848 50130 22876 51342
rect 22652 50118 22704 50124
rect 22560 47184 22612 47190
rect 22560 47126 22612 47132
rect 22560 47048 22612 47054
rect 22560 46990 22612 46996
rect 22468 46504 22520 46510
rect 22468 46446 22520 46452
rect 22284 46164 22336 46170
rect 22284 46106 22336 46112
rect 22480 46034 22508 46446
rect 22468 46028 22520 46034
rect 22468 45970 22520 45976
rect 22192 45960 22244 45966
rect 22192 45902 22244 45908
rect 22572 45880 22600 46990
rect 22480 45852 22600 45880
rect 21928 45526 22048 45554
rect 21916 45484 21968 45490
rect 21916 45426 21968 45432
rect 21928 42770 21956 45426
rect 22020 43790 22048 45526
rect 22100 45552 22152 45558
rect 22100 45494 22152 45500
rect 22480 45490 22508 45852
rect 22664 45778 22692 50118
rect 22756 50102 22876 50130
rect 22756 47054 22784 50102
rect 22834 50008 22890 50017
rect 22834 49943 22890 49952
rect 22744 47048 22796 47054
rect 22744 46990 22796 46996
rect 22744 46572 22796 46578
rect 22744 46514 22796 46520
rect 22572 45750 22692 45778
rect 22468 45484 22520 45490
rect 22468 45426 22520 45432
rect 22468 45280 22520 45286
rect 22468 45222 22520 45228
rect 22284 45076 22336 45082
rect 22284 45018 22336 45024
rect 22008 43784 22060 43790
rect 22008 43726 22060 43732
rect 22192 43648 22244 43654
rect 22192 43590 22244 43596
rect 22006 43344 22062 43353
rect 22006 43279 22062 43288
rect 21916 42764 21968 42770
rect 21916 42706 21968 42712
rect 21824 41812 21876 41818
rect 21824 41754 21876 41760
rect 21928 41274 21956 42706
rect 22020 41818 22048 43279
rect 22204 42294 22232 43590
rect 22296 42702 22324 45018
rect 22376 44804 22428 44810
rect 22376 44746 22428 44752
rect 22388 43194 22416 44746
rect 22480 43790 22508 45222
rect 22468 43784 22520 43790
rect 22468 43726 22520 43732
rect 22388 43166 22508 43194
rect 22376 43104 22428 43110
rect 22376 43046 22428 43052
rect 22284 42696 22336 42702
rect 22284 42638 22336 42644
rect 22284 42560 22336 42566
rect 22282 42528 22284 42537
rect 22336 42528 22338 42537
rect 22282 42463 22338 42472
rect 22100 42288 22152 42294
rect 22100 42230 22152 42236
rect 22192 42288 22244 42294
rect 22192 42230 22244 42236
rect 22112 41834 22140 42230
rect 22008 41812 22060 41818
rect 22112 41806 22232 41834
rect 22008 41754 22060 41760
rect 22204 41750 22232 41806
rect 22100 41744 22152 41750
rect 22098 41712 22100 41721
rect 22192 41744 22244 41750
rect 22152 41712 22154 41721
rect 22192 41686 22244 41692
rect 22098 41647 22154 41656
rect 21916 41268 21968 41274
rect 21916 41210 21968 41216
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 22020 41154 22048 41210
rect 21928 41126 22048 41154
rect 22284 41200 22336 41206
rect 22284 41142 22336 41148
rect 21548 40928 21600 40934
rect 21548 40870 21600 40876
rect 21456 40112 21508 40118
rect 21456 40054 21508 40060
rect 21468 39914 21496 40054
rect 21456 39908 21508 39914
rect 21456 39850 21508 39856
rect 21560 38350 21588 40870
rect 21652 40118 21680 40990
rect 21732 40996 21784 41002
rect 21732 40938 21784 40944
rect 21640 40112 21692 40118
rect 21640 40054 21692 40060
rect 21548 38344 21600 38350
rect 21548 38286 21600 38292
rect 21456 36236 21508 36242
rect 21652 36224 21680 40054
rect 21824 39840 21876 39846
rect 21824 39782 21876 39788
rect 21730 38312 21786 38321
rect 21730 38247 21786 38256
rect 21744 37942 21772 38247
rect 21732 37936 21784 37942
rect 21732 37878 21784 37884
rect 21732 37188 21784 37194
rect 21732 37130 21784 37136
rect 21744 36718 21772 37130
rect 21836 37126 21864 39782
rect 21928 37398 21956 41126
rect 22008 40996 22060 41002
rect 22008 40938 22060 40944
rect 21916 37392 21968 37398
rect 21916 37334 21968 37340
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21824 37120 21876 37126
rect 21824 37062 21876 37068
rect 21928 36718 21956 37198
rect 22020 37126 22048 40938
rect 22296 40526 22324 41142
rect 22100 40520 22152 40526
rect 22100 40462 22152 40468
rect 22284 40520 22336 40526
rect 22284 40462 22336 40468
rect 22112 40225 22140 40462
rect 22098 40216 22154 40225
rect 22098 40151 22154 40160
rect 22100 39908 22152 39914
rect 22100 39850 22152 39856
rect 22008 37120 22060 37126
rect 22008 37062 22060 37068
rect 22020 36786 22048 37062
rect 22112 36786 22140 39850
rect 22284 39296 22336 39302
rect 22284 39238 22336 39244
rect 22192 38480 22244 38486
rect 22192 38422 22244 38428
rect 22204 38185 22232 38422
rect 22190 38176 22246 38185
rect 22190 38111 22246 38120
rect 22296 37262 22324 39238
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22008 36780 22060 36786
rect 22008 36722 22060 36728
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 21916 36712 21968 36718
rect 21916 36654 21968 36660
rect 21824 36576 21876 36582
rect 21824 36518 21876 36524
rect 21508 36196 21680 36224
rect 21456 36178 21508 36184
rect 21364 35556 21416 35562
rect 21364 35498 21416 35504
rect 21272 32904 21324 32910
rect 21270 32872 21272 32881
rect 21324 32872 21326 32881
rect 21270 32807 21326 32816
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20732 31822 20760 32710
rect 20811 32668 21119 32688
rect 20811 32666 20817 32668
rect 20873 32666 20897 32668
rect 20953 32666 20977 32668
rect 21033 32666 21057 32668
rect 21113 32666 21119 32668
rect 20873 32614 20875 32666
rect 21055 32614 21057 32666
rect 20811 32612 20817 32614
rect 20873 32612 20897 32614
rect 20953 32612 20977 32614
rect 21033 32612 21057 32614
rect 21113 32612 21119 32614
rect 20811 32592 21119 32612
rect 21284 31822 21312 32807
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 21272 31816 21324 31822
rect 21272 31758 21324 31764
rect 20811 31580 21119 31600
rect 20811 31578 20817 31580
rect 20873 31578 20897 31580
rect 20953 31578 20977 31580
rect 21033 31578 21057 31580
rect 21113 31578 21119 31580
rect 20873 31526 20875 31578
rect 21055 31526 21057 31578
rect 20811 31524 20817 31526
rect 20873 31524 20897 31526
rect 20953 31524 20977 31526
rect 21033 31524 21057 31526
rect 21113 31524 21119 31526
rect 20811 31504 21119 31524
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20720 30660 20772 30666
rect 20720 30602 20772 30608
rect 20732 29714 20760 30602
rect 20811 30492 21119 30512
rect 20811 30490 20817 30492
rect 20873 30490 20897 30492
rect 20953 30490 20977 30492
rect 21033 30490 21057 30492
rect 21113 30490 21119 30492
rect 20873 30438 20875 30490
rect 21055 30438 21057 30490
rect 20811 30436 20817 30438
rect 20873 30436 20897 30438
rect 20953 30436 20977 30438
rect 21033 30436 21057 30438
rect 21113 30436 21119 30438
rect 20811 30416 21119 30436
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 20811 29404 21119 29424
rect 20811 29402 20817 29404
rect 20873 29402 20897 29404
rect 20953 29402 20977 29404
rect 21033 29402 21057 29404
rect 21113 29402 21119 29404
rect 20873 29350 20875 29402
rect 21055 29350 21057 29402
rect 20811 29348 20817 29350
rect 20873 29348 20897 29350
rect 20953 29348 20977 29350
rect 21033 29348 21057 29350
rect 21113 29348 21119 29350
rect 20811 29328 21119 29348
rect 20996 29232 21048 29238
rect 20996 29174 21048 29180
rect 20088 28626 20484 28642
rect 20536 28688 20588 28694
rect 20536 28630 20588 28636
rect 20076 28620 20484 28626
rect 20128 28614 20484 28620
rect 20076 28562 20128 28568
rect 19708 28552 19760 28558
rect 19708 28494 19760 28500
rect 19616 28484 19668 28490
rect 19616 28426 19668 28432
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19536 28082 19564 28358
rect 19628 28098 19656 28426
rect 19524 28076 19576 28082
rect 19628 28070 19840 28098
rect 19524 28018 19576 28024
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 19628 25362 19656 25638
rect 19616 25356 19668 25362
rect 19616 25298 19668 25304
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19260 24410 19288 24754
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19536 24206 19564 24550
rect 19812 24206 19840 28070
rect 20088 27044 20116 28426
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20180 28150 20208 28358
rect 20168 28144 20220 28150
rect 20168 28086 20220 28092
rect 20088 27016 20208 27044
rect 20180 26790 20208 27016
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20180 25974 20208 26726
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 18524 22094 18552 23666
rect 18524 22066 18644 22094
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18420 21548 18472 21554
rect 18420 21490 18472 21496
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18064 21010 18092 21286
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 18064 20466 18092 20810
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 18064 20330 18092 20402
rect 18052 20324 18104 20330
rect 18052 20266 18104 20272
rect 18156 20210 18184 21422
rect 18524 21350 18552 21966
rect 18616 21554 18644 22066
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19260 21554 19288 21830
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18064 20182 18184 20210
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18064 19310 18092 20182
rect 18248 19854 18276 20198
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18248 19378 18276 19790
rect 18616 19378 18644 21490
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20942 19380 21286
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19260 19854 19288 20402
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19260 19446 19288 19790
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18064 17338 18092 19246
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18616 17202 18644 17546
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18248 16250 18460 16266
rect 18236 16244 18472 16250
rect 18288 16238 18420 16244
rect 18236 16186 18288 16192
rect 18420 16186 18472 16192
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17914 16176 17966 16182
rect 17966 16136 18184 16164
rect 17914 16118 17966 16124
rect 18156 16130 18184 16136
rect 18156 16102 18368 16130
rect 18340 16046 18368 16102
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18052 15904 18104 15910
rect 18142 15872 18198 15881
rect 18104 15852 18142 15858
rect 18052 15846 18142 15852
rect 18064 15830 18142 15846
rect 18142 15807 18198 15816
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18432 14618 18460 15370
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18524 12238 18552 16934
rect 18708 16726 18736 17002
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18616 15978 18644 16526
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18708 16425 18736 16458
rect 18694 16416 18750 16425
rect 18694 16351 18750 16360
rect 18604 15972 18656 15978
rect 18604 15914 18656 15920
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17512 10674 17540 12038
rect 17880 11762 17908 12038
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17972 10198 18000 10678
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 18800 6914 18828 18022
rect 18984 17610 19012 19246
rect 19352 18834 19380 19994
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19536 18086 19564 24142
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 19628 21554 19656 24074
rect 19708 23520 19760 23526
rect 19708 23462 19760 23468
rect 19720 23186 19748 23462
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19246 16824 19302 16833
rect 18972 16788 19024 16794
rect 19246 16759 19248 16768
rect 18972 16730 19024 16736
rect 19300 16759 19302 16768
rect 19248 16730 19300 16736
rect 18880 16720 18932 16726
rect 18878 16688 18880 16697
rect 18932 16688 18934 16697
rect 18878 16623 18934 16632
rect 18984 16574 19012 16730
rect 18878 16552 18934 16561
rect 18984 16546 19288 16574
rect 18878 16487 18880 16496
rect 18932 16487 18934 16496
rect 18880 16458 18932 16464
rect 19260 15502 19288 16546
rect 19352 16454 19380 17070
rect 19444 16726 19472 17682
rect 19628 17678 19656 19314
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19524 17196 19576 17202
rect 19628 17184 19656 17614
rect 19708 17536 19760 17542
rect 19760 17496 19840 17524
rect 19708 17478 19760 17484
rect 19576 17156 19748 17184
rect 19524 17138 19576 17144
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19536 16674 19564 16934
rect 19536 16646 19565 16674
rect 19537 16574 19565 16646
rect 19720 16590 19748 17156
rect 19536 16561 19565 16574
rect 19708 16584 19760 16590
rect 19522 16552 19578 16561
rect 19708 16526 19760 16532
rect 19522 16487 19578 16496
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19352 16266 19380 16390
rect 19352 16238 19656 16266
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19352 15638 19380 16050
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19352 15026 19380 15574
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19444 14414 19472 14894
rect 19524 14544 19576 14550
rect 19522 14512 19524 14521
rect 19576 14512 19578 14521
rect 19522 14447 19578 14456
rect 19628 14414 19656 16238
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19720 15502 19748 15846
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19812 15094 19840 17496
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19904 16794 19932 17138
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19890 16688 19946 16697
rect 19890 16623 19892 16632
rect 19944 16623 19946 16632
rect 19892 16594 19944 16600
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 19892 16448 19944 16454
rect 19890 16416 19892 16425
rect 19944 16416 19946 16425
rect 19890 16351 19946 16360
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 20088 14958 20116 16526
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19996 14414 20024 14758
rect 20088 14618 20116 14894
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 13190 19564 14214
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19352 11898 19380 13126
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11354 19288 11698
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19352 10606 19380 11834
rect 19628 11694 19656 14350
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19996 11762 20024 11834
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19616 11280 19668 11286
rect 19614 11248 19616 11257
rect 19668 11248 19670 11257
rect 19614 11183 19670 11192
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10674 19472 11086
rect 19720 10742 19748 11494
rect 19812 11082 19840 11630
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 20088 9568 20116 14554
rect 20180 14414 20208 15438
rect 20272 14482 20300 28614
rect 20548 28218 20576 28630
rect 21008 28558 21036 29174
rect 21180 28960 21232 28966
rect 21180 28902 21232 28908
rect 21192 28558 21220 28902
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21284 28422 21312 31758
rect 21468 30870 21496 36178
rect 21836 36106 21864 36518
rect 21824 36100 21876 36106
rect 21824 36042 21876 36048
rect 21928 36038 21956 36654
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 21916 36032 21968 36038
rect 21916 35974 21968 35980
rect 21824 34944 21876 34950
rect 21824 34886 21876 34892
rect 21732 34400 21784 34406
rect 21732 34342 21784 34348
rect 21456 30864 21508 30870
rect 21456 30806 21508 30812
rect 21364 29572 21416 29578
rect 21364 29514 21416 29520
rect 21272 28416 21324 28422
rect 21272 28358 21324 28364
rect 20811 28316 21119 28336
rect 20811 28314 20817 28316
rect 20873 28314 20897 28316
rect 20953 28314 20977 28316
rect 21033 28314 21057 28316
rect 21113 28314 21119 28316
rect 20873 28262 20875 28314
rect 21055 28262 21057 28314
rect 20811 28260 20817 28262
rect 20873 28260 20897 28262
rect 20953 28260 20977 28262
rect 21033 28260 21057 28262
rect 21113 28260 21119 28262
rect 20811 28240 21119 28260
rect 20536 28212 20588 28218
rect 20536 28154 20588 28160
rect 20811 27228 21119 27248
rect 20811 27226 20817 27228
rect 20873 27226 20897 27228
rect 20953 27226 20977 27228
rect 21033 27226 21057 27228
rect 21113 27226 21119 27228
rect 20873 27174 20875 27226
rect 21055 27174 21057 27226
rect 20811 27172 20817 27174
rect 20873 27172 20897 27174
rect 20953 27172 20977 27174
rect 21033 27172 21057 27174
rect 21113 27172 21119 27174
rect 20811 27152 21119 27172
rect 20811 26140 21119 26160
rect 20811 26138 20817 26140
rect 20873 26138 20897 26140
rect 20953 26138 20977 26140
rect 21033 26138 21057 26140
rect 21113 26138 21119 26140
rect 20873 26086 20875 26138
rect 21055 26086 21057 26138
rect 20811 26084 20817 26086
rect 20873 26084 20897 26086
rect 20953 26084 20977 26086
rect 21033 26084 21057 26086
rect 21113 26084 21119 26086
rect 20811 26064 21119 26084
rect 20628 25220 20680 25226
rect 20628 25162 20680 25168
rect 20640 24954 20668 25162
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 20811 25052 21119 25072
rect 20811 25050 20817 25052
rect 20873 25050 20897 25052
rect 20953 25050 20977 25052
rect 21033 25050 21057 25052
rect 21113 25050 21119 25052
rect 20873 24998 20875 25050
rect 21055 24998 21057 25050
rect 20811 24996 20817 24998
rect 20873 24996 20897 24998
rect 20953 24996 20977 24998
rect 21033 24996 21057 24998
rect 21113 24996 21119 24998
rect 20811 24976 21119 24996
rect 20628 24948 20680 24954
rect 20628 24890 20680 24896
rect 21284 24818 21312 25094
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21376 24682 21404 29514
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21560 29170 21588 29446
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 21548 29164 21600 29170
rect 21548 29106 21600 29112
rect 21560 28422 21588 29106
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 21560 27674 21588 28358
rect 21548 27668 21600 27674
rect 21548 27610 21600 27616
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 21468 25786 21496 27338
rect 21560 26874 21588 27610
rect 21652 27470 21680 29174
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21560 26846 21680 26874
rect 21468 25758 21588 25786
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21364 24676 21416 24682
rect 21364 24618 21416 24624
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21088 24200 21140 24206
rect 21140 24148 21220 24154
rect 21088 24142 21220 24148
rect 21100 24126 21220 24142
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20732 23050 20760 24006
rect 20811 23964 21119 23984
rect 20811 23962 20817 23964
rect 20873 23962 20897 23964
rect 20953 23962 20977 23964
rect 21033 23962 21057 23964
rect 21113 23962 21119 23964
rect 20873 23910 20875 23962
rect 21055 23910 21057 23962
rect 20811 23908 20817 23910
rect 20873 23908 20897 23910
rect 20953 23908 20977 23910
rect 21033 23908 21057 23910
rect 21113 23908 21119 23910
rect 20811 23888 21119 23908
rect 21192 23730 21220 24126
rect 21284 23730 21312 24550
rect 21376 24138 21404 24618
rect 21468 24206 21496 25638
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21192 23186 21220 23666
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20811 22876 21119 22896
rect 20811 22874 20817 22876
rect 20873 22874 20897 22876
rect 20953 22874 20977 22876
rect 21033 22874 21057 22876
rect 21113 22874 21119 22876
rect 20873 22822 20875 22874
rect 21055 22822 21057 22874
rect 20811 22820 20817 22822
rect 20873 22820 20897 22822
rect 20953 22820 20977 22822
rect 21033 22820 21057 22822
rect 21113 22820 21119 22822
rect 20811 22800 21119 22820
rect 21192 22642 21220 23122
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21284 22522 21312 23666
rect 21560 23118 21588 25758
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21652 22642 21680 26846
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 21364 22568 21416 22574
rect 21284 22516 21364 22522
rect 21284 22510 21416 22516
rect 21284 22494 21404 22510
rect 21284 22438 21312 22494
rect 21272 22432 21324 22438
rect 21272 22374 21324 22380
rect 20811 21788 21119 21808
rect 20811 21786 20817 21788
rect 20873 21786 20897 21788
rect 20953 21786 20977 21788
rect 21033 21786 21057 21788
rect 21113 21786 21119 21788
rect 20873 21734 20875 21786
rect 21055 21734 21057 21786
rect 20811 21732 20817 21734
rect 20873 21732 20897 21734
rect 20953 21732 20977 21734
rect 21033 21732 21057 21734
rect 21113 21732 21119 21734
rect 20811 21712 21119 21732
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20640 20534 20668 20742
rect 20811 20700 21119 20720
rect 20811 20698 20817 20700
rect 20873 20698 20897 20700
rect 20953 20698 20977 20700
rect 21033 20698 21057 20700
rect 21113 20698 21119 20700
rect 20873 20646 20875 20698
rect 21055 20646 21057 20698
rect 20811 20644 20817 20646
rect 20873 20644 20897 20646
rect 20953 20644 20977 20646
rect 21033 20644 21057 20646
rect 21113 20644 21119 20646
rect 20811 20624 21119 20644
rect 20628 20528 20680 20534
rect 20628 20470 20680 20476
rect 20640 19854 20668 20470
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20732 18290 20760 19654
rect 20811 19612 21119 19632
rect 20811 19610 20817 19612
rect 20873 19610 20897 19612
rect 20953 19610 20977 19612
rect 21033 19610 21057 19612
rect 21113 19610 21119 19612
rect 20873 19558 20875 19610
rect 21055 19558 21057 19610
rect 20811 19556 20817 19558
rect 20873 19556 20897 19558
rect 20953 19556 20977 19558
rect 21033 19556 21057 19558
rect 21113 19556 21119 19558
rect 20811 19536 21119 19556
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 20811 18524 21119 18544
rect 20811 18522 20817 18524
rect 20873 18522 20897 18524
rect 20953 18522 20977 18524
rect 21033 18522 21057 18524
rect 21113 18522 21119 18524
rect 20873 18470 20875 18522
rect 21055 18470 21057 18522
rect 20811 18468 20817 18470
rect 20873 18468 20897 18470
rect 20953 18468 20977 18470
rect 21033 18468 21057 18470
rect 21113 18468 21119 18470
rect 20811 18448 21119 18468
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20364 17134 20392 17614
rect 20811 17436 21119 17456
rect 20811 17434 20817 17436
rect 20873 17434 20897 17436
rect 20953 17434 20977 17436
rect 21033 17434 21057 17436
rect 21113 17434 21119 17436
rect 20873 17382 20875 17434
rect 21055 17382 21057 17434
rect 20811 17380 20817 17382
rect 20873 17380 20897 17382
rect 20953 17380 20977 17382
rect 21033 17380 21057 17382
rect 21113 17380 21119 17382
rect 20811 17360 21119 17380
rect 21284 17202 21312 19314
rect 21468 17678 21496 19722
rect 21744 18630 21772 34342
rect 21836 32552 21864 34886
rect 21928 32978 21956 35974
rect 22112 35630 22140 36110
rect 22296 36106 22324 37198
rect 22284 36100 22336 36106
rect 22284 36042 22336 36048
rect 22388 35698 22416 43046
rect 22480 41274 22508 43166
rect 22468 41268 22520 41274
rect 22468 41210 22520 41216
rect 22468 41132 22520 41138
rect 22468 41074 22520 41080
rect 22480 40662 22508 41074
rect 22468 40656 22520 40662
rect 22468 40598 22520 40604
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22480 40050 22508 40462
rect 22468 40044 22520 40050
rect 22468 39986 22520 39992
rect 22572 36582 22600 45750
rect 22652 45552 22704 45558
rect 22652 45494 22704 45500
rect 22664 44878 22692 45494
rect 22652 44872 22704 44878
rect 22652 44814 22704 44820
rect 22652 44736 22704 44742
rect 22652 44678 22704 44684
rect 22664 42566 22692 44678
rect 22756 44402 22784 46514
rect 22848 46170 22876 49943
rect 22940 49094 22968 51954
rect 23032 50454 23060 52090
rect 23020 50448 23072 50454
rect 23020 50390 23072 50396
rect 23020 50312 23072 50318
rect 23020 50254 23072 50260
rect 23032 49978 23060 50254
rect 23020 49972 23072 49978
rect 23020 49914 23072 49920
rect 23018 49872 23074 49881
rect 23018 49807 23074 49816
rect 22928 49088 22980 49094
rect 22928 49030 22980 49036
rect 22940 48890 22968 49030
rect 22928 48884 22980 48890
rect 22928 48826 22980 48832
rect 22928 48612 22980 48618
rect 22928 48554 22980 48560
rect 22940 46578 22968 48554
rect 23032 48550 23060 49807
rect 23020 48544 23072 48550
rect 23020 48486 23072 48492
rect 23124 47054 23152 53450
rect 23112 47048 23164 47054
rect 23112 46990 23164 46996
rect 23020 46912 23072 46918
rect 23020 46854 23072 46860
rect 22928 46572 22980 46578
rect 22928 46514 22980 46520
rect 23032 46458 23060 46854
rect 23124 46578 23152 46990
rect 23112 46572 23164 46578
rect 23112 46514 23164 46520
rect 22940 46430 23060 46458
rect 23112 46436 23164 46442
rect 22836 46164 22888 46170
rect 22836 46106 22888 46112
rect 22836 46028 22888 46034
rect 22836 45970 22888 45976
rect 22744 44396 22796 44402
rect 22744 44338 22796 44344
rect 22652 42560 22704 42566
rect 22652 42502 22704 42508
rect 22756 41256 22784 44338
rect 22664 41228 22784 41256
rect 22664 40118 22692 41228
rect 22744 41132 22796 41138
rect 22744 41074 22796 41080
rect 22756 40186 22784 41074
rect 22744 40180 22796 40186
rect 22744 40122 22796 40128
rect 22652 40112 22704 40118
rect 22652 40054 22704 40060
rect 22664 39370 22692 40054
rect 22744 40044 22796 40050
rect 22744 39986 22796 39992
rect 22652 39364 22704 39370
rect 22652 39306 22704 39312
rect 22664 39098 22692 39306
rect 22652 39092 22704 39098
rect 22652 39034 22704 39040
rect 22664 38010 22692 39034
rect 22756 38758 22784 39986
rect 22744 38752 22796 38758
rect 22744 38694 22796 38700
rect 22652 38004 22704 38010
rect 22652 37946 22704 37952
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 22664 36224 22692 36654
rect 22480 36196 22692 36224
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22100 35624 22152 35630
rect 22100 35566 22152 35572
rect 22284 35624 22336 35630
rect 22284 35566 22336 35572
rect 22112 35086 22140 35566
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 21916 32972 21968 32978
rect 21916 32914 21968 32920
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21836 32524 21956 32552
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21836 31482 21864 32370
rect 21928 31958 21956 32524
rect 22020 32450 22048 32710
rect 22192 32496 22244 32502
rect 22020 32434 22140 32450
rect 22192 32438 22244 32444
rect 22020 32428 22152 32434
rect 22020 32422 22100 32428
rect 21916 31952 21968 31958
rect 21916 31894 21968 31900
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 21928 29306 21956 31758
rect 22020 29578 22048 32422
rect 22100 32370 22152 32376
rect 22204 32026 22232 32438
rect 22192 32020 22244 32026
rect 22192 31962 22244 31968
rect 22100 31952 22152 31958
rect 22100 31894 22152 31900
rect 22112 31822 22140 31894
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 22100 31340 22152 31346
rect 22100 31282 22152 31288
rect 22112 29889 22140 31282
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22098 29880 22154 29889
rect 22098 29815 22154 29824
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 22008 29572 22060 29578
rect 22008 29514 22060 29520
rect 21916 29300 21968 29306
rect 21916 29242 21968 29248
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21836 28558 21864 28970
rect 22008 28960 22060 28966
rect 22008 28902 22060 28908
rect 22020 28558 22048 28902
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 21836 27538 21864 28494
rect 22020 28234 22048 28494
rect 21928 28206 22048 28234
rect 21824 27532 21876 27538
rect 21824 27474 21876 27480
rect 21836 25430 21864 27474
rect 21928 27402 21956 28206
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 22020 27334 22048 28018
rect 22008 27328 22060 27334
rect 22008 27270 22060 27276
rect 21824 25424 21876 25430
rect 21824 25366 21876 25372
rect 21836 24750 21864 25366
rect 21914 24848 21970 24857
rect 21914 24783 21970 24792
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21928 23730 21956 24783
rect 22020 24750 22048 27270
rect 22112 24818 22140 29650
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22008 24744 22060 24750
rect 22008 24686 22060 24692
rect 22112 24274 22140 24754
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 22008 24132 22060 24138
rect 22008 24074 22060 24080
rect 21916 23724 21968 23730
rect 21916 23666 21968 23672
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20364 16046 20392 17070
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20364 15638 20392 15982
rect 20352 15632 20404 15638
rect 20352 15574 20404 15580
rect 20456 15502 20484 16594
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20640 15586 20668 16526
rect 20548 15570 20668 15586
rect 20536 15564 20668 15570
rect 20588 15558 20668 15564
rect 20536 15506 20588 15512
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20272 11762 20300 14418
rect 20364 13394 20392 15030
rect 20456 14346 20484 15438
rect 20628 15428 20680 15434
rect 20628 15370 20680 15376
rect 20640 14414 20668 15370
rect 20732 15026 20760 17138
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 20811 16348 21119 16368
rect 20811 16346 20817 16348
rect 20873 16346 20897 16348
rect 20953 16346 20977 16348
rect 21033 16346 21057 16348
rect 21113 16346 21119 16348
rect 20873 16294 20875 16346
rect 21055 16294 21057 16346
rect 20811 16292 20817 16294
rect 20873 16292 20897 16294
rect 20953 16292 20977 16294
rect 21033 16292 21057 16294
rect 21113 16292 21119 16294
rect 20811 16272 21119 16292
rect 21192 15881 21220 16526
rect 21178 15872 21234 15881
rect 21178 15807 21234 15816
rect 20811 15260 21119 15280
rect 20811 15258 20817 15260
rect 20873 15258 20897 15260
rect 20953 15258 20977 15260
rect 21033 15258 21057 15260
rect 21113 15258 21119 15260
rect 20873 15206 20875 15258
rect 21055 15206 21057 15258
rect 20811 15204 20817 15206
rect 20873 15204 20897 15206
rect 20953 15204 20977 15206
rect 21033 15204 21057 15206
rect 21113 15204 21119 15206
rect 20811 15184 21119 15204
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20364 12306 20392 13330
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20260 11756 20312 11762
rect 20180 11716 20260 11744
rect 20180 11218 20208 11716
rect 20260 11698 20312 11704
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20168 9580 20220 9586
rect 20088 9540 20168 9568
rect 20168 9522 20220 9528
rect 20180 8906 20208 9522
rect 20272 9178 20300 11154
rect 20364 11150 20392 12038
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20456 10826 20484 14282
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20548 13326 20576 14010
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20640 12986 20668 13194
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20732 12866 20760 14962
rect 20916 14482 20944 14962
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20811 14172 21119 14192
rect 20811 14170 20817 14172
rect 20873 14170 20897 14172
rect 20953 14170 20977 14172
rect 21033 14170 21057 14172
rect 21113 14170 21119 14172
rect 20873 14118 20875 14170
rect 21055 14118 21057 14170
rect 20811 14116 20817 14118
rect 20873 14116 20897 14118
rect 20953 14116 20977 14118
rect 21033 14116 21057 14118
rect 21113 14116 21119 14118
rect 20811 14096 21119 14116
rect 20811 13084 21119 13104
rect 20811 13082 20817 13084
rect 20873 13082 20897 13084
rect 20953 13082 20977 13084
rect 21033 13082 21057 13084
rect 21113 13082 21119 13084
rect 20873 13030 20875 13082
rect 21055 13030 21057 13082
rect 20811 13028 20817 13030
rect 20873 13028 20897 13030
rect 20953 13028 20977 13030
rect 21033 13028 21057 13030
rect 21113 13028 21119 13030
rect 20811 13008 21119 13028
rect 20628 12844 20680 12850
rect 20732 12838 20852 12866
rect 20628 12786 20680 12792
rect 20640 11898 20668 12786
rect 20824 12782 20852 12838
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20824 12594 20852 12718
rect 20824 12566 20944 12594
rect 20916 12434 20944 12566
rect 20824 12406 20944 12434
rect 20720 12232 20772 12238
rect 20824 12186 20852 12406
rect 20772 12180 20852 12186
rect 20720 12174 20852 12180
rect 20732 12158 20852 12174
rect 20811 11996 21119 12016
rect 20811 11994 20817 11996
rect 20873 11994 20897 11996
rect 20953 11994 20977 11996
rect 21033 11994 21057 11996
rect 21113 11994 21119 11996
rect 20873 11942 20875 11994
rect 21055 11942 21057 11994
rect 20811 11940 20817 11942
rect 20873 11940 20897 11942
rect 20953 11940 20977 11942
rect 21033 11940 21057 11942
rect 21113 11940 21119 11942
rect 20811 11920 21119 11940
rect 20628 11892 20680 11898
rect 20364 10810 20484 10826
rect 20352 10804 20484 10810
rect 20404 10798 20484 10804
rect 20548 11852 20628 11880
rect 20352 10746 20404 10752
rect 20364 10062 20392 10746
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20364 9722 20392 9998
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20456 9586 20484 10678
rect 20548 10674 20576 11852
rect 20628 11834 20680 11840
rect 21192 11354 21220 14962
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 12782 21312 13262
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21376 11762 21404 13126
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21376 11257 21404 11290
rect 21362 11248 21418 11257
rect 21362 11183 21418 11192
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20548 10130 20576 10610
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20456 9110 20484 9522
rect 20548 9518 20576 10066
rect 20640 9654 20668 11086
rect 21468 11082 21496 17614
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21560 15502 21588 17274
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21640 15564 21692 15570
rect 21640 15506 21692 15512
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21560 13326 21588 14894
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 20811 10908 21119 10928
rect 20811 10906 20817 10908
rect 20873 10906 20897 10908
rect 20953 10906 20977 10908
rect 21033 10906 21057 10908
rect 21113 10906 21119 10908
rect 20873 10854 20875 10906
rect 21055 10854 21057 10906
rect 20811 10852 20817 10854
rect 20873 10852 20897 10854
rect 20953 10852 20977 10854
rect 21033 10852 21057 10854
rect 21113 10852 21119 10854
rect 20811 10832 21119 10852
rect 21192 10062 21220 11018
rect 21560 10606 21588 13262
rect 21652 11218 21680 15506
rect 21836 14618 21864 16050
rect 21928 15978 21956 23530
rect 22020 17882 22048 24074
rect 22204 24070 22232 31214
rect 22296 27130 22324 35566
rect 22480 32910 22508 36196
rect 22560 36100 22612 36106
rect 22560 36042 22612 36048
rect 22468 32904 22520 32910
rect 22468 32846 22520 32852
rect 22480 32502 22508 32846
rect 22468 32496 22520 32502
rect 22468 32438 22520 32444
rect 22376 32360 22428 32366
rect 22376 32302 22428 32308
rect 22388 29170 22416 32302
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 22480 28082 22508 31826
rect 22572 31414 22600 36042
rect 22756 32434 22784 38694
rect 22848 36530 22876 45970
rect 22940 41018 22968 46430
rect 23112 46378 23164 46384
rect 23020 46368 23072 46374
rect 23020 46310 23072 46316
rect 23032 45966 23060 46310
rect 23020 45960 23072 45966
rect 23020 45902 23072 45908
rect 23020 45824 23072 45830
rect 23020 45766 23072 45772
rect 23032 41721 23060 45766
rect 23018 41712 23074 41721
rect 23018 41647 23074 41656
rect 23124 41274 23152 46378
rect 23216 41414 23244 55014
rect 23308 54194 23336 55218
rect 23400 54534 23428 56714
rect 23388 54528 23440 54534
rect 23388 54470 23440 54476
rect 23296 54188 23348 54194
rect 23296 54130 23348 54136
rect 23296 53032 23348 53038
rect 23296 52974 23348 52980
rect 23308 52698 23336 52974
rect 23296 52692 23348 52698
rect 23296 52634 23348 52640
rect 23308 51474 23336 52634
rect 23296 51468 23348 51474
rect 23492 51456 23520 56918
rect 23584 56681 23612 60454
rect 23676 58546 23704 63378
rect 23664 58540 23716 58546
rect 23664 58482 23716 58488
rect 23676 58002 23704 58482
rect 23664 57996 23716 58002
rect 23664 57938 23716 57944
rect 23664 57044 23716 57050
rect 23664 56986 23716 56992
rect 23570 56672 23626 56681
rect 23570 56607 23626 56616
rect 23572 56500 23624 56506
rect 23572 56442 23624 56448
rect 23584 55078 23612 56442
rect 23676 55418 23704 56986
rect 23664 55412 23716 55418
rect 23664 55354 23716 55360
rect 23664 55140 23716 55146
rect 23664 55082 23716 55088
rect 23572 55072 23624 55078
rect 23572 55014 23624 55020
rect 23584 52154 23612 55014
rect 23676 54874 23704 55082
rect 23664 54868 23716 54874
rect 23664 54810 23716 54816
rect 23664 54732 23716 54738
rect 23664 54674 23716 54680
rect 23676 53106 23704 54674
rect 23664 53100 23716 53106
rect 23664 53042 23716 53048
rect 23676 53009 23704 53042
rect 23662 53000 23718 53009
rect 23662 52935 23718 52944
rect 23664 52896 23716 52902
rect 23662 52864 23664 52873
rect 23716 52864 23718 52873
rect 23662 52799 23718 52808
rect 23768 52714 23796 64942
rect 23848 63368 23900 63374
rect 23848 63310 23900 63316
rect 23860 62898 23888 63310
rect 23952 63306 23980 66982
rect 24228 66570 24256 70042
rect 24768 68944 24820 68950
rect 24768 68886 24820 68892
rect 24216 66564 24268 66570
rect 24216 66506 24268 66512
rect 24124 64320 24176 64326
rect 24124 64262 24176 64268
rect 24032 63912 24084 63918
rect 24032 63854 24084 63860
rect 23940 63300 23992 63306
rect 23940 63242 23992 63248
rect 23848 62892 23900 62898
rect 23848 62834 23900 62840
rect 23860 61810 23888 62834
rect 24044 62694 24072 63854
rect 24136 63782 24164 64262
rect 24124 63776 24176 63782
rect 24124 63718 24176 63724
rect 24032 62688 24084 62694
rect 24032 62630 24084 62636
rect 23848 61804 23900 61810
rect 23848 61746 23900 61752
rect 23860 59650 23888 61746
rect 23940 61260 23992 61266
rect 23940 61202 23992 61208
rect 23952 60314 23980 61202
rect 23940 60308 23992 60314
rect 23940 60250 23992 60256
rect 23860 59634 23980 59650
rect 23860 59628 23992 59634
rect 23860 59622 23940 59628
rect 23940 59570 23992 59576
rect 23848 58948 23900 58954
rect 23848 58890 23900 58896
rect 23860 55865 23888 58890
rect 23952 57458 23980 59570
rect 23940 57452 23992 57458
rect 23940 57394 23992 57400
rect 23846 55856 23902 55865
rect 23846 55791 23902 55800
rect 23846 55176 23902 55185
rect 23846 55111 23902 55120
rect 23860 53689 23888 55111
rect 23846 53680 23902 53689
rect 23846 53615 23902 53624
rect 23676 52686 23796 52714
rect 23572 52148 23624 52154
rect 23572 52090 23624 52096
rect 23296 51410 23348 51416
rect 23400 51428 23520 51456
rect 23400 51354 23428 51428
rect 23308 51326 23428 51354
rect 23478 51368 23534 51377
rect 23308 50998 23336 51326
rect 23478 51303 23534 51312
rect 23388 51264 23440 51270
rect 23388 51206 23440 51212
rect 23492 51218 23520 51303
rect 23296 50992 23348 50998
rect 23296 50934 23348 50940
rect 23400 50862 23428 51206
rect 23492 51190 23612 51218
rect 23480 50924 23532 50930
rect 23480 50866 23532 50872
rect 23388 50856 23440 50862
rect 23388 50798 23440 50804
rect 23400 50708 23428 50798
rect 23308 50680 23428 50708
rect 23308 49706 23336 50680
rect 23386 49872 23442 49881
rect 23386 49807 23442 49816
rect 23296 49700 23348 49706
rect 23296 49642 23348 49648
rect 23400 49366 23428 49807
rect 23492 49774 23520 50866
rect 23480 49768 23532 49774
rect 23480 49710 23532 49716
rect 23388 49360 23440 49366
rect 23388 49302 23440 49308
rect 23296 49224 23348 49230
rect 23296 49166 23348 49172
rect 23308 48754 23336 49166
rect 23296 48748 23348 48754
rect 23296 48690 23348 48696
rect 23308 46442 23336 48690
rect 23480 48680 23532 48686
rect 23480 48622 23532 48628
rect 23492 47258 23520 48622
rect 23480 47252 23532 47258
rect 23480 47194 23532 47200
rect 23388 46912 23440 46918
rect 23388 46854 23440 46860
rect 23400 46646 23428 46854
rect 23388 46640 23440 46646
rect 23388 46582 23440 46588
rect 23296 46436 23348 46442
rect 23296 46378 23348 46384
rect 23400 46322 23428 46582
rect 23480 46572 23532 46578
rect 23480 46514 23532 46520
rect 23308 46294 23428 46322
rect 23308 45830 23336 46294
rect 23388 46164 23440 46170
rect 23388 46106 23440 46112
rect 23296 45824 23348 45830
rect 23296 45766 23348 45772
rect 23308 44470 23336 45766
rect 23296 44464 23348 44470
rect 23296 44406 23348 44412
rect 23296 44192 23348 44198
rect 23296 44134 23348 44140
rect 23308 43217 23336 44134
rect 23294 43208 23350 43217
rect 23294 43143 23350 43152
rect 23296 43104 23348 43110
rect 23296 43046 23348 43052
rect 23308 42770 23336 43046
rect 23296 42764 23348 42770
rect 23296 42706 23348 42712
rect 23294 42392 23350 42401
rect 23294 42327 23296 42336
rect 23348 42327 23350 42336
rect 23296 42298 23348 42304
rect 23216 41386 23336 41414
rect 23112 41268 23164 41274
rect 23112 41210 23164 41216
rect 23204 41132 23256 41138
rect 23204 41074 23256 41080
rect 22940 40990 23152 41018
rect 22928 40928 22980 40934
rect 22928 40870 22980 40876
rect 22940 39438 22968 40870
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 23020 39024 23072 39030
rect 23020 38966 23072 38972
rect 22928 38820 22980 38826
rect 22928 38762 22980 38768
rect 22940 38554 22968 38762
rect 22928 38548 22980 38554
rect 22928 38490 22980 38496
rect 22928 38412 22980 38418
rect 22928 38354 22980 38360
rect 22940 37913 22968 38354
rect 22926 37904 22982 37913
rect 22926 37839 22982 37848
rect 22926 36952 22982 36961
rect 23032 36922 23060 38966
rect 22926 36887 22982 36896
rect 23020 36916 23072 36922
rect 22940 36854 22968 36887
rect 23020 36858 23072 36864
rect 22928 36848 22980 36854
rect 22928 36790 22980 36796
rect 22848 36502 23060 36530
rect 22928 36100 22980 36106
rect 22928 36042 22980 36048
rect 22940 33114 22968 36042
rect 22928 33108 22980 33114
rect 22928 33050 22980 33056
rect 22928 32904 22980 32910
rect 22926 32872 22928 32881
rect 22980 32872 22982 32881
rect 22926 32807 22982 32816
rect 22744 32428 22796 32434
rect 22744 32370 22796 32376
rect 23032 32298 23060 36502
rect 23124 35290 23152 40990
rect 23216 40186 23244 41074
rect 23308 41018 23336 41386
rect 23400 41138 23428 46106
rect 23492 41585 23520 46514
rect 23584 41698 23612 51190
rect 23676 50182 23704 52686
rect 23756 52556 23808 52562
rect 23756 52498 23808 52504
rect 23768 50969 23796 52498
rect 23860 51814 23888 53615
rect 23952 52426 23980 57394
rect 24044 54738 24072 62630
rect 24124 61804 24176 61810
rect 24124 61746 24176 61752
rect 24136 60858 24164 61746
rect 24124 60852 24176 60858
rect 24124 60794 24176 60800
rect 24122 59120 24178 59129
rect 24122 59055 24178 59064
rect 24136 57361 24164 59055
rect 24122 57352 24178 57361
rect 24122 57287 24178 57296
rect 24124 57248 24176 57254
rect 24124 57190 24176 57196
rect 24136 56846 24164 57190
rect 24124 56840 24176 56846
rect 24124 56782 24176 56788
rect 24136 56370 24164 56782
rect 24228 56438 24256 66506
rect 24676 66496 24728 66502
rect 24676 66438 24728 66444
rect 24688 65958 24716 66438
rect 24676 65952 24728 65958
rect 24676 65894 24728 65900
rect 24308 65680 24360 65686
rect 24308 65622 24360 65628
rect 24216 56432 24268 56438
rect 24216 56374 24268 56380
rect 24124 56364 24176 56370
rect 24124 56306 24176 56312
rect 24124 56228 24176 56234
rect 24124 56170 24176 56176
rect 24032 54732 24084 54738
rect 24032 54674 24084 54680
rect 24032 53984 24084 53990
rect 24032 53926 24084 53932
rect 24044 53417 24072 53926
rect 24030 53408 24086 53417
rect 24030 53343 24086 53352
rect 23940 52420 23992 52426
rect 23940 52362 23992 52368
rect 23938 52320 23994 52329
rect 23938 52255 23994 52264
rect 23848 51808 23900 51814
rect 23848 51750 23900 51756
rect 23846 51504 23902 51513
rect 23846 51439 23902 51448
rect 23754 50960 23810 50969
rect 23754 50895 23810 50904
rect 23756 50788 23808 50794
rect 23756 50730 23808 50736
rect 23768 50425 23796 50730
rect 23754 50416 23810 50425
rect 23754 50351 23756 50360
rect 23808 50351 23810 50360
rect 23756 50322 23808 50328
rect 23756 50288 23808 50294
rect 23756 50230 23808 50236
rect 23664 50176 23716 50182
rect 23664 50118 23716 50124
rect 23662 50008 23718 50017
rect 23768 49978 23796 50230
rect 23662 49943 23718 49952
rect 23756 49972 23808 49978
rect 23676 44878 23704 49943
rect 23756 49914 23808 49920
rect 23756 49768 23808 49774
rect 23756 49710 23808 49716
rect 23768 45830 23796 49710
rect 23756 45824 23808 45830
rect 23756 45766 23808 45772
rect 23756 45484 23808 45490
rect 23756 45426 23808 45432
rect 23768 44878 23796 45426
rect 23664 44872 23716 44878
rect 23664 44814 23716 44820
rect 23756 44872 23808 44878
rect 23756 44814 23808 44820
rect 23664 44736 23716 44742
rect 23664 44678 23716 44684
rect 23676 44538 23704 44678
rect 23664 44532 23716 44538
rect 23664 44474 23716 44480
rect 23676 43858 23704 44474
rect 23756 44396 23808 44402
rect 23756 44338 23808 44344
rect 23768 43926 23796 44338
rect 23756 43920 23808 43926
rect 23756 43862 23808 43868
rect 23664 43852 23716 43858
rect 23664 43794 23716 43800
rect 23676 43314 23704 43794
rect 23756 43784 23808 43790
rect 23754 43752 23756 43761
rect 23808 43752 23810 43761
rect 23754 43687 23810 43696
rect 23756 43648 23808 43654
rect 23756 43590 23808 43596
rect 23664 43308 23716 43314
rect 23664 43250 23716 43256
rect 23664 43172 23716 43178
rect 23664 43114 23716 43120
rect 23676 42906 23704 43114
rect 23664 42900 23716 42906
rect 23664 42842 23716 42848
rect 23584 41670 23704 41698
rect 23572 41608 23624 41614
rect 23478 41576 23534 41585
rect 23572 41550 23624 41556
rect 23478 41511 23534 41520
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 23308 40990 23428 41018
rect 23584 41002 23612 41550
rect 23296 40928 23348 40934
rect 23294 40896 23296 40905
rect 23348 40896 23350 40905
rect 23294 40831 23350 40840
rect 23204 40180 23256 40186
rect 23204 40122 23256 40128
rect 23296 39976 23348 39982
rect 23296 39918 23348 39924
rect 23204 39636 23256 39642
rect 23204 39578 23256 39584
rect 23216 35698 23244 39578
rect 23308 39438 23336 39918
rect 23296 39432 23348 39438
rect 23296 39374 23348 39380
rect 23400 39250 23428 40990
rect 23572 40996 23624 41002
rect 23572 40938 23624 40944
rect 23480 40724 23532 40730
rect 23480 40666 23532 40672
rect 23492 40594 23520 40666
rect 23480 40588 23532 40594
rect 23480 40530 23532 40536
rect 23492 39982 23520 40530
rect 23572 40520 23624 40526
rect 23572 40462 23624 40468
rect 23584 40050 23612 40462
rect 23572 40044 23624 40050
rect 23572 39986 23624 39992
rect 23480 39976 23532 39982
rect 23480 39918 23532 39924
rect 23480 39840 23532 39846
rect 23480 39782 23532 39788
rect 23308 39222 23428 39250
rect 23204 35692 23256 35698
rect 23204 35634 23256 35640
rect 23112 35284 23164 35290
rect 23112 35226 23164 35232
rect 22744 32292 22796 32298
rect 22744 32234 22796 32240
rect 23020 32292 23072 32298
rect 23020 32234 23072 32240
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22560 31408 22612 31414
rect 22560 31350 22612 31356
rect 22560 30796 22612 30802
rect 22560 30738 22612 30744
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22376 27328 22428 27334
rect 22376 27270 22428 27276
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 22296 24410 22324 26930
rect 22388 26042 22416 27270
rect 22480 26858 22508 28018
rect 22572 27334 22600 30738
rect 22664 29170 22692 31962
rect 22756 29714 22784 32234
rect 23216 32201 23244 35634
rect 23308 33998 23336 39222
rect 23492 38654 23520 39782
rect 23572 39092 23624 39098
rect 23572 39034 23624 39040
rect 23584 38894 23612 39034
rect 23572 38888 23624 38894
rect 23572 38830 23624 38836
rect 23400 38626 23520 38654
rect 23400 38536 23428 38626
rect 23400 38508 23520 38536
rect 23386 38448 23442 38457
rect 23386 38383 23388 38392
rect 23440 38383 23442 38392
rect 23388 38354 23440 38360
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23202 32192 23258 32201
rect 23202 32127 23258 32136
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23112 31748 23164 31754
rect 23112 31690 23164 31696
rect 22926 31512 22982 31521
rect 23124 31482 23152 31690
rect 22926 31447 22982 31456
rect 23112 31476 23164 31482
rect 22744 29708 22796 29714
rect 22744 29650 22796 29656
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22848 29306 22876 29582
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22744 29232 22796 29238
rect 22744 29174 22796 29180
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22560 27124 22612 27130
rect 22560 27066 22612 27072
rect 22468 26852 22520 26858
rect 22468 26794 22520 26800
rect 22376 26036 22428 26042
rect 22376 25978 22428 25984
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22388 25294 22416 25842
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 22376 25152 22428 25158
rect 22376 25094 22428 25100
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22112 22710 22140 23598
rect 22204 22778 22232 23666
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21928 15570 21956 15914
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21836 14006 21864 14554
rect 21824 14000 21876 14006
rect 21824 13942 21876 13948
rect 22112 12986 22140 22170
rect 22296 22030 22324 24346
rect 22388 23225 22416 25094
rect 22374 23216 22430 23225
rect 22374 23151 22430 23160
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 22388 22710 22416 23054
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22376 22500 22428 22506
rect 22376 22442 22428 22448
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22388 21554 22416 22442
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22480 19854 22508 26794
rect 22572 22234 22600 27066
rect 22664 25974 22692 29106
rect 22652 25968 22704 25974
rect 22652 25910 22704 25916
rect 22756 25906 22784 29174
rect 22836 29096 22888 29102
rect 22836 29038 22888 29044
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 22756 25786 22784 25842
rect 22664 25758 22784 25786
rect 22664 25294 22692 25758
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22664 23866 22692 24686
rect 22756 24614 22784 25230
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22756 23730 22784 24006
rect 22848 23866 22876 29038
rect 22940 26382 22968 31447
rect 23112 31418 23164 31424
rect 23020 31340 23072 31346
rect 23020 31282 23072 31288
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 22928 26036 22980 26042
rect 22928 25978 22980 25984
rect 22940 25362 22968 25978
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 22926 24848 22982 24857
rect 22926 24783 22928 24792
rect 22980 24783 22982 24792
rect 22928 24754 22980 24760
rect 22940 24206 22968 24754
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22664 22778 22692 23258
rect 22652 22772 22704 22778
rect 22652 22714 22704 22720
rect 22650 22672 22706 22681
rect 22650 22607 22706 22616
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22572 18986 22600 21830
rect 22480 18958 22600 18986
rect 22480 18834 22508 18958
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22480 18358 22508 18770
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22388 17338 22416 18226
rect 22480 17678 22508 18294
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22480 15162 22508 17614
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22480 14618 22508 14962
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22664 13988 22692 22607
rect 22756 21962 22784 23666
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22848 18426 22876 23122
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22940 22642 22968 23054
rect 23032 22982 23060 31282
rect 23216 31142 23244 31962
rect 23308 31634 23336 32710
rect 23400 31777 23428 36518
rect 23386 31768 23442 31777
rect 23386 31703 23442 31712
rect 23308 31606 23428 31634
rect 23294 31512 23350 31521
rect 23294 31447 23350 31456
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 23204 30864 23256 30870
rect 23204 30806 23256 30812
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 23124 29170 23152 29514
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 23216 28218 23244 30806
rect 23204 28212 23256 28218
rect 23204 28154 23256 28160
rect 23112 28144 23164 28150
rect 23112 28086 23164 28092
rect 23124 23866 23152 28086
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23216 27130 23244 28018
rect 23204 27124 23256 27130
rect 23204 27066 23256 27072
rect 23308 27010 23336 31447
rect 23400 29306 23428 31606
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23492 28994 23520 38508
rect 23584 38486 23612 38830
rect 23676 38826 23704 41670
rect 23664 38820 23716 38826
rect 23664 38762 23716 38768
rect 23768 38706 23796 43590
rect 23860 39001 23888 51439
rect 23952 51066 23980 52255
rect 24032 51468 24084 51474
rect 24032 51410 24084 51416
rect 23940 51060 23992 51066
rect 23940 51002 23992 51008
rect 23940 50448 23992 50454
rect 23940 50390 23992 50396
rect 23952 50164 23980 50390
rect 24044 50318 24072 51410
rect 24032 50312 24084 50318
rect 24032 50254 24084 50260
rect 23952 50136 24072 50164
rect 23938 50008 23994 50017
rect 23938 49943 23994 49952
rect 23952 40644 23980 49943
rect 24044 47258 24072 50136
rect 24032 47252 24084 47258
rect 24032 47194 24084 47200
rect 24032 45824 24084 45830
rect 24032 45766 24084 45772
rect 24044 45422 24072 45766
rect 24032 45416 24084 45422
rect 24032 45358 24084 45364
rect 24044 43790 24072 45358
rect 24032 43784 24084 43790
rect 24032 43726 24084 43732
rect 24032 43240 24084 43246
rect 24030 43208 24032 43217
rect 24084 43208 24086 43217
rect 24030 43143 24086 43152
rect 24030 43072 24086 43081
rect 24030 43007 24086 43016
rect 24044 42265 24072 43007
rect 24030 42256 24086 42265
rect 24030 42191 24086 42200
rect 24032 41540 24084 41546
rect 24032 41482 24084 41488
rect 24044 40769 24072 41482
rect 24030 40760 24086 40769
rect 24030 40695 24086 40704
rect 23952 40616 24072 40644
rect 23846 38992 23902 39001
rect 23846 38927 23902 38936
rect 23676 38678 23796 38706
rect 23848 38752 23900 38758
rect 23848 38694 23900 38700
rect 23676 38486 23704 38678
rect 23572 38480 23624 38486
rect 23572 38422 23624 38428
rect 23664 38480 23716 38486
rect 23664 38422 23716 38428
rect 23860 38298 23888 38694
rect 24044 38418 24072 40616
rect 24032 38412 24084 38418
rect 24032 38354 24084 38360
rect 24136 38298 24164 56170
rect 24216 56160 24268 56166
rect 24216 56102 24268 56108
rect 24228 55622 24256 56102
rect 24216 55616 24268 55622
rect 24216 55558 24268 55564
rect 24214 55448 24270 55457
rect 24214 55383 24270 55392
rect 24228 55146 24256 55383
rect 24216 55140 24268 55146
rect 24216 55082 24268 55088
rect 24228 54913 24256 55082
rect 24214 54904 24270 54913
rect 24214 54839 24270 54848
rect 24216 54528 24268 54534
rect 24216 54470 24268 54476
rect 24228 51882 24256 54470
rect 24320 52562 24348 65622
rect 24584 65544 24636 65550
rect 24584 65486 24636 65492
rect 24400 64524 24452 64530
rect 24400 64466 24452 64472
rect 24412 62490 24440 64466
rect 24492 64388 24544 64394
rect 24492 64330 24544 64336
rect 24400 62484 24452 62490
rect 24400 62426 24452 62432
rect 24504 61962 24532 64330
rect 24596 63442 24624 65486
rect 24780 64394 24808 68886
rect 24964 67658 24992 75142
rect 25776 74556 26084 74576
rect 25776 74554 25782 74556
rect 25838 74554 25862 74556
rect 25918 74554 25942 74556
rect 25998 74554 26022 74556
rect 26078 74554 26084 74556
rect 25838 74502 25840 74554
rect 26020 74502 26022 74554
rect 25776 74500 25782 74502
rect 25838 74500 25862 74502
rect 25918 74500 25942 74502
rect 25998 74500 26022 74502
rect 26078 74500 26084 74502
rect 25776 74480 26084 74500
rect 26240 74248 26292 74254
rect 26240 74190 26292 74196
rect 25776 73468 26084 73488
rect 25776 73466 25782 73468
rect 25838 73466 25862 73468
rect 25918 73466 25942 73468
rect 25998 73466 26022 73468
rect 26078 73466 26084 73468
rect 25838 73414 25840 73466
rect 26020 73414 26022 73466
rect 25776 73412 25782 73414
rect 25838 73412 25862 73414
rect 25918 73412 25942 73414
rect 25998 73412 26022 73414
rect 26078 73412 26084 73414
rect 25776 73392 26084 73412
rect 26148 73092 26200 73098
rect 26148 73034 26200 73040
rect 25776 72380 26084 72400
rect 25776 72378 25782 72380
rect 25838 72378 25862 72380
rect 25918 72378 25942 72380
rect 25998 72378 26022 72380
rect 26078 72378 26084 72380
rect 25838 72326 25840 72378
rect 26020 72326 26022 72378
rect 25776 72324 25782 72326
rect 25838 72324 25862 72326
rect 25918 72324 25942 72326
rect 25998 72324 26022 72326
rect 26078 72324 26084 72326
rect 25776 72304 26084 72324
rect 25776 71292 26084 71312
rect 25776 71290 25782 71292
rect 25838 71290 25862 71292
rect 25918 71290 25942 71292
rect 25998 71290 26022 71292
rect 26078 71290 26084 71292
rect 25838 71238 25840 71290
rect 26020 71238 26022 71290
rect 25776 71236 25782 71238
rect 25838 71236 25862 71238
rect 25918 71236 25942 71238
rect 25998 71236 26022 71238
rect 26078 71236 26084 71238
rect 25776 71216 26084 71236
rect 25776 70204 26084 70224
rect 25776 70202 25782 70204
rect 25838 70202 25862 70204
rect 25918 70202 25942 70204
rect 25998 70202 26022 70204
rect 26078 70202 26084 70204
rect 25838 70150 25840 70202
rect 26020 70150 26022 70202
rect 25776 70148 25782 70150
rect 25838 70148 25862 70150
rect 25918 70148 25942 70150
rect 25998 70148 26022 70150
rect 26078 70148 26084 70150
rect 25776 70128 26084 70148
rect 25504 69760 25556 69766
rect 25504 69702 25556 69708
rect 25042 68232 25098 68241
rect 25042 68167 25098 68176
rect 24952 67652 25004 67658
rect 24952 67594 25004 67600
rect 25056 67266 25084 68167
rect 25136 67720 25188 67726
rect 25136 67662 25188 67668
rect 25412 67720 25464 67726
rect 25412 67662 25464 67668
rect 24964 67238 25084 67266
rect 25148 67250 25176 67662
rect 25228 67652 25280 67658
rect 25228 67594 25280 67600
rect 25240 67266 25268 67594
rect 25136 67244 25188 67250
rect 24860 67040 24912 67046
rect 24860 66982 24912 66988
rect 24872 64666 24900 66982
rect 24860 64660 24912 64666
rect 24860 64602 24912 64608
rect 24964 64546 24992 67238
rect 25240 67238 25360 67266
rect 25424 67250 25452 67662
rect 25136 67186 25188 67192
rect 25148 67130 25176 67186
rect 25044 67108 25096 67114
rect 25148 67102 25268 67130
rect 25044 67050 25096 67056
rect 24872 64518 24992 64546
rect 24768 64388 24820 64394
rect 24768 64330 24820 64336
rect 24676 64320 24728 64326
rect 24676 64262 24728 64268
rect 24688 64054 24716 64262
rect 24676 64048 24728 64054
rect 24872 64002 24900 64518
rect 24952 64456 25004 64462
rect 24952 64398 25004 64404
rect 24676 63990 24728 63996
rect 24780 63974 24900 64002
rect 24780 63730 24808 63974
rect 24688 63702 24808 63730
rect 24584 63436 24636 63442
rect 24584 63378 24636 63384
rect 24584 63300 24636 63306
rect 24584 63242 24636 63248
rect 24596 62830 24624 63242
rect 24584 62824 24636 62830
rect 24584 62766 24636 62772
rect 24504 61934 24624 61962
rect 24492 61804 24544 61810
rect 24492 61746 24544 61752
rect 24400 60580 24452 60586
rect 24400 60522 24452 60528
rect 24412 58954 24440 60522
rect 24400 58948 24452 58954
rect 24400 58890 24452 58896
rect 24400 58540 24452 58546
rect 24400 58482 24452 58488
rect 24412 57254 24440 58482
rect 24400 57248 24452 57254
rect 24400 57190 24452 57196
rect 24504 56982 24532 61746
rect 24596 61282 24624 61934
rect 24688 61402 24716 63702
rect 24964 63374 24992 64398
rect 25056 63866 25084 67050
rect 25240 66638 25268 67102
rect 25228 66632 25280 66638
rect 25228 66574 25280 66580
rect 25136 66564 25188 66570
rect 25136 66506 25188 66512
rect 25148 64462 25176 66506
rect 25240 66162 25268 66574
rect 25228 66156 25280 66162
rect 25228 66098 25280 66104
rect 25240 65618 25268 66098
rect 25228 65612 25280 65618
rect 25228 65554 25280 65560
rect 25228 64660 25280 64666
rect 25228 64602 25280 64608
rect 25136 64456 25188 64462
rect 25136 64398 25188 64404
rect 25148 63986 25176 64398
rect 25240 64326 25268 64602
rect 25228 64320 25280 64326
rect 25228 64262 25280 64268
rect 25136 63980 25188 63986
rect 25136 63922 25188 63928
rect 25056 63838 25176 63866
rect 24952 63368 25004 63374
rect 24952 63310 25004 63316
rect 24964 62422 24992 63310
rect 24952 62416 25004 62422
rect 24858 62384 24914 62393
rect 24952 62358 25004 62364
rect 24858 62319 24914 62328
rect 24872 62286 24900 62319
rect 24860 62280 24912 62286
rect 24860 62222 24912 62228
rect 24766 62112 24822 62121
rect 24766 62047 24822 62056
rect 24780 61946 24808 62047
rect 24768 61940 24820 61946
rect 24768 61882 24820 61888
rect 24964 61826 24992 62358
rect 25044 61940 25096 61946
rect 25044 61882 25096 61888
rect 24872 61810 24992 61826
rect 24860 61804 24992 61810
rect 24912 61798 24992 61804
rect 24860 61746 24912 61752
rect 24858 61704 24914 61713
rect 24858 61639 24914 61648
rect 24676 61396 24728 61402
rect 24676 61338 24728 61344
rect 24596 61254 24808 61282
rect 24872 61266 24900 61639
rect 24964 61606 24992 61798
rect 25056 61713 25084 61882
rect 25042 61704 25098 61713
rect 25042 61639 25098 61648
rect 24952 61600 25004 61606
rect 24952 61542 25004 61548
rect 25044 61600 25096 61606
rect 25044 61542 25096 61548
rect 24584 61056 24636 61062
rect 24584 60998 24636 61004
rect 24596 60489 24624 60998
rect 24676 60852 24728 60858
rect 24676 60794 24728 60800
rect 24582 60480 24638 60489
rect 24582 60415 24638 60424
rect 24582 60344 24638 60353
rect 24582 60279 24638 60288
rect 24492 56976 24544 56982
rect 24596 56953 24624 60279
rect 24688 60081 24716 60794
rect 24674 60072 24730 60081
rect 24674 60007 24730 60016
rect 24492 56918 24544 56924
rect 24582 56944 24638 56953
rect 24582 56879 24638 56888
rect 24584 56840 24636 56846
rect 24398 56808 24454 56817
rect 24584 56782 24636 56788
rect 24398 56743 24400 56752
rect 24452 56743 24454 56752
rect 24400 56714 24452 56720
rect 24492 56704 24544 56710
rect 24492 56646 24544 56652
rect 24400 56500 24452 56506
rect 24504 56488 24532 56646
rect 24452 56460 24532 56488
rect 24400 56442 24452 56448
rect 24400 56364 24452 56370
rect 24400 56306 24452 56312
rect 24412 55962 24440 56306
rect 24504 55962 24532 56460
rect 24596 55962 24624 56782
rect 24400 55956 24452 55962
rect 24400 55898 24452 55904
rect 24492 55956 24544 55962
rect 24492 55898 24544 55904
rect 24584 55956 24636 55962
rect 24584 55898 24636 55904
rect 24400 55820 24452 55826
rect 24400 55762 24452 55768
rect 24412 53650 24440 55762
rect 24584 55752 24636 55758
rect 24584 55694 24636 55700
rect 24492 55684 24544 55690
rect 24492 55626 24544 55632
rect 24504 55214 24532 55626
rect 24596 55282 24624 55694
rect 24584 55276 24636 55282
rect 24584 55218 24636 55224
rect 24492 55208 24544 55214
rect 24492 55150 24544 55156
rect 24504 53990 24532 55150
rect 24596 55049 24624 55218
rect 24582 55040 24638 55049
rect 24582 54975 24638 54984
rect 24584 54868 24636 54874
rect 24584 54810 24636 54816
rect 24492 53984 24544 53990
rect 24492 53926 24544 53932
rect 24400 53644 24452 53650
rect 24400 53586 24452 53592
rect 24308 52556 24360 52562
rect 24308 52498 24360 52504
rect 24308 52420 24360 52426
rect 24308 52362 24360 52368
rect 24216 51876 24268 51882
rect 24216 51818 24268 51824
rect 24216 51060 24268 51066
rect 24216 51002 24268 51008
rect 24228 41177 24256 51002
rect 24320 43994 24348 52362
rect 24400 52148 24452 52154
rect 24400 52090 24452 52096
rect 24412 51950 24440 52090
rect 24400 51944 24452 51950
rect 24400 51886 24452 51892
rect 24412 51474 24440 51886
rect 24400 51468 24452 51474
rect 24400 51410 24452 51416
rect 24400 51332 24452 51338
rect 24400 51274 24452 51280
rect 24308 43988 24360 43994
rect 24308 43930 24360 43936
rect 24306 43752 24362 43761
rect 24306 43687 24362 43696
rect 24320 41546 24348 43687
rect 24308 41540 24360 41546
rect 24308 41482 24360 41488
rect 24306 41304 24362 41313
rect 24306 41239 24362 41248
rect 24214 41168 24270 41177
rect 24214 41103 24270 41112
rect 24320 40526 24348 41239
rect 24308 40520 24360 40526
rect 24308 40462 24360 40468
rect 24308 40044 24360 40050
rect 24308 39986 24360 39992
rect 23768 38270 23888 38298
rect 23952 38270 24164 38298
rect 23570 38040 23626 38049
rect 23570 37975 23626 37984
rect 23584 32026 23612 37975
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23676 36310 23704 37810
rect 23664 36304 23716 36310
rect 23664 36246 23716 36252
rect 23676 35834 23704 36246
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 23664 32564 23716 32570
rect 23664 32506 23716 32512
rect 23572 32020 23624 32026
rect 23572 31962 23624 31968
rect 23572 31748 23624 31754
rect 23572 31690 23624 31696
rect 23584 31346 23612 31690
rect 23676 31686 23704 32506
rect 23664 31680 23716 31686
rect 23664 31622 23716 31628
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23400 28966 23520 28994
rect 23400 27112 23428 28966
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 23584 27878 23612 28154
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23400 27084 23520 27112
rect 23216 26982 23336 27010
rect 23388 26988 23440 26994
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 23112 23588 23164 23594
rect 23112 23530 23164 23536
rect 23020 22976 23072 22982
rect 23020 22918 23072 22924
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 23124 22420 23152 23530
rect 23216 22642 23244 26982
rect 23388 26930 23440 26936
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23308 23322 23336 24754
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23032 22392 23152 22420
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22940 19514 22968 19722
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22296 13960 22692 13988
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 13530 22232 13670
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22296 13410 22324 13960
rect 22376 13796 22428 13802
rect 22376 13738 22428 13744
rect 22204 13382 22324 13410
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21640 11212 21692 11218
rect 21640 11154 21692 11160
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21468 10130 21496 10406
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 20811 9820 21119 9840
rect 20811 9818 20817 9820
rect 20873 9818 20897 9820
rect 20953 9818 20977 9820
rect 21033 9818 21057 9820
rect 21113 9818 21119 9820
rect 20873 9766 20875 9818
rect 21055 9766 21057 9818
rect 20811 9764 20817 9766
rect 20873 9764 20897 9766
rect 20953 9764 20977 9766
rect 21033 9764 21057 9766
rect 21113 9764 21119 9766
rect 20811 9744 21119 9764
rect 21376 9722 21404 9998
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20548 8974 20576 9454
rect 21560 8974 21588 10542
rect 21652 10130 21680 11154
rect 21928 10266 21956 12174
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20811 8732 21119 8752
rect 20811 8730 20817 8732
rect 20873 8730 20897 8732
rect 20953 8730 20977 8732
rect 21033 8730 21057 8732
rect 21113 8730 21119 8732
rect 20873 8678 20875 8730
rect 21055 8678 21057 8730
rect 20811 8676 20817 8678
rect 20873 8676 20897 8678
rect 20953 8676 20977 8678
rect 21033 8676 21057 8678
rect 21113 8676 21119 8678
rect 20811 8656 21119 8676
rect 20811 7644 21119 7664
rect 20811 7642 20817 7644
rect 20873 7642 20897 7644
rect 20953 7642 20977 7644
rect 21033 7642 21057 7644
rect 21113 7642 21119 7644
rect 20873 7590 20875 7642
rect 21055 7590 21057 7642
rect 20811 7588 20817 7590
rect 20873 7588 20897 7590
rect 20953 7588 20977 7590
rect 21033 7588 21057 7590
rect 21113 7588 21119 7590
rect 20811 7568 21119 7588
rect 16684 6886 16804 6914
rect 18708 6886 18828 6914
rect 10880 6556 11188 6576
rect 10880 6554 10886 6556
rect 10942 6554 10966 6556
rect 11022 6554 11046 6556
rect 11102 6554 11126 6556
rect 11182 6554 11188 6556
rect 10942 6502 10944 6554
rect 11124 6502 11126 6554
rect 10880 6500 10886 6502
rect 10942 6500 10966 6502
rect 11022 6500 11046 6502
rect 11102 6500 11126 6502
rect 11182 6500 11188 6502
rect 10880 6480 11188 6500
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1582 6216 1638 6225
rect 1582 6151 1584 6160
rect 1636 6151 1638 6160
rect 1584 6122 1636 6128
rect 5915 6012 6223 6032
rect 5915 6010 5921 6012
rect 5977 6010 6001 6012
rect 6057 6010 6081 6012
rect 6137 6010 6161 6012
rect 6217 6010 6223 6012
rect 5977 5958 5979 6010
rect 6159 5958 6161 6010
rect 5915 5956 5921 5958
rect 5977 5956 6001 5958
rect 6057 5956 6081 5958
rect 6137 5956 6161 5958
rect 6217 5956 6223 5958
rect 5915 5936 6223 5956
rect 15846 6012 16154 6032
rect 15846 6010 15852 6012
rect 15908 6010 15932 6012
rect 15988 6010 16012 6012
rect 16068 6010 16092 6012
rect 16148 6010 16154 6012
rect 15908 5958 15910 6010
rect 16090 5958 16092 6010
rect 15846 5956 15852 5958
rect 15908 5956 15932 5958
rect 15988 5956 16012 5958
rect 16068 5956 16092 5958
rect 16148 5956 16154 5958
rect 15846 5936 16154 5956
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1582 5471 1638 5480
rect 2700 5234 2728 5714
rect 10880 5468 11188 5488
rect 10880 5466 10886 5468
rect 10942 5466 10966 5468
rect 11022 5466 11046 5468
rect 11102 5466 11126 5468
rect 11182 5466 11188 5468
rect 10942 5414 10944 5466
rect 11124 5414 11126 5466
rect 10880 5412 10886 5414
rect 10942 5412 10966 5414
rect 11022 5412 11046 5414
rect 11102 5412 11126 5414
rect 11182 5412 11188 5414
rect 10880 5392 11188 5412
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 1584 5024 1636 5030
rect 1582 4992 1584 5001
rect 1636 4992 1638 5001
rect 1582 4927 1638 4936
rect 5915 4924 6223 4944
rect 5915 4922 5921 4924
rect 5977 4922 6001 4924
rect 6057 4922 6081 4924
rect 6137 4922 6161 4924
rect 6217 4922 6223 4924
rect 5977 4870 5979 4922
rect 6159 4870 6161 4922
rect 5915 4868 5921 4870
rect 5977 4868 6001 4870
rect 6057 4868 6081 4870
rect 6137 4868 6161 4870
rect 6217 4868 6223 4870
rect 5915 4848 6223 4868
rect 15846 4924 16154 4944
rect 15846 4922 15852 4924
rect 15908 4922 15932 4924
rect 15988 4922 16012 4924
rect 16068 4922 16092 4924
rect 16148 4922 16154 4924
rect 15908 4870 15910 4922
rect 16090 4870 16092 4922
rect 15846 4868 15852 4870
rect 15908 4868 15932 4870
rect 15988 4868 16012 4870
rect 16068 4868 16092 4870
rect 16148 4868 16154 4870
rect 15846 4848 16154 4868
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4321 1624 4422
rect 10880 4380 11188 4400
rect 10880 4378 10886 4380
rect 10942 4378 10966 4380
rect 11022 4378 11046 4380
rect 11102 4378 11126 4380
rect 11182 4378 11188 4380
rect 10942 4326 10944 4378
rect 11124 4326 11126 4378
rect 10880 4324 10886 4326
rect 10942 4324 10966 4326
rect 11022 4324 11046 4326
rect 11102 4324 11126 4326
rect 11182 4324 11188 4326
rect 1582 4312 1638 4321
rect 10880 4304 11188 4324
rect 1582 4247 1638 4256
rect 16684 4146 16712 6886
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 1596 3641 1624 3878
rect 5915 3836 6223 3856
rect 5915 3834 5921 3836
rect 5977 3834 6001 3836
rect 6057 3834 6081 3836
rect 6137 3834 6161 3836
rect 6217 3834 6223 3836
rect 5977 3782 5979 3834
rect 6159 3782 6161 3834
rect 5915 3780 5921 3782
rect 5977 3780 6001 3782
rect 6057 3780 6081 3782
rect 6137 3780 6161 3782
rect 6217 3780 6223 3782
rect 5915 3760 6223 3780
rect 15846 3836 16154 3856
rect 15846 3834 15852 3836
rect 15908 3834 15932 3836
rect 15988 3834 16012 3836
rect 16068 3834 16092 3836
rect 16148 3834 16154 3836
rect 15908 3782 15910 3834
rect 16090 3782 16092 3834
rect 15846 3780 15852 3782
rect 15908 3780 15932 3782
rect 15988 3780 16012 3782
rect 16068 3780 16092 3782
rect 16148 3780 16154 3782
rect 15846 3760 16154 3780
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1596 2961 1624 3334
rect 1582 2952 1638 2961
rect 1582 2887 1638 2896
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 1601 1440 2790
rect 2148 2446 2176 3674
rect 10880 3292 11188 3312
rect 10880 3290 10886 3292
rect 10942 3290 10966 3292
rect 11022 3290 11046 3292
rect 11102 3290 11126 3292
rect 11182 3290 11188 3292
rect 10942 3238 10944 3290
rect 11124 3238 11126 3290
rect 10880 3236 10886 3238
rect 10942 3236 10966 3238
rect 11022 3236 11046 3238
rect 11102 3236 11126 3238
rect 11182 3236 11188 3238
rect 10880 3216 11188 3236
rect 5915 2748 6223 2768
rect 5915 2746 5921 2748
rect 5977 2746 6001 2748
rect 6057 2746 6081 2748
rect 6137 2746 6161 2748
rect 6217 2746 6223 2748
rect 5977 2694 5979 2746
rect 6159 2694 6161 2746
rect 5915 2692 5921 2694
rect 5977 2692 6001 2694
rect 6057 2692 6081 2694
rect 6137 2692 6161 2694
rect 6217 2692 6223 2694
rect 5915 2672 6223 2692
rect 15846 2748 16154 2768
rect 15846 2746 15852 2748
rect 15908 2746 15932 2748
rect 15988 2746 16012 2748
rect 16068 2746 16092 2748
rect 16148 2746 16154 2748
rect 15908 2694 15910 2746
rect 16090 2694 16092 2746
rect 15846 2692 15852 2694
rect 15908 2692 15932 2694
rect 15988 2692 16012 2694
rect 16068 2692 16092 2694
rect 16148 2692 16154 2694
rect 15846 2672 16154 2692
rect 16868 2446 16896 3878
rect 18708 2514 18736 6886
rect 21560 6798 21588 8910
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 20811 6556 21119 6576
rect 20811 6554 20817 6556
rect 20873 6554 20897 6556
rect 20953 6554 20977 6556
rect 21033 6554 21057 6556
rect 21113 6554 21119 6556
rect 20873 6502 20875 6554
rect 21055 6502 21057 6554
rect 20811 6500 20817 6502
rect 20873 6500 20897 6502
rect 20953 6500 20977 6502
rect 21033 6500 21057 6502
rect 21113 6500 21119 6502
rect 20811 6480 21119 6500
rect 22020 6254 22048 6666
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 20811 5468 21119 5488
rect 20811 5466 20817 5468
rect 20873 5466 20897 5468
rect 20953 5466 20977 5468
rect 21033 5466 21057 5468
rect 21113 5466 21119 5468
rect 20873 5414 20875 5466
rect 21055 5414 21057 5466
rect 20811 5412 20817 5414
rect 20873 5412 20897 5414
rect 20953 5412 20977 5414
rect 21033 5412 21057 5414
rect 21113 5412 21119 5414
rect 20811 5392 21119 5412
rect 20811 4380 21119 4400
rect 20811 4378 20817 4380
rect 20873 4378 20897 4380
rect 20953 4378 20977 4380
rect 21033 4378 21057 4380
rect 21113 4378 21119 4380
rect 20873 4326 20875 4378
rect 21055 4326 21057 4378
rect 20811 4324 20817 4326
rect 20873 4324 20897 4326
rect 20953 4324 20977 4326
rect 21033 4324 21057 4326
rect 21113 4324 21119 4326
rect 20811 4304 21119 4324
rect 22020 4078 22048 6190
rect 22204 5302 22232 13382
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22296 5370 22324 12922
rect 22388 9382 22416 13738
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22664 12986 22692 13194
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22664 10266 22692 10610
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22664 8974 22692 9318
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 6662 22692 7686
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 20811 3292 21119 3312
rect 20811 3290 20817 3292
rect 20873 3290 20897 3292
rect 20953 3290 20977 3292
rect 21033 3290 21057 3292
rect 21113 3290 21119 3292
rect 20873 3238 20875 3290
rect 21055 3238 21057 3290
rect 20811 3236 20817 3238
rect 20873 3236 20897 3238
rect 20953 3236 20977 3238
rect 21033 3236 21057 3238
rect 21113 3236 21119 3238
rect 20811 3216 21119 3236
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 1584 2304 1636 2310
rect 2320 2304 2372 2310
rect 1584 2246 1636 2252
rect 2318 2272 2320 2281
rect 2872 2304 2924 2310
rect 2372 2272 2374 2281
rect 1398 1592 1454 1601
rect 1398 1527 1454 1536
rect 1596 921 1624 2246
rect 2872 2246 2924 2252
rect 2318 2207 2374 2216
rect 1582 912 1638 921
rect 1582 847 1638 856
rect 2884 377 2912 2246
rect 10880 2204 11188 2224
rect 10880 2202 10886 2204
rect 10942 2202 10966 2204
rect 11022 2202 11046 2204
rect 11102 2202 11126 2204
rect 11182 2202 11188 2204
rect 10942 2150 10944 2202
rect 11124 2150 11126 2202
rect 10880 2148 10886 2150
rect 10942 2148 10966 2150
rect 11022 2148 11046 2150
rect 11102 2148 11126 2150
rect 11182 2148 11188 2150
rect 10880 2128 11188 2148
rect 20811 2204 21119 2224
rect 20811 2202 20817 2204
rect 20873 2202 20897 2204
rect 20953 2202 20977 2204
rect 21033 2202 21057 2204
rect 21113 2202 21119 2204
rect 20873 2150 20875 2202
rect 21055 2150 21057 2202
rect 20811 2148 20817 2150
rect 20873 2148 20897 2150
rect 20953 2148 20977 2150
rect 21033 2148 21057 2150
rect 21113 2148 21119 2150
rect 20811 2128 21119 2148
rect 22756 1358 22784 17818
rect 22848 17610 22876 18362
rect 22836 17604 22888 17610
rect 22836 17546 22888 17552
rect 22848 17134 22876 17546
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 23032 16946 23060 22392
rect 23400 22094 23428 26930
rect 23492 22642 23520 27084
rect 23584 24138 23612 27814
rect 23676 26790 23704 31078
rect 23664 26784 23716 26790
rect 23664 26726 23716 26732
rect 23572 24132 23624 24138
rect 23572 24074 23624 24080
rect 23584 23526 23612 24074
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23308 22066 23428 22094
rect 23112 21956 23164 21962
rect 23112 21898 23164 21904
rect 23124 18222 23152 21898
rect 23308 21690 23336 22066
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23584 21146 23612 22918
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23216 19310 23244 19994
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23204 19304 23256 19310
rect 23204 19246 23256 19252
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 23216 18970 23244 19110
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 22848 16918 23060 16946
rect 22848 12170 22876 16918
rect 23204 14952 23256 14958
rect 23204 14894 23256 14900
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22836 12164 22888 12170
rect 22836 12106 22888 12112
rect 22848 11082 22876 12106
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22940 9194 22968 13398
rect 23124 12782 23152 14350
rect 23216 13530 23244 14894
rect 23400 14822 23428 17206
rect 23492 15162 23520 19858
rect 23676 19242 23704 26726
rect 23664 19236 23716 19242
rect 23664 19178 23716 19184
rect 23768 18850 23796 38270
rect 23848 38208 23900 38214
rect 23848 38150 23900 38156
rect 23860 28082 23888 38150
rect 23952 32910 23980 38270
rect 24124 38208 24176 38214
rect 24124 38150 24176 38156
rect 24136 37874 24164 38150
rect 24124 37868 24176 37874
rect 24124 37810 24176 37816
rect 24030 37768 24086 37777
rect 24030 37703 24086 37712
rect 24044 36242 24072 37703
rect 24032 36236 24084 36242
rect 24032 36178 24084 36184
rect 24032 35828 24084 35834
rect 24032 35770 24084 35776
rect 24044 35086 24072 35770
rect 24320 35630 24348 39986
rect 24308 35624 24360 35630
rect 24308 35566 24360 35572
rect 24122 35320 24178 35329
rect 24122 35255 24124 35264
rect 24176 35255 24178 35264
rect 24124 35226 24176 35232
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 24214 33824 24270 33833
rect 24214 33759 24270 33768
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 24032 32836 24084 32842
rect 24032 32778 24084 32784
rect 24044 32434 24072 32778
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 23940 31340 23992 31346
rect 23940 31282 23992 31288
rect 23952 30734 23980 31282
rect 24044 31226 24072 31962
rect 24124 31884 24176 31890
rect 24124 31826 24176 31832
rect 24136 31346 24164 31826
rect 24124 31340 24176 31346
rect 24124 31282 24176 31288
rect 24044 31198 24164 31226
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23860 24274 23888 25978
rect 23952 25294 23980 30670
rect 24044 28218 24072 31078
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 24044 26994 24072 28154
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 24044 25838 24072 26930
rect 24136 26042 24164 31198
rect 24228 27334 24256 33759
rect 24216 27328 24268 27334
rect 24216 27270 24268 27276
rect 24320 27146 24348 35566
rect 24228 27118 24348 27146
rect 24124 26036 24176 26042
rect 24124 25978 24176 25984
rect 24124 25900 24176 25906
rect 24124 25842 24176 25848
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 23940 24948 23992 24954
rect 23940 24890 23992 24896
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23952 24206 23980 24890
rect 24136 24410 24164 25842
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 23952 23610 23980 24142
rect 24124 23656 24176 23662
rect 23952 23582 24072 23610
rect 24124 23598 24176 23604
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23584 18822 23796 18850
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23388 14816 23440 14822
rect 23308 14764 23388 14770
rect 23308 14758 23440 14764
rect 23308 14742 23428 14758
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23216 13326 23244 13466
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23216 12782 23244 13262
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 23020 11076 23072 11082
rect 23020 11018 23072 11024
rect 22848 9178 22968 9194
rect 22836 9172 22968 9178
rect 22888 9166 22968 9172
rect 22836 9114 22888 9120
rect 23032 4622 23060 11018
rect 23124 10266 23152 12718
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23216 11150 23244 11494
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23216 10810 23244 11086
rect 23204 10804 23256 10810
rect 23204 10746 23256 10752
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23124 9382 23152 10202
rect 23216 10062 23244 10746
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23308 9518 23336 14742
rect 23492 14482 23520 15098
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23400 12782 23428 13874
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23124 8838 23152 9318
rect 23308 9178 23336 9454
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 23124 8090 23152 8774
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23400 7886 23428 12718
rect 23584 12238 23612 18822
rect 23860 18714 23888 23054
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23768 18686 23888 18714
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23676 17678 23704 18022
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23768 15026 23796 18686
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 18290 23888 18566
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 23860 17882 23888 18090
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23768 12850 23796 13670
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 9586 23888 10406
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23400 7002 23428 7822
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23952 5370 23980 22578
rect 24044 20058 24072 23582
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24136 19922 24164 23598
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 24228 19802 24256 27118
rect 24308 27056 24360 27062
rect 24308 26998 24360 27004
rect 24320 24818 24348 26998
rect 24412 26994 24440 51274
rect 24504 51270 24532 53926
rect 24596 51406 24624 54810
rect 24584 51400 24636 51406
rect 24582 51368 24584 51377
rect 24636 51368 24638 51377
rect 24582 51303 24638 51312
rect 24492 51264 24544 51270
rect 24492 51206 24544 51212
rect 24490 51096 24546 51105
rect 24688 51074 24716 60007
rect 24780 51270 24808 61254
rect 24860 61260 24912 61266
rect 24860 61202 24912 61208
rect 24860 61124 24912 61130
rect 24860 61066 24912 61072
rect 24768 51264 24820 51270
rect 24768 51206 24820 51212
rect 24490 51031 24546 51040
rect 24504 50930 24532 51031
rect 24642 51020 24716 51074
rect 24688 50946 24716 51020
rect 24872 50969 24900 61066
rect 24964 60722 24992 61542
rect 24952 60716 25004 60722
rect 24952 60658 25004 60664
rect 25056 60602 25084 61542
rect 24964 60574 25084 60602
rect 24964 56914 24992 60574
rect 25042 60480 25098 60489
rect 25042 60415 25098 60424
rect 24952 56908 25004 56914
rect 24952 56850 25004 56856
rect 24952 56772 25004 56778
rect 24952 56714 25004 56720
rect 24964 55418 24992 56714
rect 25056 56506 25084 60415
rect 25044 56500 25096 56506
rect 25044 56442 25096 56448
rect 25148 55865 25176 63838
rect 25240 62393 25268 64262
rect 25226 62384 25282 62393
rect 25226 62319 25282 62328
rect 25228 62280 25280 62286
rect 25228 62222 25280 62228
rect 25240 61810 25268 62222
rect 25228 61804 25280 61810
rect 25228 61746 25280 61752
rect 25240 61198 25268 61746
rect 25228 61192 25280 61198
rect 25228 61134 25280 61140
rect 25240 60722 25268 61134
rect 25332 61062 25360 67238
rect 25412 67244 25464 67250
rect 25412 67186 25464 67192
rect 25424 66570 25452 67186
rect 25516 67182 25544 69702
rect 25776 69116 26084 69136
rect 25776 69114 25782 69116
rect 25838 69114 25862 69116
rect 25918 69114 25942 69116
rect 25998 69114 26022 69116
rect 26078 69114 26084 69116
rect 25838 69062 25840 69114
rect 26020 69062 26022 69114
rect 25776 69060 25782 69062
rect 25838 69060 25862 69062
rect 25918 69060 25942 69062
rect 25998 69060 26022 69062
rect 26078 69060 26084 69062
rect 25776 69040 26084 69060
rect 25776 68028 26084 68048
rect 25776 68026 25782 68028
rect 25838 68026 25862 68028
rect 25918 68026 25942 68028
rect 25998 68026 26022 68028
rect 26078 68026 26084 68028
rect 25838 67974 25840 68026
rect 26020 67974 26022 68026
rect 25776 67972 25782 67974
rect 25838 67972 25862 67974
rect 25918 67972 25942 67974
rect 25998 67972 26022 67974
rect 26078 67972 26084 67974
rect 25776 67952 26084 67972
rect 26056 67856 26108 67862
rect 26054 67824 26056 67833
rect 26108 67824 26110 67833
rect 26054 67759 26110 67768
rect 25686 67688 25742 67697
rect 25686 67623 25742 67632
rect 25596 67584 25648 67590
rect 25596 67526 25648 67532
rect 25504 67176 25556 67182
rect 25504 67118 25556 67124
rect 25412 66564 25464 66570
rect 25412 66506 25464 66512
rect 25412 66156 25464 66162
rect 25412 66098 25464 66104
rect 25424 66065 25452 66098
rect 25410 66056 25466 66065
rect 25410 65991 25466 66000
rect 25504 65068 25556 65074
rect 25504 65010 25556 65016
rect 25516 64462 25544 65010
rect 25504 64456 25556 64462
rect 25504 64398 25556 64404
rect 25504 64116 25556 64122
rect 25504 64058 25556 64064
rect 25412 63912 25464 63918
rect 25412 63854 25464 63860
rect 25424 63374 25452 63854
rect 25412 63368 25464 63374
rect 25412 63310 25464 63316
rect 25412 63232 25464 63238
rect 25412 63174 25464 63180
rect 25424 61606 25452 63174
rect 25412 61600 25464 61606
rect 25412 61542 25464 61548
rect 25412 61396 25464 61402
rect 25412 61338 25464 61344
rect 25320 61056 25372 61062
rect 25320 60998 25372 61004
rect 25318 60888 25374 60897
rect 25318 60823 25374 60832
rect 25332 60722 25360 60823
rect 25228 60716 25280 60722
rect 25228 60658 25280 60664
rect 25320 60716 25372 60722
rect 25320 60658 25372 60664
rect 25240 59702 25268 60658
rect 25320 60308 25372 60314
rect 25320 60250 25372 60256
rect 25228 59696 25280 59702
rect 25228 59638 25280 59644
rect 25228 59492 25280 59498
rect 25228 59434 25280 59440
rect 25240 56846 25268 59434
rect 25228 56840 25280 56846
rect 25228 56782 25280 56788
rect 25228 56704 25280 56710
rect 25226 56672 25228 56681
rect 25280 56672 25282 56681
rect 25226 56607 25282 56616
rect 25134 55856 25190 55865
rect 25134 55791 25190 55800
rect 25332 55706 25360 60250
rect 25424 57594 25452 61338
rect 25516 61062 25544 64058
rect 25608 61130 25636 67526
rect 25700 64122 25728 67623
rect 26160 67590 26188 73034
rect 26252 67930 26280 74190
rect 26240 67924 26292 67930
rect 26240 67866 26292 67872
rect 26148 67584 26200 67590
rect 26148 67526 26200 67532
rect 26160 67368 26188 67526
rect 26068 67340 26188 67368
rect 26068 67250 26096 67340
rect 26160 67250 26280 67266
rect 26056 67244 26108 67250
rect 26056 67186 26108 67192
rect 26160 67244 26292 67250
rect 26160 67238 26240 67244
rect 25776 66940 26084 66960
rect 25776 66938 25782 66940
rect 25838 66938 25862 66940
rect 25918 66938 25942 66940
rect 25998 66938 26022 66940
rect 26078 66938 26084 66940
rect 25838 66886 25840 66938
rect 26020 66886 26022 66938
rect 25776 66884 25782 66886
rect 25838 66884 25862 66886
rect 25918 66884 25942 66886
rect 25998 66884 26022 66886
rect 26078 66884 26084 66886
rect 25776 66864 26084 66884
rect 26160 66638 26188 67238
rect 26240 67186 26292 67192
rect 26238 67144 26294 67153
rect 26238 67079 26294 67088
rect 26148 66632 26200 66638
rect 26148 66574 26200 66580
rect 26148 66156 26200 66162
rect 26148 66098 26200 66104
rect 25776 65852 26084 65872
rect 25776 65850 25782 65852
rect 25838 65850 25862 65852
rect 25918 65850 25942 65852
rect 25998 65850 26022 65852
rect 26078 65850 26084 65852
rect 25838 65798 25840 65850
rect 26020 65798 26022 65850
rect 25776 65796 25782 65798
rect 25838 65796 25862 65798
rect 25918 65796 25942 65798
rect 25998 65796 26022 65798
rect 26078 65796 26084 65798
rect 25776 65776 26084 65796
rect 26160 64938 26188 66098
rect 26148 64932 26200 64938
rect 26148 64874 26200 64880
rect 25776 64764 26084 64784
rect 25776 64762 25782 64764
rect 25838 64762 25862 64764
rect 25918 64762 25942 64764
rect 25998 64762 26022 64764
rect 26078 64762 26084 64764
rect 25838 64710 25840 64762
rect 26020 64710 26022 64762
rect 25776 64708 25782 64710
rect 25838 64708 25862 64710
rect 25918 64708 25942 64710
rect 25998 64708 26022 64710
rect 26078 64708 26084 64710
rect 25776 64688 26084 64708
rect 26160 64462 26188 64874
rect 26148 64456 26200 64462
rect 26148 64398 26200 64404
rect 25688 64116 25740 64122
rect 25688 64058 25740 64064
rect 25688 63912 25740 63918
rect 25688 63854 25740 63860
rect 25700 61946 25728 63854
rect 25776 63676 26084 63696
rect 25776 63674 25782 63676
rect 25838 63674 25862 63676
rect 25918 63674 25942 63676
rect 25998 63674 26022 63676
rect 26078 63674 26084 63676
rect 25838 63622 25840 63674
rect 26020 63622 26022 63674
rect 25776 63620 25782 63622
rect 25838 63620 25862 63622
rect 25918 63620 25942 63622
rect 25998 63620 26022 63622
rect 26078 63620 26084 63622
rect 25776 63600 26084 63620
rect 26160 63238 26188 64398
rect 26148 63232 26200 63238
rect 26148 63174 26200 63180
rect 25776 62588 26084 62608
rect 25776 62586 25782 62588
rect 25838 62586 25862 62588
rect 25918 62586 25942 62588
rect 25998 62586 26022 62588
rect 26078 62586 26084 62588
rect 25838 62534 25840 62586
rect 26020 62534 26022 62586
rect 25776 62532 25782 62534
rect 25838 62532 25862 62534
rect 25918 62532 25942 62534
rect 25998 62532 26022 62534
rect 26078 62532 26084 62534
rect 25776 62512 26084 62532
rect 26148 62348 26200 62354
rect 26148 62290 26200 62296
rect 25964 62144 26016 62150
rect 25964 62086 26016 62092
rect 25688 61940 25740 61946
rect 25688 61882 25740 61888
rect 25976 61878 26004 62086
rect 25964 61872 26016 61878
rect 25964 61814 26016 61820
rect 25688 61804 25740 61810
rect 25688 61746 25740 61752
rect 25700 61198 25728 61746
rect 25776 61500 26084 61520
rect 25776 61498 25782 61500
rect 25838 61498 25862 61500
rect 25918 61498 25942 61500
rect 25998 61498 26022 61500
rect 26078 61498 26084 61500
rect 25838 61446 25840 61498
rect 26020 61446 26022 61498
rect 25776 61444 25782 61446
rect 25838 61444 25862 61446
rect 25918 61444 25942 61446
rect 25998 61444 26022 61446
rect 26078 61444 26084 61446
rect 25776 61424 26084 61444
rect 25688 61192 25740 61198
rect 25964 61192 26016 61198
rect 25688 61134 25740 61140
rect 25778 61160 25834 61169
rect 25596 61124 25648 61130
rect 25964 61134 26016 61140
rect 25778 61095 25780 61104
rect 25596 61066 25648 61072
rect 25832 61095 25834 61104
rect 25780 61066 25832 61072
rect 25504 61056 25556 61062
rect 25504 60998 25556 61004
rect 25688 61056 25740 61062
rect 25688 60998 25740 61004
rect 25594 60888 25650 60897
rect 25594 60823 25650 60832
rect 25504 60648 25556 60654
rect 25504 60590 25556 60596
rect 25412 57588 25464 57594
rect 25412 57530 25464 57536
rect 25412 56500 25464 56506
rect 25412 56442 25464 56448
rect 25148 55678 25360 55706
rect 25044 55616 25096 55622
rect 25044 55558 25096 55564
rect 25056 55457 25084 55558
rect 25042 55448 25098 55457
rect 24952 55412 25004 55418
rect 25042 55383 25098 55392
rect 24952 55354 25004 55360
rect 25044 55208 25096 55214
rect 24950 55176 25006 55185
rect 25044 55150 25096 55156
rect 24950 55111 25006 55120
rect 24964 51649 24992 55111
rect 25056 54913 25084 55150
rect 25042 54904 25098 54913
rect 25042 54839 25098 54848
rect 25044 54120 25096 54126
rect 25044 54062 25096 54068
rect 24950 51640 25006 51649
rect 24950 51575 25006 51584
rect 24952 51332 25004 51338
rect 24952 51274 25004 51280
rect 24858 50960 24914 50969
rect 24492 50924 24544 50930
rect 24688 50918 24808 50946
rect 24492 50866 24544 50872
rect 24504 49774 24532 50866
rect 24780 50674 24808 50918
rect 24858 50895 24914 50904
rect 24860 50856 24912 50862
rect 24860 50798 24912 50804
rect 24872 50697 24900 50798
rect 24964 50794 24992 51274
rect 24952 50788 25004 50794
rect 24952 50730 25004 50736
rect 24688 50646 24808 50674
rect 24858 50688 24914 50697
rect 24584 50448 24636 50454
rect 24584 50390 24636 50396
rect 24596 49842 24624 50390
rect 24688 50318 24716 50646
rect 24914 50646 24992 50674
rect 24858 50623 24914 50632
rect 24858 50552 24914 50561
rect 24768 50516 24820 50522
rect 24858 50487 24914 50496
rect 24768 50458 24820 50464
rect 24676 50312 24728 50318
rect 24676 50254 24728 50260
rect 24780 50164 24808 50458
rect 24688 50136 24808 50164
rect 24584 49836 24636 49842
rect 24584 49778 24636 49784
rect 24492 49768 24544 49774
rect 24492 49710 24544 49716
rect 24504 48890 24532 49710
rect 24596 48890 24624 49778
rect 24492 48884 24544 48890
rect 24492 48826 24544 48832
rect 24584 48884 24636 48890
rect 24584 48826 24636 48832
rect 24490 48784 24546 48793
rect 24490 48719 24546 48728
rect 24504 45014 24532 48719
rect 24582 48512 24638 48521
rect 24582 48447 24638 48456
rect 24492 45008 24544 45014
rect 24492 44950 24544 44956
rect 24492 44872 24544 44878
rect 24492 44814 24544 44820
rect 24504 44538 24532 44814
rect 24492 44532 24544 44538
rect 24492 44474 24544 44480
rect 24492 44260 24544 44266
rect 24492 44202 24544 44208
rect 24504 44033 24532 44202
rect 24490 44024 24546 44033
rect 24490 43959 24546 43968
rect 24492 43852 24544 43858
rect 24492 43794 24544 43800
rect 24504 43246 24532 43794
rect 24596 43450 24624 48447
rect 24688 45626 24716 50136
rect 24766 50008 24822 50017
rect 24766 49943 24768 49952
rect 24820 49943 24822 49952
rect 24768 49914 24820 49920
rect 24768 49836 24820 49842
rect 24768 49778 24820 49784
rect 24780 49706 24808 49778
rect 24768 49700 24820 49706
rect 24768 49642 24820 49648
rect 24768 48748 24820 48754
rect 24768 48690 24820 48696
rect 24780 47190 24808 48690
rect 24768 47184 24820 47190
rect 24768 47126 24820 47132
rect 24768 46980 24820 46986
rect 24768 46922 24820 46928
rect 24676 45620 24728 45626
rect 24676 45562 24728 45568
rect 24780 45558 24808 46922
rect 24768 45552 24820 45558
rect 24768 45494 24820 45500
rect 24768 45416 24820 45422
rect 24768 45358 24820 45364
rect 24676 45280 24728 45286
rect 24676 45222 24728 45228
rect 24688 45121 24716 45222
rect 24674 45112 24730 45121
rect 24674 45047 24730 45056
rect 24780 44810 24808 45358
rect 24768 44804 24820 44810
rect 24768 44746 24820 44752
rect 24676 44464 24728 44470
rect 24676 44406 24728 44412
rect 24688 43858 24716 44406
rect 24676 43852 24728 43858
rect 24676 43794 24728 43800
rect 24584 43444 24636 43450
rect 24584 43386 24636 43392
rect 24492 43240 24544 43246
rect 24492 43182 24544 43188
rect 24504 43081 24532 43182
rect 24584 43172 24636 43178
rect 24584 43114 24636 43120
rect 24490 43072 24546 43081
rect 24490 43007 24546 43016
rect 24492 42764 24544 42770
rect 24492 42706 24544 42712
rect 24504 39574 24532 42706
rect 24596 39846 24624 43114
rect 24688 42906 24716 43794
rect 24780 43790 24808 44746
rect 24768 43784 24820 43790
rect 24768 43726 24820 43732
rect 24780 43314 24808 43726
rect 24768 43308 24820 43314
rect 24768 43250 24820 43256
rect 24766 43208 24822 43217
rect 24766 43143 24822 43152
rect 24780 43110 24808 43143
rect 24768 43104 24820 43110
rect 24768 43046 24820 43052
rect 24766 42936 24822 42945
rect 24676 42900 24728 42906
rect 24766 42871 24822 42880
rect 24676 42842 24728 42848
rect 24780 42838 24808 42871
rect 24768 42832 24820 42838
rect 24768 42774 24820 42780
rect 24674 42664 24730 42673
rect 24674 42599 24730 42608
rect 24688 42566 24716 42599
rect 24676 42560 24728 42566
rect 24676 42502 24728 42508
rect 24780 42208 24808 42774
rect 24872 42673 24900 50487
rect 24964 50454 24992 50646
rect 24952 50448 25004 50454
rect 24952 50390 25004 50396
rect 24950 49736 25006 49745
rect 24950 49671 25006 49680
rect 24964 46714 24992 49671
rect 24952 46708 25004 46714
rect 24952 46650 25004 46656
rect 25056 46152 25084 54062
rect 25148 51218 25176 55678
rect 25320 55616 25372 55622
rect 25320 55558 25372 55564
rect 25332 55214 25360 55558
rect 25424 55350 25452 56442
rect 25516 55865 25544 60590
rect 25608 57050 25636 60823
rect 25596 57044 25648 57050
rect 25596 56986 25648 56992
rect 25596 56908 25648 56914
rect 25596 56850 25648 56856
rect 25502 55856 25558 55865
rect 25502 55791 25558 55800
rect 25504 55684 25556 55690
rect 25504 55626 25556 55632
rect 25412 55344 25464 55350
rect 25412 55286 25464 55292
rect 25320 55208 25372 55214
rect 25320 55150 25372 55156
rect 25228 55140 25280 55146
rect 25228 55082 25280 55088
rect 25240 54194 25268 55082
rect 25332 55078 25360 55150
rect 25320 55072 25372 55078
rect 25320 55014 25372 55020
rect 25320 54324 25372 54330
rect 25320 54266 25372 54272
rect 25228 54188 25280 54194
rect 25228 54130 25280 54136
rect 25240 54097 25268 54130
rect 25226 54088 25282 54097
rect 25226 54023 25282 54032
rect 25332 53174 25360 54266
rect 25320 53168 25372 53174
rect 25320 53110 25372 53116
rect 25332 51542 25360 53110
rect 25412 51876 25464 51882
rect 25412 51818 25464 51824
rect 25320 51536 25372 51542
rect 25320 51478 25372 51484
rect 25320 51400 25372 51406
rect 25320 51342 25372 51348
rect 25148 51190 25268 51218
rect 25134 51096 25190 51105
rect 25134 51031 25190 51040
rect 24964 46124 25084 46152
rect 24964 45558 24992 46124
rect 25044 46028 25096 46034
rect 25044 45970 25096 45976
rect 24952 45552 25004 45558
rect 24952 45494 25004 45500
rect 25056 45422 25084 45970
rect 25044 45416 25096 45422
rect 25044 45358 25096 45364
rect 24952 45280 25004 45286
rect 24952 45222 25004 45228
rect 24858 42664 24914 42673
rect 24858 42599 24914 42608
rect 24688 42180 24808 42208
rect 24688 42022 24716 42180
rect 24768 42084 24820 42090
rect 24768 42026 24820 42032
rect 24676 42016 24728 42022
rect 24676 41958 24728 41964
rect 24780 41614 24808 42026
rect 24768 41608 24820 41614
rect 24768 41550 24820 41556
rect 24860 41472 24912 41478
rect 24860 41414 24912 41420
rect 24766 41304 24822 41313
rect 24766 41239 24822 41248
rect 24780 41070 24808 41239
rect 24768 41064 24820 41070
rect 24768 41006 24820 41012
rect 24676 40996 24728 41002
rect 24676 40938 24728 40944
rect 24688 39846 24716 40938
rect 24780 39914 24808 41006
rect 24768 39908 24820 39914
rect 24768 39850 24820 39856
rect 24584 39840 24636 39846
rect 24584 39782 24636 39788
rect 24676 39840 24728 39846
rect 24676 39782 24728 39788
rect 24492 39568 24544 39574
rect 24492 39510 24544 39516
rect 24584 39432 24636 39438
rect 24584 39374 24636 39380
rect 24596 38962 24624 39374
rect 24768 39364 24820 39370
rect 24768 39306 24820 39312
rect 24676 39296 24728 39302
rect 24676 39238 24728 39244
rect 24584 38956 24636 38962
rect 24584 38898 24636 38904
rect 24596 38865 24624 38898
rect 24582 38856 24638 38865
rect 24582 38791 24638 38800
rect 24688 38677 24716 39238
rect 24780 39098 24808 39306
rect 24768 39092 24820 39098
rect 24768 39034 24820 39040
rect 24674 38668 24730 38677
rect 24674 38603 24730 38612
rect 24582 38448 24638 38457
rect 24582 38383 24638 38392
rect 24596 37942 24624 38383
rect 24674 38312 24730 38321
rect 24674 38247 24730 38256
rect 24584 37936 24636 37942
rect 24584 37878 24636 37884
rect 24492 37732 24544 37738
rect 24492 37674 24544 37680
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24400 25764 24452 25770
rect 24400 25706 24452 25712
rect 24412 25498 24440 25706
rect 24400 25492 24452 25498
rect 24400 25434 24452 25440
rect 24400 25356 24452 25362
rect 24400 25298 24452 25304
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24412 24750 24440 25298
rect 24400 24744 24452 24750
rect 24306 24712 24362 24721
rect 24400 24686 24452 24692
rect 24306 24647 24362 24656
rect 24320 22642 24348 24647
rect 24308 22636 24360 22642
rect 24308 22578 24360 22584
rect 24412 22094 24440 24686
rect 24136 19774 24256 19802
rect 24320 22066 24440 22094
rect 24032 19236 24084 19242
rect 24032 19178 24084 19184
rect 24044 18290 24072 19178
rect 24136 18358 24164 19774
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24228 19514 24256 19654
rect 24216 19508 24268 19514
rect 24216 19450 24268 19456
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24044 17882 24072 18226
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24044 16998 24072 17818
rect 24228 17202 24256 18022
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 24044 14822 24072 14962
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24136 13938 24164 17070
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24136 13394 24164 13874
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24228 13190 24256 15370
rect 24320 15314 24348 22066
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21418 24440 21830
rect 24400 21412 24452 21418
rect 24400 21354 24452 21360
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24412 19378 24440 19654
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24504 15502 24532 37674
rect 24596 37330 24624 37878
rect 24584 37324 24636 37330
rect 24584 37266 24636 37272
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24596 27470 24624 37062
rect 24688 33522 24716 38247
rect 24780 37670 24808 39034
rect 24872 38677 24900 41414
rect 24964 38962 24992 45222
rect 25056 44946 25084 45358
rect 25044 44940 25096 44946
rect 25044 44882 25096 44888
rect 25148 44742 25176 51031
rect 25240 50522 25268 51190
rect 25228 50516 25280 50522
rect 25228 50458 25280 50464
rect 25228 50244 25280 50250
rect 25228 50186 25280 50192
rect 25240 49910 25268 50186
rect 25228 49904 25280 49910
rect 25228 49846 25280 49852
rect 25228 49632 25280 49638
rect 25228 49574 25280 49580
rect 25240 49366 25268 49574
rect 25228 49360 25280 49366
rect 25228 49302 25280 49308
rect 25228 49224 25280 49230
rect 25228 49166 25280 49172
rect 25240 48754 25268 49166
rect 25228 48748 25280 48754
rect 25228 48690 25280 48696
rect 25240 48074 25268 48690
rect 25332 48278 25360 51342
rect 25320 48272 25372 48278
rect 25320 48214 25372 48220
rect 25320 48136 25372 48142
rect 25320 48078 25372 48084
rect 25228 48068 25280 48074
rect 25228 48010 25280 48016
rect 25228 47592 25280 47598
rect 25228 47534 25280 47540
rect 25240 46209 25268 47534
rect 25226 46200 25282 46209
rect 25226 46135 25282 46144
rect 25228 46096 25280 46102
rect 25228 46038 25280 46044
rect 25044 44736 25096 44742
rect 25044 44678 25096 44684
rect 25136 44736 25188 44742
rect 25136 44678 25188 44684
rect 24952 38956 25004 38962
rect 24952 38898 25004 38904
rect 24952 38820 25004 38826
rect 24952 38762 25004 38768
rect 24858 38668 24914 38677
rect 24858 38603 24914 38612
rect 24964 38570 24992 38762
rect 24872 38542 24992 38570
rect 24872 38468 24900 38542
rect 24872 38440 24992 38468
rect 24858 38176 24914 38185
rect 24858 38111 24914 38120
rect 24872 37942 24900 38111
rect 24872 37936 24930 37942
rect 24872 37913 24878 37936
rect 24858 37904 24878 37913
rect 24914 37878 24930 37884
rect 24858 37839 24914 37848
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 24858 37632 24914 37641
rect 24780 37398 24808 37606
rect 24858 37567 24914 37576
rect 24768 37392 24820 37398
rect 24768 37334 24820 37340
rect 24768 36712 24820 36718
rect 24768 36654 24820 36660
rect 24780 36310 24808 36654
rect 24768 36304 24820 36310
rect 24768 36246 24820 36252
rect 24768 36168 24820 36174
rect 24766 36136 24768 36145
rect 24820 36136 24822 36145
rect 24766 36071 24822 36080
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 24780 35698 24808 35770
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 24768 35216 24820 35222
rect 24768 35158 24820 35164
rect 24780 34406 24808 35158
rect 24768 34400 24820 34406
rect 24768 34342 24820 34348
rect 24872 34218 24900 37567
rect 24964 36174 24992 38440
rect 25056 37874 25084 44678
rect 25136 43648 25188 43654
rect 25136 43590 25188 43596
rect 25148 43382 25176 43590
rect 25136 43376 25188 43382
rect 25136 43318 25188 43324
rect 25148 43178 25176 43318
rect 25136 43172 25188 43178
rect 25136 43114 25188 43120
rect 25134 43072 25190 43081
rect 25134 43007 25190 43016
rect 25148 42838 25176 43007
rect 25136 42832 25188 42838
rect 25136 42774 25188 42780
rect 25136 42696 25188 42702
rect 25136 42638 25188 42644
rect 25148 41546 25176 42638
rect 25136 41540 25188 41546
rect 25136 41482 25188 41488
rect 25136 40996 25188 41002
rect 25136 40938 25188 40944
rect 25148 40497 25176 40938
rect 25240 40905 25268 46038
rect 25332 45830 25360 48078
rect 25424 46102 25452 51818
rect 25516 51218 25544 55626
rect 25608 52018 25636 56850
rect 25700 56506 25728 60998
rect 25872 60852 25924 60858
rect 25872 60794 25924 60800
rect 25884 60761 25912 60794
rect 25870 60752 25926 60761
rect 25780 60722 25832 60728
rect 25870 60687 25926 60696
rect 25780 60664 25832 60670
rect 25792 60636 25820 60664
rect 25792 60608 25912 60636
rect 25976 60625 26004 61134
rect 26160 60704 26188 62290
rect 26252 61169 26280 67079
rect 26344 64666 26372 76366
rect 27172 74534 27200 77386
rect 26988 74506 27200 74534
rect 26792 73160 26844 73166
rect 26792 73102 26844 73108
rect 26424 68332 26476 68338
rect 26424 68274 26476 68280
rect 26332 64660 26384 64666
rect 26332 64602 26384 64608
rect 26332 64456 26384 64462
rect 26330 64424 26332 64433
rect 26384 64424 26386 64433
rect 26330 64359 26386 64368
rect 26436 62150 26464 68274
rect 26516 68196 26568 68202
rect 26516 68138 26568 68144
rect 26528 66774 26556 68138
rect 26608 67856 26660 67862
rect 26608 67798 26660 67804
rect 26516 66768 26568 66774
rect 26516 66710 26568 66716
rect 26516 64388 26568 64394
rect 26516 64330 26568 64336
rect 26528 63073 26556 64330
rect 26514 63064 26570 63073
rect 26514 62999 26570 63008
rect 26516 62824 26568 62830
rect 26516 62766 26568 62772
rect 26424 62144 26476 62150
rect 26424 62086 26476 62092
rect 26332 61804 26384 61810
rect 26332 61746 26384 61752
rect 26344 61198 26372 61746
rect 26332 61192 26384 61198
rect 26238 61160 26294 61169
rect 26332 61134 26384 61140
rect 26238 61095 26294 61104
rect 26240 61056 26292 61062
rect 26240 60998 26292 61004
rect 26068 60676 26188 60704
rect 25884 60500 25912 60608
rect 25962 60616 26018 60625
rect 25962 60551 26018 60560
rect 26068 60500 26096 60676
rect 26148 60580 26200 60586
rect 26148 60522 26200 60528
rect 25884 60472 26096 60500
rect 25776 60412 26084 60432
rect 25776 60410 25782 60412
rect 25838 60410 25862 60412
rect 25918 60410 25942 60412
rect 25998 60410 26022 60412
rect 26078 60410 26084 60412
rect 25838 60358 25840 60410
rect 26020 60358 26022 60410
rect 25776 60356 25782 60358
rect 25838 60356 25862 60358
rect 25918 60356 25942 60358
rect 25998 60356 26022 60358
rect 26078 60356 26084 60358
rect 25776 60336 26084 60356
rect 26160 60296 26188 60522
rect 26068 60268 26188 60296
rect 25778 60208 25834 60217
rect 25778 60143 25834 60152
rect 25872 60172 25924 60178
rect 25792 60110 25820 60143
rect 25872 60114 25924 60120
rect 25780 60104 25832 60110
rect 25780 60046 25832 60052
rect 25792 59498 25820 60046
rect 25884 59945 25912 60114
rect 25870 59936 25926 59945
rect 25870 59871 25926 59880
rect 25872 59764 25924 59770
rect 25872 59706 25924 59712
rect 25884 59673 25912 59706
rect 26068 59673 26096 60268
rect 26146 60208 26202 60217
rect 26146 60143 26202 60152
rect 25870 59664 25926 59673
rect 25870 59599 25926 59608
rect 26054 59664 26110 59673
rect 26054 59599 26110 59608
rect 25780 59492 25832 59498
rect 25780 59434 25832 59440
rect 25776 59324 26084 59344
rect 25776 59322 25782 59324
rect 25838 59322 25862 59324
rect 25918 59322 25942 59324
rect 25998 59322 26022 59324
rect 26078 59322 26084 59324
rect 25838 59270 25840 59322
rect 26020 59270 26022 59322
rect 25776 59268 25782 59270
rect 25838 59268 25862 59270
rect 25918 59268 25942 59270
rect 25998 59268 26022 59270
rect 26078 59268 26084 59270
rect 25776 59248 26084 59268
rect 25776 58236 26084 58256
rect 25776 58234 25782 58236
rect 25838 58234 25862 58236
rect 25918 58234 25942 58236
rect 25998 58234 26022 58236
rect 26078 58234 26084 58236
rect 25838 58182 25840 58234
rect 26020 58182 26022 58234
rect 25776 58180 25782 58182
rect 25838 58180 25862 58182
rect 25918 58180 25942 58182
rect 25998 58180 26022 58182
rect 26078 58180 26084 58182
rect 25776 58160 26084 58180
rect 25872 58064 25924 58070
rect 25872 58006 25924 58012
rect 25962 58032 26018 58041
rect 25884 57390 25912 58006
rect 25962 57967 26018 57976
rect 25872 57384 25924 57390
rect 25976 57361 26004 57967
rect 26054 57488 26110 57497
rect 26054 57423 26056 57432
rect 26108 57423 26110 57432
rect 26056 57394 26108 57400
rect 25872 57326 25924 57332
rect 25962 57352 26018 57361
rect 25962 57287 26018 57296
rect 25776 57148 26084 57168
rect 25776 57146 25782 57148
rect 25838 57146 25862 57148
rect 25918 57146 25942 57148
rect 25998 57146 26022 57148
rect 26078 57146 26084 57148
rect 25838 57094 25840 57146
rect 26020 57094 26022 57146
rect 25776 57092 25782 57094
rect 25838 57092 25862 57094
rect 25918 57092 25942 57094
rect 25998 57092 26022 57094
rect 26078 57092 26084 57094
rect 25776 57072 26084 57092
rect 26054 56944 26110 56953
rect 26054 56879 26110 56888
rect 25964 56840 26016 56846
rect 25964 56782 26016 56788
rect 25872 56704 25924 56710
rect 25872 56646 25924 56652
rect 25884 56506 25912 56646
rect 25688 56500 25740 56506
rect 25688 56442 25740 56448
rect 25872 56500 25924 56506
rect 25872 56442 25924 56448
rect 25976 56370 26004 56782
rect 26068 56710 26096 56879
rect 26056 56704 26108 56710
rect 26056 56646 26108 56652
rect 25964 56364 26016 56370
rect 25964 56306 26016 56312
rect 25776 56060 26084 56080
rect 25776 56058 25782 56060
rect 25838 56058 25862 56060
rect 25918 56058 25942 56060
rect 25998 56058 26022 56060
rect 26078 56058 26084 56060
rect 25838 56006 25840 56058
rect 26020 56006 26022 56058
rect 25776 56004 25782 56006
rect 25838 56004 25862 56006
rect 25918 56004 25942 56006
rect 25998 56004 26022 56006
rect 26078 56004 26084 56006
rect 25776 55984 26084 56004
rect 25688 55956 25740 55962
rect 25688 55898 25740 55904
rect 25700 55690 25728 55898
rect 25962 55856 26018 55865
rect 25962 55791 25964 55800
rect 26016 55791 26018 55800
rect 25964 55762 26016 55768
rect 25688 55684 25740 55690
rect 25688 55626 25740 55632
rect 25964 55684 26016 55690
rect 25964 55626 26016 55632
rect 25870 55448 25926 55457
rect 25780 55412 25832 55418
rect 25870 55383 25926 55392
rect 25780 55354 25832 55360
rect 25792 55321 25820 55354
rect 25884 55350 25912 55383
rect 25872 55344 25924 55350
rect 25778 55312 25834 55321
rect 25872 55286 25924 55292
rect 25778 55247 25834 55256
rect 25976 55185 26004 55626
rect 25962 55176 26018 55185
rect 25962 55111 26018 55120
rect 25776 54972 26084 54992
rect 25776 54970 25782 54972
rect 25838 54970 25862 54972
rect 25918 54970 25942 54972
rect 25998 54970 26022 54972
rect 26078 54970 26084 54972
rect 25838 54918 25840 54970
rect 26020 54918 26022 54970
rect 25776 54916 25782 54918
rect 25838 54916 25862 54918
rect 25918 54916 25942 54918
rect 25998 54916 26022 54918
rect 26078 54916 26084 54918
rect 25776 54896 26084 54916
rect 26160 54874 26188 60143
rect 26252 56930 26280 60998
rect 26344 60586 26372 61134
rect 26422 61024 26478 61033
rect 26422 60959 26478 60968
rect 26332 60580 26384 60586
rect 26332 60522 26384 60528
rect 26344 60110 26372 60522
rect 26332 60104 26384 60110
rect 26332 60046 26384 60052
rect 26332 59628 26384 59634
rect 26332 59570 26384 59576
rect 26344 58614 26372 59570
rect 26332 58608 26384 58614
rect 26330 58576 26332 58585
rect 26384 58576 26386 58585
rect 26330 58511 26386 58520
rect 26332 58404 26384 58410
rect 26332 58346 26384 58352
rect 26344 57633 26372 58346
rect 26330 57624 26386 57633
rect 26330 57559 26386 57568
rect 26332 57452 26384 57458
rect 26332 57394 26384 57400
rect 26344 57050 26372 57394
rect 26332 57044 26384 57050
rect 26332 56986 26384 56992
rect 26252 56902 26372 56930
rect 26240 56840 26292 56846
rect 26240 56782 26292 56788
rect 26252 56370 26280 56782
rect 26240 56364 26292 56370
rect 26240 56306 26292 56312
rect 26252 55078 26280 56306
rect 26240 55072 26292 55078
rect 26240 55014 26292 55020
rect 26148 54868 26200 54874
rect 26148 54810 26200 54816
rect 26056 54800 26108 54806
rect 26056 54742 26108 54748
rect 26146 54768 26202 54777
rect 26068 54233 26096 54742
rect 26146 54703 26202 54712
rect 26160 54534 26188 54703
rect 26252 54670 26280 55014
rect 26240 54664 26292 54670
rect 26240 54606 26292 54612
rect 26148 54528 26200 54534
rect 26148 54470 26200 54476
rect 26146 54360 26202 54369
rect 26146 54295 26202 54304
rect 26054 54224 26110 54233
rect 26054 54159 26110 54168
rect 25776 53884 26084 53904
rect 25776 53882 25782 53884
rect 25838 53882 25862 53884
rect 25918 53882 25942 53884
rect 25998 53882 26022 53884
rect 26078 53882 26084 53884
rect 25838 53830 25840 53882
rect 26020 53830 26022 53882
rect 25776 53828 25782 53830
rect 25838 53828 25862 53830
rect 25918 53828 25942 53830
rect 25998 53828 26022 53830
rect 26078 53828 26084 53830
rect 25776 53808 26084 53828
rect 25872 53644 25924 53650
rect 25872 53586 25924 53592
rect 25884 52970 25912 53586
rect 26160 53582 26188 54295
rect 26148 53576 26200 53582
rect 26148 53518 26200 53524
rect 25964 53440 26016 53446
rect 25964 53382 26016 53388
rect 25976 53145 26004 53382
rect 25962 53136 26018 53145
rect 26160 53106 26188 53518
rect 25962 53071 26018 53080
rect 26148 53100 26200 53106
rect 26148 53042 26200 53048
rect 25872 52964 25924 52970
rect 25872 52906 25924 52912
rect 25776 52796 26084 52816
rect 25776 52794 25782 52796
rect 25838 52794 25862 52796
rect 25918 52794 25942 52796
rect 25998 52794 26022 52796
rect 26078 52794 26084 52796
rect 25838 52742 25840 52794
rect 26020 52742 26022 52794
rect 25776 52740 25782 52742
rect 25838 52740 25862 52742
rect 25918 52740 25942 52742
rect 25998 52740 26022 52742
rect 26078 52740 26084 52742
rect 25776 52720 26084 52740
rect 26160 52494 26188 53042
rect 26148 52488 26200 52494
rect 26148 52430 26200 52436
rect 25964 52352 26016 52358
rect 25964 52294 26016 52300
rect 25976 52154 26004 52294
rect 25964 52148 26016 52154
rect 25964 52090 26016 52096
rect 25688 52080 25740 52086
rect 25688 52022 25740 52028
rect 25596 52012 25648 52018
rect 25596 51954 25648 51960
rect 25608 51338 25636 51954
rect 25596 51332 25648 51338
rect 25596 51274 25648 51280
rect 25516 51190 25636 51218
rect 25504 50924 25556 50930
rect 25504 50866 25556 50872
rect 25516 49434 25544 50866
rect 25504 49428 25556 49434
rect 25504 49370 25556 49376
rect 25504 49088 25556 49094
rect 25504 49030 25556 49036
rect 25516 48929 25544 49030
rect 25502 48920 25558 48929
rect 25502 48855 25558 48864
rect 25504 48816 25556 48822
rect 25504 48758 25556 48764
rect 25516 47462 25544 48758
rect 25504 47456 25556 47462
rect 25504 47398 25556 47404
rect 25504 46504 25556 46510
rect 25502 46472 25504 46481
rect 25556 46472 25558 46481
rect 25502 46407 25558 46416
rect 25504 46368 25556 46374
rect 25504 46310 25556 46316
rect 25412 46096 25464 46102
rect 25412 46038 25464 46044
rect 25412 45892 25464 45898
rect 25516 45880 25544 46310
rect 25464 45852 25544 45880
rect 25412 45834 25464 45840
rect 25320 45824 25372 45830
rect 25320 45766 25372 45772
rect 25320 45620 25372 45626
rect 25320 45562 25372 45568
rect 25332 45422 25360 45562
rect 25320 45416 25372 45422
rect 25320 45358 25372 45364
rect 25332 44946 25360 45358
rect 25320 44940 25372 44946
rect 25320 44882 25372 44888
rect 25332 44334 25360 44882
rect 25320 44328 25372 44334
rect 25320 44270 25372 44276
rect 25332 43314 25360 44270
rect 25320 43308 25372 43314
rect 25320 43250 25372 43256
rect 25320 43172 25372 43178
rect 25320 43114 25372 43120
rect 25332 42566 25360 43114
rect 25320 42560 25372 42566
rect 25320 42502 25372 42508
rect 25332 42401 25360 42502
rect 25318 42392 25374 42401
rect 25318 42327 25374 42336
rect 25424 42226 25452 45834
rect 25504 45552 25556 45558
rect 25504 45494 25556 45500
rect 25516 44402 25544 45494
rect 25504 44396 25556 44402
rect 25504 44338 25556 44344
rect 25412 42220 25464 42226
rect 25412 42162 25464 42168
rect 25320 42016 25372 42022
rect 25320 41958 25372 41964
rect 25332 41682 25360 41958
rect 25320 41676 25372 41682
rect 25320 41618 25372 41624
rect 25318 41576 25374 41585
rect 25318 41511 25374 41520
rect 25226 40896 25282 40905
rect 25226 40831 25282 40840
rect 25226 40760 25282 40769
rect 25226 40695 25282 40704
rect 25134 40488 25190 40497
rect 25134 40423 25190 40432
rect 25136 39840 25188 39846
rect 25136 39782 25188 39788
rect 25044 37868 25096 37874
rect 25044 37810 25096 37816
rect 25044 37664 25096 37670
rect 25044 37606 25096 37612
rect 24952 36168 25004 36174
rect 24952 36110 25004 36116
rect 24964 34678 24992 36110
rect 24952 34672 25004 34678
rect 24952 34614 25004 34620
rect 24780 34190 24900 34218
rect 25056 34202 25084 37606
rect 25148 36786 25176 39782
rect 25240 38962 25268 40695
rect 25228 38956 25280 38962
rect 25228 38898 25280 38904
rect 25240 38554 25268 38898
rect 25228 38548 25280 38554
rect 25228 38490 25280 38496
rect 25228 38412 25280 38418
rect 25228 38354 25280 38360
rect 25240 38010 25268 38354
rect 25228 38004 25280 38010
rect 25228 37946 25280 37952
rect 25228 37800 25280 37806
rect 25228 37742 25280 37748
rect 25240 37505 25268 37742
rect 25226 37496 25282 37505
rect 25226 37431 25282 37440
rect 25136 36780 25188 36786
rect 25136 36722 25188 36728
rect 25148 36174 25176 36722
rect 25228 36576 25280 36582
rect 25228 36518 25280 36524
rect 25136 36168 25188 36174
rect 25136 36110 25188 36116
rect 25044 34196 25096 34202
rect 24780 33658 24808 34190
rect 25044 34138 25096 34144
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24676 33516 24728 33522
rect 24676 33458 24728 33464
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 24676 33380 24728 33386
rect 24676 33322 24728 33328
rect 24688 32026 24716 33322
rect 24676 32020 24728 32026
rect 24676 31962 24728 31968
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 24688 31142 24716 31758
rect 24780 31482 24808 33458
rect 24872 31482 24900 34002
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 25056 33522 25084 33934
rect 25136 33584 25188 33590
rect 25136 33526 25188 33532
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 24952 32836 25004 32842
rect 24952 32778 25004 32784
rect 24964 31634 24992 32778
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 25056 31736 25084 32710
rect 25148 32065 25176 33526
rect 25134 32056 25190 32065
rect 25134 31991 25190 32000
rect 25056 31708 25176 31736
rect 24964 31606 25084 31634
rect 24768 31476 24820 31482
rect 24768 31418 24820 31424
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24858 31376 24914 31385
rect 24858 31311 24914 31320
rect 24676 31136 24728 31142
rect 24676 31078 24728 31084
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24676 27396 24728 27402
rect 24676 27338 24728 27344
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24596 24857 24624 27270
rect 24582 24848 24638 24857
rect 24582 24783 24638 24792
rect 24584 24744 24636 24750
rect 24584 24686 24636 24692
rect 24596 23730 24624 24686
rect 24688 23866 24716 27338
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24584 23724 24636 23730
rect 24584 23666 24636 23672
rect 24596 23118 24624 23666
rect 24676 23520 24728 23526
rect 24676 23462 24728 23468
rect 24688 23118 24716 23462
rect 24780 23322 24808 28426
rect 24872 26874 24900 31311
rect 25056 30870 25084 31606
rect 25148 31249 25176 31708
rect 25134 31240 25190 31249
rect 25134 31175 25190 31184
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 25044 30864 25096 30870
rect 25044 30806 25096 30812
rect 25148 30802 25176 31078
rect 25136 30796 25188 30802
rect 25136 30738 25188 30744
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 25042 30696 25098 30705
rect 24964 27130 24992 30670
rect 25042 30631 25098 30640
rect 25056 28665 25084 30631
rect 25148 30122 25176 30738
rect 25136 30116 25188 30122
rect 25136 30058 25188 30064
rect 25136 29300 25188 29306
rect 25136 29242 25188 29248
rect 25148 28762 25176 29242
rect 25136 28756 25188 28762
rect 25136 28698 25188 28704
rect 25042 28656 25098 28665
rect 25042 28591 25098 28600
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 25044 28484 25096 28490
rect 25044 28426 25096 28432
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 24872 26846 24992 26874
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24872 25401 24900 26726
rect 24858 25392 24914 25401
rect 24858 25327 24914 25336
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24872 24614 24900 25230
rect 24860 24608 24912 24614
rect 24860 24550 24912 24556
rect 24872 23526 24900 24550
rect 24964 24177 24992 26846
rect 24950 24168 25006 24177
rect 24950 24103 25006 24112
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24964 23730 24992 24006
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 24768 22976 24820 22982
rect 24768 22918 24820 22924
rect 24780 21690 24808 22918
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24584 21616 24636 21622
rect 24872 21570 24900 23258
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24964 22250 24992 22986
rect 25056 22409 25084 28426
rect 25148 28082 25176 28494
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25148 27470 25176 28018
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25148 26994 25176 27406
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25134 26888 25190 26897
rect 25134 26823 25190 26832
rect 25148 23050 25176 26823
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 25042 22400 25098 22409
rect 25042 22335 25098 22344
rect 24964 22222 25084 22250
rect 24950 22128 25006 22137
rect 24950 22063 25006 22072
rect 24964 21842 24992 22063
rect 25056 22001 25084 22222
rect 25042 21992 25098 22001
rect 25042 21927 25098 21936
rect 24964 21814 25084 21842
rect 24950 21720 25006 21729
rect 24950 21655 25006 21664
rect 24584 21558 24636 21564
rect 24596 20942 24624 21558
rect 24688 21542 24900 21570
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24596 19854 24624 20878
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24596 18766 24624 19790
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24596 18086 24624 18702
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24688 15434 24716 21542
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24872 20942 24900 21422
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24872 19854 24900 20878
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24872 18766 24900 19790
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24872 18290 24900 18702
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24320 15286 24716 15314
rect 24400 14340 24452 14346
rect 24400 14282 24452 14288
rect 24412 13530 24440 14282
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24596 13326 24624 13806
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24596 12434 24624 13262
rect 24412 12406 24624 12434
rect 24412 11150 24440 12406
rect 24688 12322 24716 15286
rect 24504 12294 24716 12322
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24044 10674 24072 11086
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 24228 10742 24256 10950
rect 24216 10736 24268 10742
rect 24216 10678 24268 10684
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 24044 9722 24072 10610
rect 24412 10130 24440 10950
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24044 8498 24072 9658
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24044 7954 24072 8230
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 24504 7410 24532 12294
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 24688 11898 24716 12106
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24584 9036 24636 9042
rect 24584 8978 24636 8984
rect 24596 8498 24624 8978
rect 24780 8498 24808 18226
rect 24858 18184 24914 18193
rect 24858 18119 24914 18128
rect 24872 14618 24900 18119
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24872 12986 24900 14282
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24872 11762 24900 12786
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24596 7410 24624 8434
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24136 6390 24164 7142
rect 24504 6458 24532 7346
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24596 5234 24624 7346
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24780 5642 24808 6054
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24676 5296 24728 5302
rect 24676 5238 24728 5244
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 24584 5228 24636 5234
rect 24584 5170 24636 5176
rect 23216 4826 23244 5170
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23492 4486 23520 4558
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23400 4214 23428 4422
rect 23388 4208 23440 4214
rect 23388 4150 23440 4156
rect 23492 4026 23520 4422
rect 24044 4214 24072 4966
rect 24596 4758 24624 5170
rect 24584 4752 24636 4758
rect 24584 4694 24636 4700
rect 24596 4622 24624 4694
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 23400 4010 23520 4026
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23388 4004 23520 4010
rect 23440 3998 23520 4004
rect 23388 3946 23440 3952
rect 23952 3602 23980 4014
rect 24688 3942 24716 5238
rect 24964 5098 24992 21655
rect 25056 16522 25084 21814
rect 25148 21554 25176 22510
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25134 21448 25190 21457
rect 25134 21383 25190 21392
rect 25148 19854 25176 21383
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25148 18222 25176 19246
rect 25240 18306 25268 36518
rect 25332 25378 25360 41511
rect 25424 41274 25452 42162
rect 25516 41546 25544 44338
rect 25504 41540 25556 41546
rect 25504 41482 25556 41488
rect 25502 41440 25558 41449
rect 25502 41375 25558 41384
rect 25412 41268 25464 41274
rect 25412 41210 25464 41216
rect 25410 41168 25466 41177
rect 25410 41103 25466 41112
rect 25424 32881 25452 41103
rect 25516 38554 25544 41375
rect 25608 38593 25636 51190
rect 25700 48890 25728 52022
rect 25776 51708 26084 51728
rect 25776 51706 25782 51708
rect 25838 51706 25862 51708
rect 25918 51706 25942 51708
rect 25998 51706 26022 51708
rect 26078 51706 26084 51708
rect 25838 51654 25840 51706
rect 26020 51654 26022 51706
rect 25776 51652 25782 51654
rect 25838 51652 25862 51654
rect 25918 51652 25942 51654
rect 25998 51652 26022 51654
rect 26078 51652 26084 51654
rect 25776 51632 26084 51652
rect 25964 51536 26016 51542
rect 25964 51478 26016 51484
rect 25778 51096 25834 51105
rect 25976 51066 26004 51478
rect 26148 51468 26200 51474
rect 26148 51410 26200 51416
rect 26056 51332 26108 51338
rect 26056 51274 26108 51280
rect 25778 51031 25780 51040
rect 25832 51031 25834 51040
rect 25964 51060 26016 51066
rect 25780 51002 25832 51008
rect 25964 51002 26016 51008
rect 26068 50998 26096 51274
rect 26056 50992 26108 50998
rect 26056 50934 26108 50940
rect 25778 50824 25834 50833
rect 25778 50759 25780 50768
rect 25832 50759 25834 50768
rect 25780 50730 25832 50736
rect 25776 50620 26084 50640
rect 25776 50618 25782 50620
rect 25838 50618 25862 50620
rect 25918 50618 25942 50620
rect 25998 50618 26022 50620
rect 26078 50618 26084 50620
rect 25838 50566 25840 50618
rect 26020 50566 26022 50618
rect 25776 50564 25782 50566
rect 25838 50564 25862 50566
rect 25918 50564 25942 50566
rect 25998 50564 26022 50566
rect 26078 50564 26084 50566
rect 25776 50544 26084 50564
rect 25870 50280 25926 50289
rect 25870 50215 25926 50224
rect 25778 50008 25834 50017
rect 25778 49943 25780 49952
rect 25832 49943 25834 49952
rect 25780 49914 25832 49920
rect 25884 49774 25912 50215
rect 25872 49768 25924 49774
rect 25872 49710 25924 49716
rect 25776 49532 26084 49552
rect 25776 49530 25782 49532
rect 25838 49530 25862 49532
rect 25918 49530 25942 49532
rect 25998 49530 26022 49532
rect 26078 49530 26084 49532
rect 25838 49478 25840 49530
rect 26020 49478 26022 49530
rect 25776 49476 25782 49478
rect 25838 49476 25862 49478
rect 25918 49476 25942 49478
rect 25998 49476 26022 49478
rect 26078 49476 26084 49478
rect 25776 49456 26084 49476
rect 25780 49292 25832 49298
rect 25780 49234 25832 49240
rect 25688 48884 25740 48890
rect 25688 48826 25740 48832
rect 25792 48686 25820 49234
rect 25872 49224 25924 49230
rect 25872 49166 25924 49172
rect 25884 48890 25912 49166
rect 25872 48884 25924 48890
rect 25872 48826 25924 48832
rect 25964 48884 26016 48890
rect 25964 48826 26016 48832
rect 25780 48680 25832 48686
rect 25976 48657 26004 48826
rect 26160 48793 26188 51410
rect 26146 48784 26202 48793
rect 26252 48770 26280 54606
rect 26344 53009 26372 56902
rect 26436 55434 26464 60959
rect 26528 55622 26556 62766
rect 26620 61305 26648 67798
rect 26700 67720 26752 67726
rect 26700 67662 26752 67668
rect 26606 61296 26662 61305
rect 26606 61231 26662 61240
rect 26712 61146 26740 67662
rect 26804 64122 26832 73102
rect 26884 67720 26936 67726
rect 26884 67662 26936 67668
rect 26896 67386 26924 67662
rect 26884 67380 26936 67386
rect 26884 67322 26936 67328
rect 26884 67108 26936 67114
rect 26884 67050 26936 67056
rect 26896 66881 26924 67050
rect 26882 66872 26938 66881
rect 26988 66842 27016 74506
rect 27264 70394 27292 77454
rect 27436 74860 27488 74866
rect 27436 74802 27488 74808
rect 27344 73772 27396 73778
rect 27344 73714 27396 73720
rect 27172 70366 27292 70394
rect 27068 68264 27120 68270
rect 27068 68206 27120 68212
rect 27080 67862 27108 68206
rect 27068 67856 27120 67862
rect 27068 67798 27120 67804
rect 27068 67720 27120 67726
rect 27068 67662 27120 67668
rect 27080 67182 27108 67662
rect 27068 67176 27120 67182
rect 27068 67118 27120 67124
rect 26882 66807 26938 66816
rect 26976 66836 27028 66842
rect 26976 66778 27028 66784
rect 27172 66722 27200 70366
rect 27252 68808 27304 68814
rect 27252 68750 27304 68756
rect 27264 67289 27292 68750
rect 27250 67280 27306 67289
rect 27250 67215 27306 67224
rect 26896 66694 27200 66722
rect 27252 66700 27304 66706
rect 26792 64116 26844 64122
rect 26792 64058 26844 64064
rect 26792 63232 26844 63238
rect 26792 63174 26844 63180
rect 26804 61441 26832 63174
rect 26790 61432 26846 61441
rect 26790 61367 26846 61376
rect 26620 61118 26740 61146
rect 26620 60314 26648 61118
rect 26896 60840 26924 66694
rect 27252 66642 27304 66648
rect 26976 66632 27028 66638
rect 27028 66592 27200 66620
rect 26976 66574 27028 66580
rect 26976 66496 27028 66502
rect 26976 66438 27028 66444
rect 26988 64462 27016 66438
rect 27068 64524 27120 64530
rect 27068 64466 27120 64472
rect 26976 64456 27028 64462
rect 26976 64398 27028 64404
rect 26988 63034 27016 64398
rect 27080 63986 27108 64466
rect 27068 63980 27120 63986
rect 27068 63922 27120 63928
rect 26976 63028 27028 63034
rect 26976 62970 27028 62976
rect 27080 62778 27108 63922
rect 26988 62750 27108 62778
rect 26988 62286 27016 62750
rect 27172 62694 27200 66592
rect 27160 62688 27212 62694
rect 27160 62630 27212 62636
rect 27264 62393 27292 66642
rect 27356 65754 27384 73714
rect 27448 67930 27476 74802
rect 27528 68332 27580 68338
rect 27528 68274 27580 68280
rect 27540 68241 27568 68274
rect 27526 68232 27582 68241
rect 27526 68167 27582 68176
rect 27436 67924 27488 67930
rect 27436 67866 27488 67872
rect 27620 67856 27672 67862
rect 27526 67824 27582 67833
rect 27620 67798 27672 67804
rect 27526 67759 27582 67768
rect 27540 67232 27568 67759
rect 27632 67726 27660 67798
rect 27620 67720 27672 67726
rect 27620 67662 27672 67668
rect 27632 67590 27660 67662
rect 27620 67584 27672 67590
rect 27620 67526 27672 67532
rect 27632 67386 27660 67526
rect 27620 67380 27672 67386
rect 27620 67322 27672 67328
rect 27620 67244 27672 67250
rect 27540 67204 27620 67232
rect 27620 67186 27672 67192
rect 27436 67108 27488 67114
rect 27436 67050 27488 67056
rect 27344 65748 27396 65754
rect 27344 65690 27396 65696
rect 27448 63753 27476 67050
rect 27620 66700 27672 66706
rect 27620 66642 27672 66648
rect 27632 66298 27660 66642
rect 27620 66292 27672 66298
rect 27620 66234 27672 66240
rect 27620 65544 27672 65550
rect 27620 65486 27672 65492
rect 27632 64530 27660 65486
rect 27620 64524 27672 64530
rect 27620 64466 27672 64472
rect 27724 64122 27752 77454
rect 28552 77178 28580 78639
rect 28540 77172 28592 77178
rect 28540 77114 28592 77120
rect 28356 77036 28408 77042
rect 28356 76978 28408 76984
rect 28368 74534 28396 76978
rect 28828 76634 28856 79183
rect 29274 77752 29330 77761
rect 29274 77687 29330 77696
rect 28908 77376 28960 77382
rect 28906 77344 28908 77353
rect 28960 77344 28962 77353
rect 28906 77279 28962 77288
rect 29288 77178 29316 77687
rect 29368 77512 29420 77518
rect 29368 77454 29420 77460
rect 29380 77294 29408 77454
rect 30104 77376 30156 77382
rect 30104 77318 30156 77324
rect 29380 77266 29500 77294
rect 29276 77172 29328 77178
rect 29276 77114 29328 77120
rect 29092 77036 29144 77042
rect 29092 76978 29144 76984
rect 29000 76968 29052 76974
rect 29000 76910 29052 76916
rect 28816 76628 28868 76634
rect 28816 76570 28868 76576
rect 28368 74506 28580 74534
rect 28448 69420 28500 69426
rect 28448 69362 28500 69368
rect 27804 67720 27856 67726
rect 27802 67688 27804 67697
rect 27856 67688 27858 67697
rect 27802 67623 27858 67632
rect 27804 67584 27856 67590
rect 27802 67552 27804 67561
rect 27856 67552 27858 67561
rect 27802 67487 27858 67496
rect 27804 67380 27856 67386
rect 27804 67322 27856 67328
rect 27816 66706 27844 67322
rect 27896 67312 27948 67318
rect 27896 67254 27948 67260
rect 27804 66700 27856 66706
rect 27804 66642 27856 66648
rect 27804 66564 27856 66570
rect 27804 66506 27856 66512
rect 27816 65754 27844 66506
rect 27804 65748 27856 65754
rect 27804 65690 27856 65696
rect 27816 64462 27844 65690
rect 27908 65657 27936 67254
rect 28264 67244 28316 67250
rect 28264 67186 28316 67192
rect 27988 66156 28040 66162
rect 27988 66098 28040 66104
rect 27894 65648 27950 65657
rect 27894 65583 27950 65592
rect 27896 65544 27948 65550
rect 27896 65486 27948 65492
rect 27908 65210 27936 65486
rect 27896 65204 27948 65210
rect 27896 65146 27948 65152
rect 27804 64456 27856 64462
rect 27896 64456 27948 64462
rect 27804 64398 27856 64404
rect 27894 64424 27896 64433
rect 27948 64424 27950 64433
rect 27712 64116 27764 64122
rect 27712 64058 27764 64064
rect 27528 64048 27580 64054
rect 27528 63990 27580 63996
rect 27434 63744 27490 63753
rect 27434 63679 27490 63688
rect 27540 62937 27568 63990
rect 27712 63844 27764 63850
rect 27712 63786 27764 63792
rect 27724 63578 27752 63786
rect 27712 63572 27764 63578
rect 27712 63514 27764 63520
rect 27712 63368 27764 63374
rect 27712 63310 27764 63316
rect 27620 63300 27672 63306
rect 27620 63242 27672 63248
rect 27632 63209 27660 63242
rect 27618 63200 27674 63209
rect 27618 63135 27674 63144
rect 27526 62928 27582 62937
rect 27526 62863 27582 62872
rect 27620 62892 27672 62898
rect 27620 62834 27672 62840
rect 27344 62688 27396 62694
rect 27344 62630 27396 62636
rect 27250 62384 27306 62393
rect 27250 62319 27306 62328
rect 26976 62280 27028 62286
rect 27252 62280 27304 62286
rect 26976 62222 27028 62228
rect 27172 62240 27252 62268
rect 26988 61810 27016 62222
rect 26976 61804 27028 61810
rect 26976 61746 27028 61752
rect 26988 61198 27016 61746
rect 26976 61192 27028 61198
rect 26976 61134 27028 61140
rect 27172 61033 27200 62240
rect 27252 62222 27304 62228
rect 27356 62132 27384 62630
rect 27436 62280 27488 62286
rect 27632 62257 27660 62834
rect 27724 62801 27752 63310
rect 27710 62792 27766 62801
rect 27710 62727 27766 62736
rect 27712 62348 27764 62354
rect 27712 62290 27764 62296
rect 27436 62222 27488 62228
rect 27618 62248 27674 62257
rect 27264 62104 27384 62132
rect 27448 62121 27476 62222
rect 27618 62183 27674 62192
rect 27434 62112 27490 62121
rect 26974 61024 27030 61033
rect 26974 60959 27030 60968
rect 27158 61024 27214 61033
rect 27158 60959 27214 60968
rect 26712 60812 26924 60840
rect 26712 60314 26740 60812
rect 26988 60734 27016 60959
rect 26896 60706 27016 60734
rect 27068 60716 27120 60722
rect 26792 60648 26844 60654
rect 26792 60590 26844 60596
rect 26608 60308 26660 60314
rect 26608 60250 26660 60256
rect 26700 60308 26752 60314
rect 26700 60250 26752 60256
rect 26804 60194 26832 60590
rect 26712 60166 26832 60194
rect 26608 60104 26660 60110
rect 26606 60072 26608 60081
rect 26660 60072 26662 60081
rect 26606 60007 26662 60016
rect 26608 59968 26660 59974
rect 26608 59910 26660 59916
rect 26620 57633 26648 59910
rect 26712 57798 26740 60166
rect 26790 60072 26846 60081
rect 26790 60007 26846 60016
rect 26804 59974 26832 60007
rect 26792 59968 26844 59974
rect 26792 59910 26844 59916
rect 26896 59770 26924 60706
rect 27068 60658 27120 60664
rect 26974 60616 27030 60625
rect 27080 60586 27108 60658
rect 26974 60551 27030 60560
rect 27068 60580 27120 60586
rect 26884 59764 26936 59770
rect 26884 59706 26936 59712
rect 26988 59650 27016 60551
rect 27068 60522 27120 60528
rect 27066 60344 27122 60353
rect 27066 60279 27122 60288
rect 26804 59622 27016 59650
rect 26700 57792 26752 57798
rect 26700 57734 26752 57740
rect 26606 57624 26662 57633
rect 26606 57559 26662 57568
rect 26608 57520 26660 57526
rect 26608 57462 26660 57468
rect 26620 56166 26648 57462
rect 26608 56160 26660 56166
rect 26608 56102 26660 56108
rect 26516 55616 26568 55622
rect 26516 55558 26568 55564
rect 26436 55406 26648 55434
rect 26424 55344 26476 55350
rect 26424 55286 26476 55292
rect 26330 53000 26386 53009
rect 26330 52935 26386 52944
rect 26332 52896 26384 52902
rect 26332 52838 26384 52844
rect 26344 51270 26372 52838
rect 26332 51264 26384 51270
rect 26436 51241 26464 55286
rect 26516 53440 26568 53446
rect 26516 53382 26568 53388
rect 26528 53174 26556 53382
rect 26516 53168 26568 53174
rect 26516 53110 26568 53116
rect 26620 52698 26648 55406
rect 26608 52692 26660 52698
rect 26608 52634 26660 52640
rect 26712 52442 26740 57734
rect 26804 56001 26832 59622
rect 26884 59560 26936 59566
rect 26884 59502 26936 59508
rect 26974 59528 27030 59537
rect 26790 55992 26846 56001
rect 26790 55927 26846 55936
rect 26792 55616 26844 55622
rect 26792 55558 26844 55564
rect 26528 52414 26740 52442
rect 26332 51206 26384 51212
rect 26422 51232 26478 51241
rect 26422 51167 26478 51176
rect 26424 51060 26476 51066
rect 26424 51002 26476 51008
rect 26332 49836 26384 49842
rect 26332 49778 26384 49784
rect 26344 49076 26372 49778
rect 26436 49230 26464 51002
rect 26528 49230 26556 52414
rect 26700 52352 26752 52358
rect 26700 52294 26752 52300
rect 26608 52080 26660 52086
rect 26606 52048 26608 52057
rect 26660 52048 26662 52057
rect 26606 51983 26662 51992
rect 26608 51944 26660 51950
rect 26608 51886 26660 51892
rect 26424 49224 26476 49230
rect 26424 49166 26476 49172
rect 26516 49224 26568 49230
rect 26516 49166 26568 49172
rect 26424 49088 26476 49094
rect 26344 49048 26424 49076
rect 26424 49030 26476 49036
rect 26330 48784 26386 48793
rect 26252 48742 26330 48770
rect 26146 48719 26202 48728
rect 26436 48754 26464 49030
rect 26330 48719 26386 48728
rect 26424 48748 26476 48754
rect 26424 48690 26476 48696
rect 26148 48680 26200 48686
rect 25780 48622 25832 48628
rect 25962 48648 26018 48657
rect 25792 48532 25820 48622
rect 26528 48634 26556 49166
rect 26148 48622 26200 48628
rect 25962 48583 26018 48592
rect 25700 48504 25820 48532
rect 25700 48142 25728 48504
rect 25776 48444 26084 48464
rect 25776 48442 25782 48444
rect 25838 48442 25862 48444
rect 25918 48442 25942 48444
rect 25998 48442 26022 48444
rect 26078 48442 26084 48444
rect 25838 48390 25840 48442
rect 26020 48390 26022 48442
rect 25776 48388 25782 48390
rect 25838 48388 25862 48390
rect 25918 48388 25942 48390
rect 25998 48388 26022 48390
rect 26078 48388 26084 48390
rect 25776 48368 26084 48388
rect 26160 48362 26188 48622
rect 26344 48606 26556 48634
rect 26160 48346 26280 48362
rect 26160 48340 26292 48346
rect 26160 48334 26240 48340
rect 26344 48328 26372 48606
rect 26516 48544 26568 48550
rect 26516 48486 26568 48492
rect 26528 48346 26556 48486
rect 26424 48340 26476 48346
rect 26344 48300 26424 48328
rect 26240 48282 26292 48288
rect 26424 48282 26476 48288
rect 26516 48340 26568 48346
rect 26516 48282 26568 48288
rect 26148 48272 26200 48278
rect 26148 48214 26200 48220
rect 26330 48240 26386 48249
rect 25688 48136 25740 48142
rect 25688 48078 25740 48084
rect 26056 48136 26108 48142
rect 26056 48078 26108 48084
rect 25700 46034 25728 48078
rect 25962 47832 26018 47841
rect 25962 47767 25964 47776
rect 26016 47767 26018 47776
rect 25964 47738 26016 47744
rect 26068 47734 26096 48078
rect 26056 47728 26108 47734
rect 26056 47670 26108 47676
rect 26160 47666 26188 48214
rect 26330 48175 26386 48184
rect 26238 48104 26294 48113
rect 26238 48039 26294 48048
rect 26148 47660 26200 47666
rect 26148 47602 26200 47608
rect 25776 47356 26084 47376
rect 25776 47354 25782 47356
rect 25838 47354 25862 47356
rect 25918 47354 25942 47356
rect 25998 47354 26022 47356
rect 26078 47354 26084 47356
rect 25838 47302 25840 47354
rect 26020 47302 26022 47354
rect 25776 47300 25782 47302
rect 25838 47300 25862 47302
rect 25918 47300 25942 47302
rect 25998 47300 26022 47302
rect 26078 47300 26084 47302
rect 25776 47280 26084 47300
rect 26056 47184 26108 47190
rect 26056 47126 26108 47132
rect 26068 46510 26096 47126
rect 26160 47122 26188 47602
rect 26148 47116 26200 47122
rect 26148 47058 26200 47064
rect 26148 46980 26200 46986
rect 26148 46922 26200 46928
rect 25780 46504 25832 46510
rect 25778 46472 25780 46481
rect 26056 46504 26108 46510
rect 25832 46472 25834 46481
rect 26056 46446 26108 46452
rect 25778 46407 25834 46416
rect 25776 46268 26084 46288
rect 25776 46266 25782 46268
rect 25838 46266 25862 46268
rect 25918 46266 25942 46268
rect 25998 46266 26022 46268
rect 26078 46266 26084 46268
rect 25838 46214 25840 46266
rect 26020 46214 26022 46266
rect 25776 46212 25782 46214
rect 25838 46212 25862 46214
rect 25918 46212 25942 46214
rect 25998 46212 26022 46214
rect 26078 46212 26084 46214
rect 25776 46192 26084 46212
rect 25688 46028 25740 46034
rect 25688 45970 25740 45976
rect 25688 45824 25740 45830
rect 25688 45766 25740 45772
rect 25700 42888 25728 45766
rect 25776 45180 26084 45200
rect 25776 45178 25782 45180
rect 25838 45178 25862 45180
rect 25918 45178 25942 45180
rect 25998 45178 26022 45180
rect 26078 45178 26084 45180
rect 25838 45126 25840 45178
rect 26020 45126 26022 45178
rect 25776 45124 25782 45126
rect 25838 45124 25862 45126
rect 25918 45124 25942 45126
rect 25998 45124 26022 45126
rect 26078 45124 26084 45126
rect 25776 45104 26084 45124
rect 25776 44092 26084 44112
rect 25776 44090 25782 44092
rect 25838 44090 25862 44092
rect 25918 44090 25942 44092
rect 25998 44090 26022 44092
rect 26078 44090 26084 44092
rect 25838 44038 25840 44090
rect 26020 44038 26022 44090
rect 25776 44036 25782 44038
rect 25838 44036 25862 44038
rect 25918 44036 25942 44038
rect 25998 44036 26022 44038
rect 26078 44036 26084 44038
rect 25776 44016 26084 44036
rect 25776 43004 26084 43024
rect 25776 43002 25782 43004
rect 25838 43002 25862 43004
rect 25918 43002 25942 43004
rect 25998 43002 26022 43004
rect 26078 43002 26084 43004
rect 25838 42950 25840 43002
rect 26020 42950 26022 43002
rect 25776 42948 25782 42950
rect 25838 42948 25862 42950
rect 25918 42948 25942 42950
rect 25998 42948 26022 42950
rect 26078 42948 26084 42950
rect 25776 42928 26084 42948
rect 25700 42860 26004 42888
rect 25870 42800 25926 42809
rect 25780 42764 25832 42770
rect 25870 42735 25926 42744
rect 25780 42706 25832 42712
rect 25688 42628 25740 42634
rect 25688 42570 25740 42576
rect 25700 41682 25728 42570
rect 25792 42537 25820 42706
rect 25884 42634 25912 42735
rect 25872 42628 25924 42634
rect 25872 42570 25924 42576
rect 25778 42528 25834 42537
rect 25778 42463 25834 42472
rect 25780 42356 25832 42362
rect 25780 42298 25832 42304
rect 25792 42158 25820 42298
rect 25884 42265 25912 42570
rect 25976 42566 26004 42860
rect 25964 42560 26016 42566
rect 25964 42502 26016 42508
rect 26056 42560 26108 42566
rect 26056 42502 26108 42508
rect 25870 42256 25926 42265
rect 25870 42191 25926 42200
rect 25780 42152 25832 42158
rect 25780 42094 25832 42100
rect 25976 42090 26004 42502
rect 26068 42090 26096 42502
rect 25964 42084 26016 42090
rect 25964 42026 26016 42032
rect 26056 42084 26108 42090
rect 26056 42026 26108 42032
rect 25776 41916 26084 41936
rect 25776 41914 25782 41916
rect 25838 41914 25862 41916
rect 25918 41914 25942 41916
rect 25998 41914 26022 41916
rect 26078 41914 26084 41916
rect 25838 41862 25840 41914
rect 26020 41862 26022 41914
rect 25776 41860 25782 41862
rect 25838 41860 25862 41862
rect 25918 41860 25942 41862
rect 25998 41860 26022 41862
rect 26078 41860 26084 41862
rect 25776 41840 26084 41860
rect 25964 41744 26016 41750
rect 25964 41686 26016 41692
rect 25688 41676 25740 41682
rect 25688 41618 25740 41624
rect 25686 41576 25742 41585
rect 25686 41511 25742 41520
rect 25594 38584 25650 38593
rect 25504 38548 25556 38554
rect 25594 38519 25650 38528
rect 25504 38490 25556 38496
rect 25700 38400 25728 41511
rect 25780 41472 25832 41478
rect 25780 41414 25832 41420
rect 25792 41274 25820 41414
rect 25780 41268 25832 41274
rect 25780 41210 25832 41216
rect 25792 40916 25820 41210
rect 25976 41041 26004 41686
rect 26056 41540 26108 41546
rect 26056 41482 26108 41488
rect 25962 41032 26018 41041
rect 25962 40967 26018 40976
rect 26068 40984 26096 41482
rect 26160 41449 26188 46922
rect 26252 42702 26280 48039
rect 26344 45121 26372 48175
rect 26424 47456 26476 47462
rect 26424 47398 26476 47404
rect 26436 45558 26464 47398
rect 26620 47258 26648 51886
rect 26712 49434 26740 52294
rect 26700 49428 26752 49434
rect 26700 49370 26752 49376
rect 26700 49292 26752 49298
rect 26700 49234 26752 49240
rect 26712 48686 26740 49234
rect 26804 49201 26832 55558
rect 26896 52358 26924 59502
rect 26974 59463 26976 59472
rect 27028 59463 27030 59472
rect 26976 59434 27028 59440
rect 26976 58540 27028 58546
rect 26976 58482 27028 58488
rect 26988 58342 27016 58482
rect 26976 58336 27028 58342
rect 26976 58278 27028 58284
rect 26976 57860 27028 57866
rect 26976 57802 27028 57808
rect 26988 57458 27016 57802
rect 26976 57452 27028 57458
rect 26976 57394 27028 57400
rect 26988 54874 27016 57394
rect 26976 54868 27028 54874
rect 26976 54810 27028 54816
rect 26974 54768 27030 54777
rect 26974 54703 26976 54712
rect 27028 54703 27030 54712
rect 26976 54674 27028 54680
rect 26976 53576 27028 53582
rect 26976 53518 27028 53524
rect 26988 53038 27016 53518
rect 26976 53032 27028 53038
rect 26976 52974 27028 52980
rect 26988 52494 27016 52974
rect 26976 52488 27028 52494
rect 26976 52430 27028 52436
rect 26884 52352 26936 52358
rect 26884 52294 26936 52300
rect 26988 52000 27016 52430
rect 26896 51972 27016 52000
rect 26896 49609 26924 51972
rect 26976 51876 27028 51882
rect 26976 51818 27028 51824
rect 26882 49600 26938 49609
rect 26882 49535 26938 49544
rect 26988 49473 27016 51818
rect 26974 49464 27030 49473
rect 26974 49399 27030 49408
rect 27080 49201 27108 60279
rect 27160 60240 27212 60246
rect 27158 60208 27160 60217
rect 27212 60208 27214 60217
rect 27158 60143 27214 60152
rect 27160 60104 27212 60110
rect 27160 60046 27212 60052
rect 27172 59634 27200 60046
rect 27160 59628 27212 59634
rect 27160 59570 27212 59576
rect 27158 58848 27214 58857
rect 27158 58783 27214 58792
rect 27172 58070 27200 58783
rect 27160 58064 27212 58070
rect 27160 58006 27212 58012
rect 27160 57928 27212 57934
rect 27160 57870 27212 57876
rect 27172 56302 27200 57870
rect 27160 56296 27212 56302
rect 27160 56238 27212 56244
rect 27172 55690 27200 56238
rect 27160 55684 27212 55690
rect 27160 55626 27212 55632
rect 27172 53990 27200 55626
rect 27160 53984 27212 53990
rect 27160 53926 27212 53932
rect 27172 49722 27200 53926
rect 27264 51762 27292 62104
rect 27434 62047 27490 62056
rect 27528 61804 27580 61810
rect 27344 61788 27396 61794
rect 27528 61746 27580 61752
rect 27344 61730 27396 61736
rect 27356 61033 27384 61730
rect 27436 61600 27488 61606
rect 27436 61542 27488 61548
rect 27448 61402 27476 61542
rect 27436 61396 27488 61402
rect 27436 61338 27488 61344
rect 27342 61024 27398 61033
rect 27342 60959 27398 60968
rect 27540 60858 27568 61746
rect 27724 61248 27752 62290
rect 27632 61220 27752 61248
rect 27528 60852 27580 60858
rect 27528 60794 27580 60800
rect 27436 60716 27488 60722
rect 27436 60658 27488 60664
rect 27344 60512 27396 60518
rect 27344 60454 27396 60460
rect 27356 59634 27384 60454
rect 27344 59628 27396 59634
rect 27344 59570 27396 59576
rect 27344 59424 27396 59430
rect 27344 59366 27396 59372
rect 27356 58546 27384 59366
rect 27448 59090 27476 60658
rect 27632 60466 27660 61220
rect 27710 61160 27766 61169
rect 27710 61095 27766 61104
rect 27540 60438 27660 60466
rect 27436 59084 27488 59090
rect 27436 59026 27488 59032
rect 27436 58948 27488 58954
rect 27436 58890 27488 58896
rect 27344 58540 27396 58546
rect 27344 58482 27396 58488
rect 27448 58426 27476 58890
rect 27356 58398 27476 58426
rect 27356 57866 27384 58398
rect 27344 57860 27396 57866
rect 27344 57802 27396 57808
rect 27356 57390 27384 57802
rect 27436 57792 27488 57798
rect 27434 57760 27436 57769
rect 27488 57760 27490 57769
rect 27434 57695 27490 57704
rect 27434 57488 27490 57497
rect 27434 57423 27490 57432
rect 27344 57384 27396 57390
rect 27344 57326 27396 57332
rect 27356 57225 27384 57326
rect 27342 57216 27398 57225
rect 27342 57151 27398 57160
rect 27342 57080 27398 57089
rect 27342 57015 27398 57024
rect 27356 56982 27384 57015
rect 27344 56976 27396 56982
rect 27344 56918 27396 56924
rect 27448 56914 27476 57423
rect 27436 56908 27488 56914
rect 27436 56850 27488 56856
rect 27344 56840 27396 56846
rect 27344 56782 27396 56788
rect 27356 56234 27384 56782
rect 27344 56228 27396 56234
rect 27344 56170 27396 56176
rect 27448 55826 27476 56850
rect 27436 55820 27488 55826
rect 27356 55780 27436 55808
rect 27356 55146 27384 55780
rect 27436 55762 27488 55768
rect 27434 55584 27490 55593
rect 27434 55519 27490 55528
rect 27344 55140 27396 55146
rect 27344 55082 27396 55088
rect 27356 54602 27384 55082
rect 27448 54806 27476 55519
rect 27540 55418 27568 60438
rect 27724 60194 27752 61095
rect 27816 60858 27844 64398
rect 27894 64359 27950 64368
rect 27896 62144 27948 62150
rect 27894 62112 27896 62121
rect 27948 62112 27950 62121
rect 27894 62047 27950 62056
rect 27896 61668 27948 61674
rect 27896 61610 27948 61616
rect 27908 61198 27936 61610
rect 27896 61192 27948 61198
rect 27896 61134 27948 61140
rect 27894 61024 27950 61033
rect 27894 60959 27950 60968
rect 27804 60852 27856 60858
rect 27804 60794 27856 60800
rect 27632 60166 27752 60194
rect 27632 58682 27660 60166
rect 27804 60104 27856 60110
rect 27804 60046 27856 60052
rect 27712 59628 27764 59634
rect 27712 59570 27764 59576
rect 27724 58682 27752 59570
rect 27620 58676 27672 58682
rect 27620 58618 27672 58624
rect 27712 58676 27764 58682
rect 27712 58618 27764 58624
rect 27618 58576 27674 58585
rect 27618 58511 27674 58520
rect 27528 55412 27580 55418
rect 27528 55354 27580 55360
rect 27436 54800 27488 54806
rect 27632 54754 27660 58511
rect 27436 54742 27488 54748
rect 27448 54641 27476 54742
rect 27540 54726 27660 54754
rect 27434 54632 27490 54641
rect 27344 54596 27396 54602
rect 27434 54567 27490 54576
rect 27344 54538 27396 54544
rect 27356 54330 27384 54538
rect 27434 54496 27490 54505
rect 27434 54431 27490 54440
rect 27344 54324 27396 54330
rect 27344 54266 27396 54272
rect 27448 54194 27476 54431
rect 27436 54188 27488 54194
rect 27436 54130 27488 54136
rect 27344 53100 27396 53106
rect 27344 53042 27396 53048
rect 27356 52494 27384 53042
rect 27540 52986 27568 54726
rect 27620 54596 27672 54602
rect 27620 54538 27672 54544
rect 27632 54126 27660 54538
rect 27620 54120 27672 54126
rect 27620 54062 27672 54068
rect 27724 53530 27752 58618
rect 27632 53502 27752 53530
rect 27632 53106 27660 53502
rect 27712 53440 27764 53446
rect 27712 53382 27764 53388
rect 27724 53281 27752 53382
rect 27710 53272 27766 53281
rect 27710 53207 27766 53216
rect 27620 53100 27672 53106
rect 27620 53042 27672 53048
rect 27540 52958 27660 52986
rect 27528 52624 27580 52630
rect 27632 52601 27660 52958
rect 27712 52964 27764 52970
rect 27712 52906 27764 52912
rect 27528 52566 27580 52572
rect 27618 52592 27674 52601
rect 27344 52488 27396 52494
rect 27344 52430 27396 52436
rect 27356 52018 27384 52430
rect 27436 52352 27488 52358
rect 27436 52294 27488 52300
rect 27448 52154 27476 52294
rect 27436 52148 27488 52154
rect 27436 52090 27488 52096
rect 27344 52012 27396 52018
rect 27344 51954 27396 51960
rect 27264 51734 27384 51762
rect 27252 50176 27304 50182
rect 27252 50118 27304 50124
rect 27264 49842 27292 50118
rect 27252 49836 27304 49842
rect 27252 49778 27304 49784
rect 27172 49694 27292 49722
rect 27160 49360 27212 49366
rect 27160 49302 27212 49308
rect 26790 49192 26846 49201
rect 26790 49127 26846 49136
rect 27066 49192 27122 49201
rect 27066 49127 27122 49136
rect 26976 49088 27028 49094
rect 26976 49030 27028 49036
rect 26988 48890 27016 49030
rect 26976 48884 27028 48890
rect 26976 48826 27028 48832
rect 27172 48754 27200 49302
rect 27264 48906 27292 49694
rect 27356 49065 27384 51734
rect 27434 49736 27490 49745
rect 27434 49671 27436 49680
rect 27488 49671 27490 49680
rect 27436 49642 27488 49648
rect 27434 49464 27490 49473
rect 27434 49399 27490 49408
rect 27448 49366 27476 49399
rect 27436 49360 27488 49366
rect 27436 49302 27488 49308
rect 27436 49224 27488 49230
rect 27436 49166 27488 49172
rect 27342 49056 27398 49065
rect 27342 48991 27398 49000
rect 27264 48878 27384 48906
rect 26884 48748 26936 48754
rect 26884 48690 26936 48696
rect 27160 48748 27212 48754
rect 27160 48690 27212 48696
rect 26700 48680 26752 48686
rect 26700 48622 26752 48628
rect 26712 48142 26740 48622
rect 26896 48550 26924 48690
rect 27066 48648 27122 48657
rect 26988 48606 27066 48634
rect 26884 48544 26936 48550
rect 26790 48512 26846 48521
rect 26884 48486 26936 48492
rect 26790 48447 26846 48456
rect 26700 48136 26752 48142
rect 26700 48078 26752 48084
rect 26608 47252 26660 47258
rect 26608 47194 26660 47200
rect 26608 47116 26660 47122
rect 26608 47058 26660 47064
rect 26528 46918 26556 46949
rect 26516 46912 26568 46918
rect 26514 46880 26516 46889
rect 26568 46880 26570 46889
rect 26514 46815 26570 46824
rect 26528 46714 26556 46815
rect 26516 46708 26568 46714
rect 26516 46650 26568 46656
rect 26516 46504 26568 46510
rect 26516 46446 26568 46452
rect 26424 45552 26476 45558
rect 26424 45494 26476 45500
rect 26330 45112 26386 45121
rect 26330 45047 26386 45056
rect 26332 45008 26384 45014
rect 26332 44950 26384 44956
rect 26344 43994 26372 44950
rect 26332 43988 26384 43994
rect 26332 43930 26384 43936
rect 26424 43648 26476 43654
rect 26424 43590 26476 43596
rect 26436 43110 26464 43590
rect 26424 43104 26476 43110
rect 26424 43046 26476 43052
rect 26240 42696 26292 42702
rect 26240 42638 26292 42644
rect 26240 42288 26292 42294
rect 26240 42230 26292 42236
rect 26424 42288 26476 42294
rect 26424 42230 26476 42236
rect 26146 41440 26202 41449
rect 26146 41375 26202 41384
rect 26252 41274 26280 42230
rect 26332 42084 26384 42090
rect 26332 42026 26384 42032
rect 26240 41268 26292 41274
rect 26240 41210 26292 41216
rect 26068 40956 26280 40984
rect 25792 40888 26188 40916
rect 25776 40828 26084 40848
rect 25776 40826 25782 40828
rect 25838 40826 25862 40828
rect 25918 40826 25942 40828
rect 25998 40826 26022 40828
rect 26078 40826 26084 40828
rect 25838 40774 25840 40826
rect 26020 40774 26022 40826
rect 25776 40772 25782 40774
rect 25838 40772 25862 40774
rect 25918 40772 25942 40774
rect 25998 40772 26022 40774
rect 26078 40772 26084 40774
rect 25776 40752 26084 40772
rect 25780 40588 25832 40594
rect 25780 40530 25832 40536
rect 25792 40361 25820 40530
rect 25870 40488 25926 40497
rect 25870 40423 25872 40432
rect 25924 40423 25926 40432
rect 26054 40488 26110 40497
rect 26054 40423 26056 40432
rect 25872 40394 25924 40400
rect 26108 40423 26110 40432
rect 26056 40394 26108 40400
rect 25778 40352 25834 40361
rect 25778 40287 25834 40296
rect 26056 40180 26108 40186
rect 26056 40122 26108 40128
rect 26068 39828 26096 40122
rect 26160 39896 26188 40888
rect 26252 40186 26280 40956
rect 26344 40497 26372 42026
rect 26436 41750 26464 42230
rect 26528 42226 26556 46446
rect 26516 42220 26568 42226
rect 26516 42162 26568 42168
rect 26424 41744 26476 41750
rect 26424 41686 26476 41692
rect 26528 41596 26556 42162
rect 26436 41568 26556 41596
rect 26436 41070 26464 41568
rect 26516 41472 26568 41478
rect 26514 41440 26516 41449
rect 26568 41440 26570 41449
rect 26514 41375 26570 41384
rect 26514 41304 26570 41313
rect 26514 41239 26570 41248
rect 26424 41064 26476 41070
rect 26424 41006 26476 41012
rect 26330 40488 26386 40497
rect 26330 40423 26386 40432
rect 26332 40384 26384 40390
rect 26332 40326 26384 40332
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 26160 39868 26280 39896
rect 26068 39800 26188 39828
rect 25776 39740 26084 39760
rect 25776 39738 25782 39740
rect 25838 39738 25862 39740
rect 25918 39738 25942 39740
rect 25998 39738 26022 39740
rect 26078 39738 26084 39740
rect 25838 39686 25840 39738
rect 26020 39686 26022 39738
rect 25776 39684 25782 39686
rect 25838 39684 25862 39686
rect 25918 39684 25942 39686
rect 25998 39684 26022 39686
rect 26078 39684 26084 39686
rect 25776 39664 26084 39684
rect 26160 39624 26188 39800
rect 26068 39596 26188 39624
rect 25962 39400 26018 39409
rect 25872 39364 25924 39370
rect 25962 39335 26018 39344
rect 25872 39306 25924 39312
rect 25884 39001 25912 39306
rect 25976 39098 26004 39335
rect 26068 39098 26096 39596
rect 26146 39536 26202 39545
rect 26146 39471 26202 39480
rect 25964 39092 26016 39098
rect 25964 39034 26016 39040
rect 26056 39092 26108 39098
rect 26056 39034 26108 39040
rect 25870 38992 25926 39001
rect 25870 38927 25926 38936
rect 25872 38888 25924 38894
rect 25870 38856 25872 38865
rect 25924 38856 25926 38865
rect 26068 38826 26096 39034
rect 25870 38791 25926 38800
rect 26056 38820 26108 38826
rect 26056 38762 26108 38768
rect 25776 38652 26084 38672
rect 25776 38650 25782 38652
rect 25838 38650 25862 38652
rect 25918 38650 25942 38652
rect 25998 38650 26022 38652
rect 26078 38650 26084 38652
rect 25838 38598 25840 38650
rect 26020 38598 26022 38650
rect 25776 38596 25782 38598
rect 25838 38596 25862 38598
rect 25918 38596 25942 38598
rect 25998 38596 26022 38598
rect 26078 38596 26084 38598
rect 25776 38576 26084 38596
rect 25608 38372 25728 38400
rect 25778 38448 25834 38457
rect 26054 38448 26110 38457
rect 25778 38383 25834 38392
rect 25872 38412 25924 38418
rect 25608 38298 25636 38372
rect 25792 38350 25820 38383
rect 26054 38383 26110 38392
rect 25872 38354 25924 38360
rect 25780 38344 25832 38350
rect 25504 38276 25556 38282
rect 25608 38270 25728 38298
rect 25780 38286 25832 38292
rect 25504 38218 25556 38224
rect 25516 37330 25544 38218
rect 25594 38176 25650 38185
rect 25594 38111 25650 38120
rect 25504 37324 25556 37330
rect 25504 37266 25556 37272
rect 25502 37224 25558 37233
rect 25502 37159 25558 37168
rect 25410 32872 25466 32881
rect 25410 32807 25466 32816
rect 25412 31884 25464 31890
rect 25412 31826 25464 31832
rect 25424 30734 25452 31826
rect 25516 31346 25544 37159
rect 25608 36582 25636 38111
rect 25700 36689 25728 38270
rect 25884 37942 25912 38354
rect 26068 38282 26096 38383
rect 26056 38276 26108 38282
rect 26056 38218 26108 38224
rect 26068 38010 26096 38218
rect 26056 38004 26108 38010
rect 26056 37946 26108 37952
rect 25872 37936 25924 37942
rect 25872 37878 25924 37884
rect 25776 37564 26084 37584
rect 25776 37562 25782 37564
rect 25838 37562 25862 37564
rect 25918 37562 25942 37564
rect 25998 37562 26022 37564
rect 26078 37562 26084 37564
rect 25838 37510 25840 37562
rect 26020 37510 26022 37562
rect 25776 37508 25782 37510
rect 25838 37508 25862 37510
rect 25918 37508 25942 37510
rect 25998 37508 26022 37510
rect 26078 37508 26084 37510
rect 25776 37488 26084 37508
rect 26056 37120 26108 37126
rect 26054 37088 26056 37097
rect 26108 37088 26110 37097
rect 26054 37023 26110 37032
rect 26160 36802 26188 39471
rect 26252 39438 26280 39868
rect 26240 39432 26292 39438
rect 26240 39374 26292 39380
rect 26252 38282 26280 39374
rect 26344 39137 26372 40326
rect 26436 39273 26464 41006
rect 26422 39264 26478 39273
rect 26422 39199 26478 39208
rect 26330 39128 26386 39137
rect 26330 39063 26386 39072
rect 26528 39001 26556 41239
rect 26620 39642 26648 47058
rect 26712 42090 26740 48078
rect 26700 42084 26752 42090
rect 26700 42026 26752 42032
rect 26698 41984 26754 41993
rect 26698 41919 26754 41928
rect 26608 39636 26660 39642
rect 26608 39578 26660 39584
rect 26514 38992 26570 39001
rect 26514 38927 26570 38936
rect 26514 38856 26570 38865
rect 26514 38791 26570 38800
rect 26330 38720 26386 38729
rect 26330 38655 26386 38664
rect 26240 38276 26292 38282
rect 26240 38218 26292 38224
rect 26240 37800 26292 37806
rect 26240 37742 26292 37748
rect 26068 36774 26188 36802
rect 25780 36712 25832 36718
rect 25686 36680 25742 36689
rect 25780 36654 25832 36660
rect 25686 36615 25742 36624
rect 25596 36576 25648 36582
rect 25792 36564 25820 36654
rect 26068 36650 26096 36774
rect 26148 36712 26200 36718
rect 26148 36654 26200 36660
rect 26056 36644 26108 36650
rect 26056 36586 26108 36592
rect 25596 36518 25648 36524
rect 25700 36536 25820 36564
rect 25700 36360 25728 36536
rect 25776 36476 26084 36496
rect 25776 36474 25782 36476
rect 25838 36474 25862 36476
rect 25918 36474 25942 36476
rect 25998 36474 26022 36476
rect 26078 36474 26084 36476
rect 25838 36422 25840 36474
rect 26020 36422 26022 36474
rect 25776 36420 25782 36422
rect 25838 36420 25862 36422
rect 25918 36420 25942 36422
rect 25998 36420 26022 36422
rect 26078 36420 26084 36422
rect 25776 36400 26084 36420
rect 25700 36332 25912 36360
rect 25780 36168 25832 36174
rect 25594 36136 25650 36145
rect 25780 36110 25832 36116
rect 25594 36071 25650 36080
rect 25608 34134 25636 36071
rect 25792 35737 25820 36110
rect 25884 36106 25912 36332
rect 25964 36304 26016 36310
rect 25964 36246 26016 36252
rect 25872 36100 25924 36106
rect 25872 36042 25924 36048
rect 25884 35873 25912 36042
rect 25870 35864 25926 35873
rect 25976 35834 26004 36246
rect 26056 36032 26108 36038
rect 26054 36000 26056 36009
rect 26160 36020 26188 36654
rect 26252 36106 26280 37742
rect 26240 36100 26292 36106
rect 26240 36042 26292 36048
rect 26108 36000 26188 36020
rect 26110 35992 26188 36000
rect 26054 35935 26110 35944
rect 25870 35799 25926 35808
rect 25964 35828 26016 35834
rect 25964 35770 26016 35776
rect 25778 35728 25834 35737
rect 25778 35663 25834 35672
rect 26344 35494 26372 38655
rect 26422 38584 26478 38593
rect 26422 38519 26478 38528
rect 26436 36922 26464 38519
rect 26424 36916 26476 36922
rect 26424 36858 26476 36864
rect 26424 36780 26476 36786
rect 26424 36722 26476 36728
rect 26436 36689 26464 36722
rect 26422 36680 26478 36689
rect 26422 36615 26478 36624
rect 26528 36394 26556 38791
rect 26620 38350 26648 39578
rect 26608 38344 26660 38350
rect 26608 38286 26660 38292
rect 26608 38208 26660 38214
rect 26606 38176 26608 38185
rect 26660 38176 26662 38185
rect 26606 38111 26662 38120
rect 26608 37936 26660 37942
rect 26608 37878 26660 37884
rect 26620 36530 26648 37878
rect 26712 36689 26740 41919
rect 26698 36680 26754 36689
rect 26698 36615 26754 36624
rect 26620 36502 26740 36530
rect 26436 36366 26556 36394
rect 26606 36408 26662 36417
rect 26332 35488 26384 35494
rect 26332 35430 26384 35436
rect 25776 35388 26084 35408
rect 25776 35386 25782 35388
rect 25838 35386 25862 35388
rect 25918 35386 25942 35388
rect 25998 35386 26022 35388
rect 26078 35386 26084 35388
rect 25838 35334 25840 35386
rect 26020 35334 26022 35386
rect 25776 35332 25782 35334
rect 25838 35332 25862 35334
rect 25918 35332 25942 35334
rect 25998 35332 26022 35334
rect 26078 35332 26084 35334
rect 25776 35312 26084 35332
rect 26332 35148 26384 35154
rect 26332 35090 26384 35096
rect 26240 34536 26292 34542
rect 26240 34478 26292 34484
rect 25776 34300 26084 34320
rect 25776 34298 25782 34300
rect 25838 34298 25862 34300
rect 25918 34298 25942 34300
rect 25998 34298 26022 34300
rect 26078 34298 26084 34300
rect 25838 34246 25840 34298
rect 26020 34246 26022 34298
rect 25776 34244 25782 34246
rect 25838 34244 25862 34246
rect 25918 34244 25942 34246
rect 25998 34244 26022 34246
rect 26078 34244 26084 34246
rect 25776 34224 26084 34244
rect 25596 34128 25648 34134
rect 25964 34128 26016 34134
rect 25596 34070 25648 34076
rect 25778 34096 25834 34105
rect 25964 34070 26016 34076
rect 25778 34031 25834 34040
rect 25792 33998 25820 34031
rect 25780 33992 25832 33998
rect 25780 33934 25832 33940
rect 25688 33924 25740 33930
rect 25688 33866 25740 33872
rect 25596 32768 25648 32774
rect 25596 32710 25648 32716
rect 25608 31890 25636 32710
rect 25596 31884 25648 31890
rect 25596 31826 25648 31832
rect 25594 31784 25650 31793
rect 25594 31719 25650 31728
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25608 31226 25636 31719
rect 25516 31198 25636 31226
rect 25412 30728 25464 30734
rect 25412 30670 25464 30676
rect 25412 30252 25464 30258
rect 25412 30194 25464 30200
rect 25424 27606 25452 30194
rect 25412 27600 25464 27606
rect 25412 27542 25464 27548
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25424 27169 25452 27406
rect 25410 27160 25466 27169
rect 25410 27095 25466 27104
rect 25412 26988 25464 26994
rect 25412 26930 25464 26936
rect 25424 26466 25452 26930
rect 25516 26874 25544 31198
rect 25596 31136 25648 31142
rect 25596 31078 25648 31084
rect 25608 30938 25636 31078
rect 25596 30932 25648 30938
rect 25596 30874 25648 30880
rect 25596 30796 25648 30802
rect 25596 30738 25648 30744
rect 25608 30190 25636 30738
rect 25596 30184 25648 30190
rect 25594 30152 25596 30161
rect 25648 30152 25650 30161
rect 25594 30087 25650 30096
rect 25596 30048 25648 30054
rect 25596 29990 25648 29996
rect 25608 29714 25636 29990
rect 25700 29850 25728 33866
rect 25872 33584 25924 33590
rect 25872 33526 25924 33532
rect 25884 33386 25912 33526
rect 25976 33454 26004 34070
rect 26252 33658 26280 34478
rect 26240 33652 26292 33658
rect 26240 33594 26292 33600
rect 26148 33584 26200 33590
rect 26148 33526 26200 33532
rect 25964 33448 26016 33454
rect 25964 33390 26016 33396
rect 25872 33380 25924 33386
rect 25872 33322 25924 33328
rect 25776 33212 26084 33232
rect 25776 33210 25782 33212
rect 25838 33210 25862 33212
rect 25918 33210 25942 33212
rect 25998 33210 26022 33212
rect 26078 33210 26084 33212
rect 25838 33158 25840 33210
rect 26020 33158 26022 33210
rect 25776 33156 25782 33158
rect 25838 33156 25862 33158
rect 25918 33156 25942 33158
rect 25998 33156 26022 33158
rect 26078 33156 26084 33158
rect 25776 33136 26084 33156
rect 25780 33040 25832 33046
rect 25778 33008 25780 33017
rect 25832 33008 25834 33017
rect 25778 32943 25834 32952
rect 25872 32904 25924 32910
rect 25872 32846 25924 32852
rect 25884 32366 25912 32846
rect 25872 32360 25924 32366
rect 25872 32302 25924 32308
rect 25776 32124 26084 32144
rect 25776 32122 25782 32124
rect 25838 32122 25862 32124
rect 25918 32122 25942 32124
rect 25998 32122 26022 32124
rect 26078 32122 26084 32124
rect 25838 32070 25840 32122
rect 26020 32070 26022 32122
rect 25776 32068 25782 32070
rect 25838 32068 25862 32070
rect 25918 32068 25942 32070
rect 25998 32068 26022 32070
rect 26078 32068 26084 32070
rect 25776 32048 26084 32068
rect 26056 31952 26108 31958
rect 26054 31920 26056 31929
rect 26108 31920 26110 31929
rect 26054 31855 26110 31864
rect 26160 31385 26188 33526
rect 26344 33318 26372 35090
rect 26332 33312 26384 33318
rect 26332 33254 26384 33260
rect 26332 32428 26384 32434
rect 26332 32370 26384 32376
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 26252 31822 26280 32166
rect 26240 31816 26292 31822
rect 26240 31758 26292 31764
rect 26238 31648 26294 31657
rect 26238 31583 26294 31592
rect 26146 31376 26202 31385
rect 26146 31311 26202 31320
rect 26148 31204 26200 31210
rect 26148 31146 26200 31152
rect 25776 31036 26084 31056
rect 25776 31034 25782 31036
rect 25838 31034 25862 31036
rect 25918 31034 25942 31036
rect 25998 31034 26022 31036
rect 26078 31034 26084 31036
rect 25838 30982 25840 31034
rect 26020 30982 26022 31034
rect 25776 30980 25782 30982
rect 25838 30980 25862 30982
rect 25918 30980 25942 30982
rect 25998 30980 26022 30982
rect 26078 30980 26084 30982
rect 25776 30960 26084 30980
rect 26160 30938 26188 31146
rect 26148 30932 26200 30938
rect 26148 30874 26200 30880
rect 26054 30832 26110 30841
rect 26054 30767 26110 30776
rect 26068 30172 26096 30767
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26160 30326 26188 30670
rect 26148 30320 26200 30326
rect 26148 30262 26200 30268
rect 26068 30144 26188 30172
rect 25776 29948 26084 29968
rect 25776 29946 25782 29948
rect 25838 29946 25862 29948
rect 25918 29946 25942 29948
rect 25998 29946 26022 29948
rect 26078 29946 26084 29948
rect 25838 29894 25840 29946
rect 26020 29894 26022 29946
rect 25776 29892 25782 29894
rect 25838 29892 25862 29894
rect 25918 29892 25942 29894
rect 25998 29892 26022 29894
rect 26078 29892 26084 29894
rect 25776 29872 26084 29892
rect 25688 29844 25740 29850
rect 25688 29786 25740 29792
rect 25964 29776 26016 29782
rect 25778 29744 25834 29753
rect 25596 29708 25648 29714
rect 25964 29718 26016 29724
rect 25778 29679 25834 29688
rect 25596 29650 25648 29656
rect 25596 29232 25648 29238
rect 25596 29174 25648 29180
rect 25608 28218 25636 29174
rect 25792 28948 25820 29679
rect 25872 29640 25924 29646
rect 25872 29582 25924 29588
rect 25884 29510 25912 29582
rect 25872 29504 25924 29510
rect 25976 29481 26004 29718
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 25872 29446 25924 29452
rect 25962 29472 26018 29481
rect 25962 29407 26018 29416
rect 26068 29345 26096 29514
rect 26054 29336 26110 29345
rect 26054 29271 26110 29280
rect 26054 29200 26110 29209
rect 26054 29135 26056 29144
rect 26108 29135 26110 29144
rect 26056 29106 26108 29112
rect 25700 28920 25820 28948
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25594 27976 25650 27985
rect 25594 27911 25650 27920
rect 25608 27062 25636 27911
rect 25596 27056 25648 27062
rect 25700 27033 25728 28920
rect 25776 28860 26084 28880
rect 25776 28858 25782 28860
rect 25838 28858 25862 28860
rect 25918 28858 25942 28860
rect 25998 28858 26022 28860
rect 26078 28858 26084 28860
rect 25838 28806 25840 28858
rect 26020 28806 26022 28858
rect 25776 28804 25782 28806
rect 25838 28804 25862 28806
rect 25918 28804 25942 28806
rect 25998 28804 26022 28806
rect 26078 28804 26084 28806
rect 25776 28784 26084 28804
rect 25776 27772 26084 27792
rect 25776 27770 25782 27772
rect 25838 27770 25862 27772
rect 25918 27770 25942 27772
rect 25998 27770 26022 27772
rect 26078 27770 26084 27772
rect 25838 27718 25840 27770
rect 26020 27718 26022 27770
rect 25776 27716 25782 27718
rect 25838 27716 25862 27718
rect 25918 27716 25942 27718
rect 25998 27716 26022 27718
rect 26078 27716 26084 27718
rect 25776 27696 26084 27716
rect 25780 27600 25832 27606
rect 26160 27554 26188 30144
rect 25780 27542 25832 27548
rect 25792 27470 25820 27542
rect 26068 27526 26188 27554
rect 25780 27464 25832 27470
rect 25780 27406 25832 27412
rect 25872 27056 25924 27062
rect 25596 26998 25648 27004
rect 25686 27024 25742 27033
rect 25872 26998 25924 27004
rect 25686 26959 25742 26968
rect 25516 26846 25728 26874
rect 25884 26858 25912 26998
rect 26068 26858 26096 27526
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 25424 26438 25636 26466
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25516 25498 25544 26250
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25332 25350 25544 25378
rect 25318 25256 25374 25265
rect 25318 25191 25374 25200
rect 25332 24750 25360 25191
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25332 23322 25360 24686
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25424 23866 25452 24142
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 25320 23316 25372 23322
rect 25320 23258 25372 23264
rect 25424 23202 25452 23598
rect 25332 23174 25452 23202
rect 25332 22982 25360 23174
rect 25412 23112 25464 23118
rect 25410 23080 25412 23089
rect 25464 23080 25466 23089
rect 25410 23015 25466 23024
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25332 22030 25360 22374
rect 25320 22024 25372 22030
rect 25320 21966 25372 21972
rect 25318 21856 25374 21865
rect 25318 21791 25374 21800
rect 25332 18465 25360 21791
rect 25424 21690 25452 22578
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25424 19446 25452 21490
rect 25516 19786 25544 25350
rect 25608 22545 25636 26438
rect 25594 22536 25650 22545
rect 25594 22471 25650 22480
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25608 21962 25636 22374
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25608 20942 25636 21558
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25700 19530 25728 26846
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 26056 26852 26108 26858
rect 26056 26794 26108 26800
rect 25776 26684 26084 26704
rect 25776 26682 25782 26684
rect 25838 26682 25862 26684
rect 25918 26682 25942 26684
rect 25998 26682 26022 26684
rect 26078 26682 26084 26684
rect 25838 26630 25840 26682
rect 26020 26630 26022 26682
rect 25776 26628 25782 26630
rect 25838 26628 25862 26630
rect 25918 26628 25942 26630
rect 25998 26628 26022 26630
rect 26078 26628 26084 26630
rect 25776 26608 26084 26628
rect 26054 26480 26110 26489
rect 26054 26415 26110 26424
rect 26068 25684 26096 26415
rect 26160 26382 26188 27406
rect 26252 27130 26280 31583
rect 26344 31346 26372 32370
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 26332 31136 26384 31142
rect 26332 31078 26384 31084
rect 26344 30666 26372 31078
rect 26332 30660 26384 30666
rect 26332 30602 26384 30608
rect 26332 30320 26384 30326
rect 26332 30262 26384 30268
rect 26344 29510 26372 30262
rect 26332 29504 26384 29510
rect 26332 29446 26384 29452
rect 26240 27124 26292 27130
rect 26240 27066 26292 27072
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26252 26489 26280 26726
rect 26238 26480 26294 26489
rect 26238 26415 26294 26424
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26068 25656 26188 25684
rect 25776 25596 26084 25616
rect 25776 25594 25782 25596
rect 25838 25594 25862 25596
rect 25918 25594 25942 25596
rect 25998 25594 26022 25596
rect 26078 25594 26084 25596
rect 25838 25542 25840 25594
rect 26020 25542 26022 25594
rect 25776 25540 25782 25542
rect 25838 25540 25862 25542
rect 25918 25540 25942 25542
rect 25998 25540 26022 25542
rect 26078 25540 26084 25542
rect 25776 25520 26084 25540
rect 25776 24508 26084 24528
rect 25776 24506 25782 24508
rect 25838 24506 25862 24508
rect 25918 24506 25942 24508
rect 25998 24506 26022 24508
rect 26078 24506 26084 24508
rect 25838 24454 25840 24506
rect 26020 24454 26022 24506
rect 25776 24452 25782 24454
rect 25838 24452 25862 24454
rect 25918 24452 25942 24454
rect 25998 24452 26022 24454
rect 26078 24452 26084 24454
rect 25776 24432 26084 24452
rect 25776 23420 26084 23440
rect 25776 23418 25782 23420
rect 25838 23418 25862 23420
rect 25918 23418 25942 23420
rect 25998 23418 26022 23420
rect 26078 23418 26084 23420
rect 25838 23366 25840 23418
rect 26020 23366 26022 23418
rect 25776 23364 25782 23366
rect 25838 23364 25862 23366
rect 25918 23364 25942 23366
rect 25998 23364 26022 23366
rect 26078 23364 26084 23366
rect 25776 23344 26084 23364
rect 26160 23118 26188 25656
rect 26252 24818 26280 26318
rect 26344 25362 26372 29446
rect 26332 25356 26384 25362
rect 26332 25298 26384 25304
rect 26332 25152 26384 25158
rect 26332 25094 26384 25100
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 26238 24712 26294 24721
rect 26238 24647 26294 24656
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25776 22332 26084 22352
rect 25776 22330 25782 22332
rect 25838 22330 25862 22332
rect 25918 22330 25942 22332
rect 25998 22330 26022 22332
rect 26078 22330 26084 22332
rect 25838 22278 25840 22330
rect 26020 22278 26022 22330
rect 25776 22276 25782 22278
rect 25838 22276 25862 22278
rect 25918 22276 25942 22278
rect 25998 22276 26022 22278
rect 26078 22276 26084 22278
rect 25776 22256 26084 22276
rect 26160 22080 26188 23054
rect 26252 22642 26280 24647
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26252 22234 26280 22578
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 25976 22052 26188 22080
rect 26238 22128 26294 22137
rect 26238 22063 26240 22072
rect 25976 21622 26004 22052
rect 26292 22063 26294 22072
rect 26240 22034 26292 22040
rect 26148 21956 26200 21962
rect 26148 21898 26200 21904
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 25964 21616 26016 21622
rect 25964 21558 26016 21564
rect 26068 21332 26096 21626
rect 26160 21570 26188 21898
rect 26252 21690 26280 22034
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26160 21542 26280 21570
rect 26068 21304 26188 21332
rect 25776 21244 26084 21264
rect 25776 21242 25782 21244
rect 25838 21242 25862 21244
rect 25918 21242 25942 21244
rect 25998 21242 26022 21244
rect 26078 21242 26084 21244
rect 25838 21190 25840 21242
rect 26020 21190 26022 21242
rect 25776 21188 25782 21190
rect 25838 21188 25862 21190
rect 25918 21188 25942 21190
rect 25998 21188 26022 21190
rect 26078 21188 26084 21190
rect 25776 21168 26084 21188
rect 25778 21040 25834 21049
rect 25778 20975 25834 20984
rect 25792 20330 25820 20975
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25776 20156 26084 20176
rect 25776 20154 25782 20156
rect 25838 20154 25862 20156
rect 25918 20154 25942 20156
rect 25998 20154 26022 20156
rect 26078 20154 26084 20156
rect 25838 20102 25840 20154
rect 26020 20102 26022 20154
rect 25776 20100 25782 20102
rect 25838 20100 25862 20102
rect 25918 20100 25942 20102
rect 25998 20100 26022 20102
rect 26078 20100 26084 20102
rect 25776 20080 26084 20100
rect 26160 20040 26188 21304
rect 25976 20012 26188 20040
rect 25976 19922 26004 20012
rect 25964 19916 26016 19922
rect 25516 19502 25728 19530
rect 25884 19876 25964 19904
rect 25412 19440 25464 19446
rect 25412 19382 25464 19388
rect 25412 18896 25464 18902
rect 25412 18838 25464 18844
rect 25318 18456 25374 18465
rect 25318 18391 25374 18400
rect 25240 18278 25360 18306
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 25044 16516 25096 16522
rect 25044 16458 25096 16464
rect 25042 16144 25098 16153
rect 25042 16079 25044 16088
rect 25096 16079 25098 16088
rect 25044 16050 25096 16056
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25056 12646 25084 14758
rect 25148 14226 25176 18158
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 16998 25268 18022
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25240 15094 25268 16050
rect 25228 15088 25280 15094
rect 25228 15030 25280 15036
rect 25332 14414 25360 18278
rect 25424 18154 25452 18838
rect 25412 18148 25464 18154
rect 25412 18090 25464 18096
rect 25516 17218 25544 19502
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25608 17678 25636 19314
rect 25792 19258 25820 19314
rect 25700 19230 25820 19258
rect 25884 19242 25912 19876
rect 25964 19858 26016 19864
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 26068 19258 26096 19858
rect 25872 19236 25924 19242
rect 25700 18850 25728 19230
rect 26068 19230 26188 19258
rect 25872 19178 25924 19184
rect 25776 19068 26084 19088
rect 25776 19066 25782 19068
rect 25838 19066 25862 19068
rect 25918 19066 25942 19068
rect 25998 19066 26022 19068
rect 26078 19066 26084 19068
rect 25838 19014 25840 19066
rect 26020 19014 26022 19066
rect 25776 19012 25782 19014
rect 25838 19012 25862 19014
rect 25918 19012 25942 19014
rect 25998 19012 26022 19014
rect 26078 19012 26084 19014
rect 25776 18992 26084 19012
rect 25700 18822 25820 18850
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25700 17882 25728 18634
rect 25792 18193 25820 18822
rect 25962 18728 26018 18737
rect 25962 18663 25964 18672
rect 26016 18663 26018 18672
rect 25964 18634 26016 18640
rect 25976 18222 26004 18634
rect 25964 18216 26016 18222
rect 25778 18184 25834 18193
rect 25964 18158 26016 18164
rect 25778 18119 25834 18128
rect 25776 17980 26084 18000
rect 25776 17978 25782 17980
rect 25838 17978 25862 17980
rect 25918 17978 25942 17980
rect 25998 17978 26022 17980
rect 26078 17978 26084 17980
rect 25838 17926 25840 17978
rect 26020 17926 26022 17978
rect 25776 17924 25782 17926
rect 25838 17924 25862 17926
rect 25918 17924 25942 17926
rect 25998 17924 26022 17926
rect 26078 17924 26084 17926
rect 25776 17904 26084 17924
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25596 17672 25648 17678
rect 26056 17672 26108 17678
rect 25596 17614 25648 17620
rect 26054 17640 26056 17649
rect 26108 17640 26110 17649
rect 26054 17575 26110 17584
rect 25516 17190 25728 17218
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25412 15428 25464 15434
rect 25412 15370 25464 15376
rect 25424 15162 25452 15370
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 25424 14822 25452 14962
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25148 14198 25360 14226
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 25056 12102 25084 12582
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 11694 25084 12038
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 25148 11218 25176 13330
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25148 10810 25176 11154
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24952 5092 25004 5098
rect 24952 5034 25004 5040
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 25056 2378 25084 8434
rect 25240 7750 25268 13874
rect 25332 11150 25360 14198
rect 25424 13326 25452 14554
rect 25516 13938 25544 16458
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25608 15502 25636 16050
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25594 15328 25650 15337
rect 25594 15263 25650 15272
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25412 12980 25464 12986
rect 25412 12922 25464 12928
rect 25424 12850 25452 12922
rect 25516 12850 25544 13126
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25332 9382 25360 11086
rect 25424 11082 25452 11630
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25516 9994 25544 11494
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25332 8974 25360 9318
rect 25320 8968 25372 8974
rect 25320 8910 25372 8916
rect 25516 8650 25544 9930
rect 25608 9586 25636 15263
rect 25700 11082 25728 17190
rect 25776 16892 26084 16912
rect 25776 16890 25782 16892
rect 25838 16890 25862 16892
rect 25918 16890 25942 16892
rect 25998 16890 26022 16892
rect 26078 16890 26084 16892
rect 25838 16838 25840 16890
rect 26020 16838 26022 16890
rect 25776 16836 25782 16838
rect 25838 16836 25862 16838
rect 25918 16836 25942 16838
rect 25998 16836 26022 16838
rect 26078 16836 26084 16838
rect 25776 16816 26084 16836
rect 26160 15978 26188 19230
rect 26252 17678 26280 21542
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 26148 15972 26200 15978
rect 26148 15914 26200 15920
rect 25776 15804 26084 15824
rect 25776 15802 25782 15804
rect 25838 15802 25862 15804
rect 25918 15802 25942 15804
rect 25998 15802 26022 15804
rect 26078 15802 26084 15804
rect 25838 15750 25840 15802
rect 26020 15750 26022 15802
rect 25776 15748 25782 15750
rect 25838 15748 25862 15750
rect 25918 15748 25942 15750
rect 25998 15748 26022 15750
rect 26078 15748 26084 15750
rect 25776 15728 26084 15748
rect 26252 15502 26280 16118
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 25776 14716 26084 14736
rect 25776 14714 25782 14716
rect 25838 14714 25862 14716
rect 25918 14714 25942 14716
rect 25998 14714 26022 14716
rect 26078 14714 26084 14716
rect 25838 14662 25840 14714
rect 26020 14662 26022 14714
rect 25776 14660 25782 14662
rect 25838 14660 25862 14662
rect 25918 14660 25942 14662
rect 25998 14660 26022 14662
rect 26078 14660 26084 14662
rect 25776 14640 26084 14660
rect 26160 14414 26188 15438
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25792 14113 25820 14214
rect 25778 14104 25834 14113
rect 25778 14039 25834 14048
rect 26160 13870 26188 14350
rect 26252 14006 26280 15438
rect 26344 14822 26372 25094
rect 26436 20874 26464 36366
rect 26606 36343 26662 36352
rect 26516 36304 26568 36310
rect 26514 36272 26516 36281
rect 26568 36272 26570 36281
rect 26514 36207 26570 36216
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 26528 27538 26556 35430
rect 26516 27532 26568 27538
rect 26516 27474 26568 27480
rect 26516 27396 26568 27402
rect 26516 27338 26568 27344
rect 26424 20868 26476 20874
rect 26424 20810 26476 20816
rect 26422 20768 26478 20777
rect 26422 20703 26478 20712
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26240 14000 26292 14006
rect 26240 13942 26292 13948
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 25776 13628 26084 13648
rect 25776 13626 25782 13628
rect 25838 13626 25862 13628
rect 25918 13626 25942 13628
rect 25998 13626 26022 13628
rect 26078 13626 26084 13628
rect 25838 13574 25840 13626
rect 26020 13574 26022 13626
rect 25776 13572 25782 13574
rect 25838 13572 25862 13574
rect 25918 13572 25942 13574
rect 25998 13572 26022 13574
rect 26078 13572 26084 13574
rect 25776 13552 26084 13572
rect 26160 13326 26188 13806
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26252 13394 26280 13738
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 25776 12540 26084 12560
rect 25776 12538 25782 12540
rect 25838 12538 25862 12540
rect 25918 12538 25942 12540
rect 25998 12538 26022 12540
rect 26078 12538 26084 12540
rect 25838 12486 25840 12538
rect 26020 12486 26022 12538
rect 25776 12484 25782 12486
rect 25838 12484 25862 12486
rect 25918 12484 25942 12486
rect 25998 12484 26022 12486
rect 26078 12484 26084 12486
rect 25776 12464 26084 12484
rect 26160 12238 26188 13262
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 25964 12164 26016 12170
rect 25964 12106 26016 12112
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25884 11626 25912 12038
rect 25976 11762 26004 12106
rect 26146 12064 26202 12073
rect 26146 11999 26202 12008
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25872 11620 25924 11626
rect 25872 11562 25924 11568
rect 25776 11452 26084 11472
rect 25776 11450 25782 11452
rect 25838 11450 25862 11452
rect 25918 11450 25942 11452
rect 25998 11450 26022 11452
rect 26078 11450 26084 11452
rect 25838 11398 25840 11450
rect 26020 11398 26022 11450
rect 25776 11396 25782 11398
rect 25838 11396 25862 11398
rect 25918 11396 25942 11398
rect 25998 11396 26022 11398
rect 26078 11396 26084 11398
rect 25776 11376 26084 11396
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25776 10364 26084 10384
rect 25776 10362 25782 10364
rect 25838 10362 25862 10364
rect 25918 10362 25942 10364
rect 25998 10362 26022 10364
rect 26078 10362 26084 10364
rect 25838 10310 25840 10362
rect 26020 10310 26022 10362
rect 25776 10308 25782 10310
rect 25838 10308 25862 10310
rect 25918 10308 25942 10310
rect 25998 10308 26022 10310
rect 26078 10308 26084 10310
rect 25776 10288 26084 10308
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25332 8622 25544 8650
rect 25228 7744 25280 7750
rect 25228 7686 25280 7692
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 4622 25268 7142
rect 25332 6746 25360 8622
rect 25608 8566 25636 9522
rect 25776 9276 26084 9296
rect 25776 9274 25782 9276
rect 25838 9274 25862 9276
rect 25918 9274 25942 9276
rect 25998 9274 26022 9276
rect 26078 9274 26084 9276
rect 25838 9222 25840 9274
rect 26020 9222 26022 9274
rect 25776 9220 25782 9222
rect 25838 9220 25862 9222
rect 25918 9220 25942 9222
rect 25998 9220 26022 9222
rect 26078 9220 26084 9222
rect 25776 9200 26084 9220
rect 26160 8906 26188 11999
rect 26252 11898 26280 13194
rect 26344 12986 26372 14758
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26240 11892 26292 11898
rect 26240 11834 26292 11840
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26252 9994 26280 11018
rect 26344 10266 26372 12786
rect 26436 12442 26464 20703
rect 26528 19825 26556 27338
rect 26514 19816 26570 19825
rect 26514 19751 26570 19760
rect 26514 19680 26570 19689
rect 26514 19615 26570 19624
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26528 11200 26556 19615
rect 26620 18986 26648 36343
rect 26712 34202 26740 36502
rect 26700 34196 26752 34202
rect 26700 34138 26752 34144
rect 26700 34060 26752 34066
rect 26700 34002 26752 34008
rect 26712 31498 26740 34002
rect 26804 31686 26832 48447
rect 26882 48328 26938 48337
rect 26882 48263 26938 48272
rect 26896 46170 26924 48263
rect 26884 46164 26936 46170
rect 26884 46106 26936 46112
rect 26884 44736 26936 44742
rect 26884 44678 26936 44684
rect 26896 44402 26924 44678
rect 26884 44396 26936 44402
rect 26884 44338 26936 44344
rect 26896 43790 26924 44338
rect 26884 43784 26936 43790
rect 26884 43726 26936 43732
rect 26896 41585 26924 43726
rect 26882 41576 26938 41585
rect 26882 41511 26938 41520
rect 26988 41414 27016 48606
rect 27066 48583 27122 48592
rect 27066 48512 27122 48521
rect 27066 48447 27122 48456
rect 26896 41386 27016 41414
rect 26896 37108 26924 41386
rect 26974 41168 27030 41177
rect 26974 41103 27030 41112
rect 26988 37874 27016 41103
rect 26976 37868 27028 37874
rect 26976 37810 27028 37816
rect 26988 37398 27016 37810
rect 26976 37392 27028 37398
rect 26976 37334 27028 37340
rect 27080 37346 27108 48447
rect 27356 48226 27384 48878
rect 27448 48736 27476 49166
rect 27540 49094 27568 52566
rect 27618 52527 27674 52536
rect 27618 52456 27674 52465
rect 27618 52391 27674 52400
rect 27632 51610 27660 52391
rect 27724 52018 27752 52906
rect 27712 52012 27764 52018
rect 27712 51954 27764 51960
rect 27620 51604 27672 51610
rect 27620 51546 27672 51552
rect 27816 51338 27844 60046
rect 27908 53825 27936 60959
rect 28000 60636 28028 66098
rect 28080 65952 28132 65958
rect 28080 65894 28132 65900
rect 28172 65952 28224 65958
rect 28172 65894 28224 65900
rect 28092 65521 28120 65894
rect 28078 65512 28134 65521
rect 28078 65447 28134 65456
rect 28080 65000 28132 65006
rect 28078 64968 28080 64977
rect 28132 64968 28134 64977
rect 28078 64903 28134 64912
rect 28184 64161 28212 65894
rect 28170 64152 28226 64161
rect 28170 64087 28226 64096
rect 28276 64025 28304 67186
rect 28460 65657 28488 69362
rect 28446 65648 28502 65657
rect 28446 65583 28502 65592
rect 28448 65476 28500 65482
rect 28448 65418 28500 65424
rect 28356 65408 28408 65414
rect 28356 65350 28408 65356
rect 28368 65074 28396 65350
rect 28356 65068 28408 65074
rect 28356 65010 28408 65016
rect 28356 64932 28408 64938
rect 28356 64874 28408 64880
rect 28368 64326 28396 64874
rect 28356 64320 28408 64326
rect 28356 64262 28408 64268
rect 28262 64016 28318 64025
rect 28172 63980 28224 63986
rect 28368 63986 28396 64262
rect 28262 63951 28318 63960
rect 28356 63980 28408 63986
rect 28172 63922 28224 63928
rect 28356 63922 28408 63928
rect 28080 63912 28132 63918
rect 28078 63880 28080 63889
rect 28132 63880 28134 63889
rect 28078 63815 28134 63824
rect 28080 63504 28132 63510
rect 28080 63446 28132 63452
rect 28092 62762 28120 63446
rect 28080 62756 28132 62762
rect 28080 62698 28132 62704
rect 28092 61033 28120 62698
rect 28078 61024 28134 61033
rect 28078 60959 28134 60968
rect 28000 60608 28120 60636
rect 28092 60568 28120 60608
rect 28000 60540 28120 60568
rect 27894 53816 27950 53825
rect 27894 53751 27950 53760
rect 28000 53666 28028 60540
rect 28078 60208 28134 60217
rect 28078 60143 28134 60152
rect 28092 60042 28120 60143
rect 28080 60036 28132 60042
rect 28080 59978 28132 59984
rect 28078 59664 28134 59673
rect 28078 59599 28080 59608
rect 28132 59599 28134 59608
rect 28080 59570 28132 59576
rect 28078 59528 28134 59537
rect 28078 59463 28134 59472
rect 27908 53638 28028 53666
rect 27908 53242 27936 53638
rect 27988 53576 28040 53582
rect 27988 53518 28040 53524
rect 27896 53236 27948 53242
rect 27896 53178 27948 53184
rect 27896 53100 27948 53106
rect 27896 53042 27948 53048
rect 27620 51332 27672 51338
rect 27620 51274 27672 51280
rect 27804 51332 27856 51338
rect 27804 51274 27856 51280
rect 27632 49434 27660 51274
rect 27802 51232 27858 51241
rect 27802 51167 27858 51176
rect 27710 51096 27766 51105
rect 27710 51031 27766 51040
rect 27620 49428 27672 49434
rect 27620 49370 27672 49376
rect 27528 49088 27580 49094
rect 27528 49030 27580 49036
rect 27620 49088 27672 49094
rect 27620 49030 27672 49036
rect 27632 48793 27660 49030
rect 27618 48784 27674 48793
rect 27528 48748 27580 48754
rect 27448 48708 27528 48736
rect 27618 48719 27674 48728
rect 27528 48690 27580 48696
rect 27434 48512 27490 48521
rect 27434 48447 27490 48456
rect 27283 48198 27384 48226
rect 27283 48192 27311 48198
rect 27172 48164 27311 48192
rect 27172 47122 27200 48164
rect 27250 48104 27306 48113
rect 27250 48039 27306 48048
rect 27264 47598 27292 48039
rect 27342 47968 27398 47977
rect 27342 47903 27398 47912
rect 27252 47592 27304 47598
rect 27252 47534 27304 47540
rect 27264 47190 27292 47534
rect 27252 47184 27304 47190
rect 27252 47126 27304 47132
rect 27160 47116 27212 47122
rect 27160 47058 27212 47064
rect 27172 44878 27200 47058
rect 27252 46164 27304 46170
rect 27252 46106 27304 46112
rect 27160 44872 27212 44878
rect 27160 44814 27212 44820
rect 27160 44532 27212 44538
rect 27160 44474 27212 44480
rect 27172 37466 27200 44474
rect 27264 38010 27292 46106
rect 27252 38004 27304 38010
rect 27252 37946 27304 37952
rect 27160 37460 27212 37466
rect 27160 37402 27212 37408
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 26988 37244 27016 37334
rect 27080 37318 27200 37346
rect 26988 37216 27108 37244
rect 26896 37080 27016 37108
rect 26884 36644 26936 36650
rect 26884 36586 26936 36592
rect 26896 36378 26924 36586
rect 26884 36372 26936 36378
rect 26884 36314 26936 36320
rect 26884 36168 26936 36174
rect 26884 36110 26936 36116
rect 26896 34406 26924 36110
rect 26884 34400 26936 34406
rect 26884 34342 26936 34348
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26896 33590 26924 33934
rect 26884 33584 26936 33590
rect 26884 33526 26936 33532
rect 26896 32910 26924 33526
rect 26884 32904 26936 32910
rect 26884 32846 26936 32852
rect 26988 32201 27016 37080
rect 27080 35086 27108 37216
rect 27068 35080 27120 35086
rect 27068 35022 27120 35028
rect 27068 34604 27120 34610
rect 27068 34546 27120 34552
rect 26974 32192 27030 32201
rect 26974 32127 27030 32136
rect 27080 31940 27108 34546
rect 27172 34474 27200 37318
rect 27160 34468 27212 34474
rect 27160 34410 27212 34416
rect 27264 34082 27292 37402
rect 27172 34054 27292 34082
rect 27172 33561 27200 34054
rect 27252 33924 27304 33930
rect 27252 33866 27304 33872
rect 27158 33552 27214 33561
rect 27158 33487 27214 33496
rect 27160 33448 27212 33454
rect 27160 33390 27212 33396
rect 26896 31912 27108 31940
rect 26792 31680 26844 31686
rect 26792 31622 26844 31628
rect 26712 31470 26832 31498
rect 26700 31340 26752 31346
rect 26700 31282 26752 31288
rect 26712 27674 26740 31282
rect 26804 30433 26832 31470
rect 26790 30424 26846 30433
rect 26790 30359 26846 30368
rect 26792 30116 26844 30122
rect 26792 30058 26844 30064
rect 26804 29850 26832 30058
rect 26792 29844 26844 29850
rect 26792 29786 26844 29792
rect 26790 29744 26846 29753
rect 26790 29679 26846 29688
rect 26804 28490 26832 29679
rect 26792 28484 26844 28490
rect 26792 28426 26844 28432
rect 26792 28144 26844 28150
rect 26792 28086 26844 28092
rect 26700 27668 26752 27674
rect 26700 27610 26752 27616
rect 26700 27532 26752 27538
rect 26700 27474 26752 27480
rect 26712 26042 26740 27474
rect 26700 26036 26752 26042
rect 26700 25978 26752 25984
rect 26700 25288 26752 25294
rect 26804 25265 26832 28086
rect 26896 26926 26924 31912
rect 26974 31784 27030 31793
rect 26974 31719 27030 31728
rect 27068 31748 27120 31754
rect 26988 31482 27016 31719
rect 27068 31690 27120 31696
rect 26976 31476 27028 31482
rect 26976 31418 27028 31424
rect 27080 31346 27108 31690
rect 26976 31340 27028 31346
rect 26976 31282 27028 31288
rect 27068 31340 27120 31346
rect 27068 31282 27120 31288
rect 26988 31226 27016 31282
rect 26988 31198 27108 31226
rect 27080 30734 27108 31198
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 27080 29889 27108 30670
rect 27066 29880 27122 29889
rect 27066 29815 27122 29824
rect 27172 29730 27200 33390
rect 27264 31890 27292 33866
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 27264 31498 27292 31826
rect 27356 31754 27384 47903
rect 27448 44538 27476 48447
rect 27540 48142 27568 48690
rect 27618 48328 27674 48337
rect 27618 48263 27674 48272
rect 27528 48136 27580 48142
rect 27528 48078 27580 48084
rect 27540 47598 27568 48078
rect 27528 47592 27580 47598
rect 27528 47534 27580 47540
rect 27540 47054 27568 47534
rect 27528 47048 27580 47054
rect 27528 46990 27580 46996
rect 27528 46912 27580 46918
rect 27528 46854 27580 46860
rect 27436 44532 27488 44538
rect 27436 44474 27488 44480
rect 27434 44432 27490 44441
rect 27434 44367 27490 44376
rect 27448 42401 27476 44367
rect 27434 42392 27490 42401
rect 27434 42327 27490 42336
rect 27436 42288 27488 42294
rect 27436 42230 27488 42236
rect 27448 42158 27476 42230
rect 27436 42152 27488 42158
rect 27436 42094 27488 42100
rect 27436 42016 27488 42022
rect 27436 41958 27488 41964
rect 27448 41002 27476 41958
rect 27540 41721 27568 46854
rect 27632 42265 27660 48263
rect 27724 42673 27752 51031
rect 27816 46934 27844 51167
rect 27908 50454 27936 53042
rect 28000 52873 28028 53518
rect 27986 52864 28042 52873
rect 27986 52799 28042 52808
rect 27986 52728 28042 52737
rect 27986 52663 28042 52672
rect 28000 52562 28028 52663
rect 27988 52556 28040 52562
rect 27988 52498 28040 52504
rect 27988 52420 28040 52426
rect 27988 52362 28040 52368
rect 28000 50969 28028 52362
rect 27986 50960 28042 50969
rect 27986 50895 28042 50904
rect 27896 50448 27948 50454
rect 27896 50390 27948 50396
rect 27988 50312 28040 50318
rect 27988 50254 28040 50260
rect 27896 50244 27948 50250
rect 27896 50186 27948 50192
rect 27908 49450 27936 50186
rect 28000 49609 28028 50254
rect 27986 49600 28042 49609
rect 27986 49535 28042 49544
rect 27908 49422 28028 49450
rect 27896 49292 27948 49298
rect 27896 49234 27948 49240
rect 27908 48278 27936 49234
rect 27896 48272 27948 48278
rect 27896 48214 27948 48220
rect 27896 48136 27948 48142
rect 27896 48078 27948 48084
rect 27908 47122 27936 48078
rect 27896 47116 27948 47122
rect 27896 47058 27948 47064
rect 27816 46906 27936 46934
rect 27804 45552 27856 45558
rect 27804 45494 27856 45500
rect 27816 44713 27844 45494
rect 27802 44704 27858 44713
rect 27802 44639 27858 44648
rect 27804 43104 27856 43110
rect 27804 43046 27856 43052
rect 27710 42664 27766 42673
rect 27710 42599 27766 42608
rect 27712 42288 27764 42294
rect 27618 42256 27674 42265
rect 27712 42230 27764 42236
rect 27618 42191 27674 42200
rect 27620 42084 27672 42090
rect 27620 42026 27672 42032
rect 27526 41712 27582 41721
rect 27526 41647 27582 41656
rect 27528 41608 27580 41614
rect 27632 41596 27660 42026
rect 27580 41568 27660 41596
rect 27528 41550 27580 41556
rect 27632 41138 27660 41568
rect 27724 41546 27752 42230
rect 27816 42226 27844 43046
rect 27804 42220 27856 42226
rect 27804 42162 27856 42168
rect 27802 41984 27858 41993
rect 27802 41919 27858 41928
rect 27712 41540 27764 41546
rect 27712 41482 27764 41488
rect 27712 41268 27764 41274
rect 27712 41210 27764 41216
rect 27724 41177 27752 41210
rect 27710 41168 27766 41177
rect 27620 41132 27672 41138
rect 27710 41103 27766 41112
rect 27620 41074 27672 41080
rect 27526 41032 27582 41041
rect 27436 40996 27488 41002
rect 27526 40967 27582 40976
rect 27710 41032 27766 41041
rect 27710 40967 27766 40976
rect 27436 40938 27488 40944
rect 27540 40934 27568 40967
rect 27528 40928 27580 40934
rect 27580 40876 27660 40882
rect 27528 40870 27660 40876
rect 27540 40854 27660 40870
rect 27540 40805 27568 40854
rect 27528 40520 27580 40526
rect 27528 40462 27580 40468
rect 27436 40384 27488 40390
rect 27436 40326 27488 40332
rect 27448 40050 27476 40326
rect 27540 40186 27568 40462
rect 27632 40186 27660 40854
rect 27528 40180 27580 40186
rect 27528 40122 27580 40128
rect 27620 40180 27672 40186
rect 27620 40122 27672 40128
rect 27436 40044 27488 40050
rect 27436 39986 27488 39992
rect 27448 36174 27476 39986
rect 27620 39908 27672 39914
rect 27620 39850 27672 39856
rect 27528 39840 27580 39846
rect 27528 39782 27580 39788
rect 27540 39114 27568 39782
rect 27632 39681 27660 39850
rect 27618 39672 27674 39681
rect 27618 39607 27674 39616
rect 27540 39086 27660 39114
rect 27528 38956 27580 38962
rect 27528 38898 27580 38904
rect 27540 37466 27568 38898
rect 27632 38010 27660 39086
rect 27620 38004 27672 38010
rect 27620 37946 27672 37952
rect 27528 37460 27580 37466
rect 27528 37402 27580 37408
rect 27620 37256 27672 37262
rect 27620 37198 27672 37204
rect 27528 37120 27580 37126
rect 27528 37062 27580 37068
rect 27436 36168 27488 36174
rect 27436 36110 27488 36116
rect 27436 36032 27488 36038
rect 27436 35974 27488 35980
rect 27344 31748 27396 31754
rect 27344 31690 27396 31696
rect 27264 31470 27384 31498
rect 27252 31340 27304 31346
rect 27252 31282 27304 31288
rect 26988 29702 27200 29730
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26884 26784 26936 26790
rect 26884 26726 26936 26732
rect 26700 25230 26752 25236
rect 26790 25256 26846 25265
rect 26712 24954 26740 25230
rect 26790 25191 26846 25200
rect 26896 25106 26924 26726
rect 26804 25078 26924 25106
rect 26700 24948 26752 24954
rect 26700 24890 26752 24896
rect 26712 24206 26740 24890
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26712 22982 26740 24006
rect 26700 22976 26752 22982
rect 26700 22918 26752 22924
rect 26698 22808 26754 22817
rect 26698 22743 26754 22752
rect 26712 22710 26740 22743
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 26700 22432 26752 22438
rect 26700 22374 26752 22380
rect 26712 19378 26740 22374
rect 26804 22234 26832 25078
rect 26882 24984 26938 24993
rect 26882 24919 26938 24928
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26790 22128 26846 22137
rect 26790 22063 26846 22072
rect 26804 21554 26832 22063
rect 26896 22001 26924 24919
rect 26882 21992 26938 22001
rect 26882 21927 26938 21936
rect 26792 21548 26844 21554
rect 26792 21490 26844 21496
rect 26884 20868 26936 20874
rect 26884 20810 26936 20816
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26620 18958 26740 18986
rect 26608 18896 26660 18902
rect 26608 18838 26660 18844
rect 26620 17746 26648 18838
rect 26608 17740 26660 17746
rect 26608 17682 26660 17688
rect 26606 17640 26662 17649
rect 26606 17575 26662 17584
rect 26620 16658 26648 17575
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26620 13530 26648 15506
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 26712 13394 26740 18958
rect 26804 14278 26832 19722
rect 26896 15570 26924 20810
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26790 14104 26846 14113
rect 26790 14039 26846 14048
rect 26700 13388 26752 13394
rect 26700 13330 26752 13336
rect 26804 13326 26832 14039
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26700 13252 26752 13258
rect 26700 13194 26752 13200
rect 26712 11626 26740 13194
rect 26804 12374 26832 13262
rect 26792 12368 26844 12374
rect 26792 12310 26844 12316
rect 26700 11620 26752 11626
rect 26700 11562 26752 11568
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26436 11172 26556 11200
rect 26436 10962 26464 11172
rect 26620 11150 26648 11494
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26436 10934 26648 10962
rect 26514 10840 26570 10849
rect 26514 10775 26570 10784
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 26344 9674 26372 10202
rect 26344 9646 26464 9674
rect 26148 8900 26200 8906
rect 26148 8842 26200 8848
rect 26160 8634 26188 8842
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 25596 8560 25648 8566
rect 25516 8508 25596 8514
rect 25516 8502 25648 8508
rect 25516 8486 25636 8502
rect 25516 7954 25544 8486
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25504 7336 25556 7342
rect 25504 7278 25556 7284
rect 25424 6866 25452 7278
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25516 6798 25544 7278
rect 25608 6934 25636 8366
rect 26436 8362 26464 9646
rect 26528 8566 26556 10775
rect 26620 8566 26648 10934
rect 26712 10690 26740 11562
rect 26804 10849 26832 12310
rect 26896 12102 26924 15370
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26790 10840 26846 10849
rect 26790 10775 26846 10784
rect 26712 10674 26832 10690
rect 26712 10668 26844 10674
rect 26712 10662 26792 10668
rect 26792 10610 26844 10616
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 26712 8378 26740 9454
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 26620 8350 26740 8378
rect 25776 8188 26084 8208
rect 25776 8186 25782 8188
rect 25838 8186 25862 8188
rect 25918 8186 25942 8188
rect 25998 8186 26022 8188
rect 26078 8186 26084 8188
rect 25838 8134 25840 8186
rect 26020 8134 26022 8186
rect 25776 8132 25782 8134
rect 25838 8132 25862 8134
rect 25918 8132 25942 8134
rect 25998 8132 26022 8134
rect 26078 8132 26084 8134
rect 25776 8112 26084 8132
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 25700 7410 25728 7822
rect 25964 7812 26016 7818
rect 25964 7754 26016 7760
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25596 6928 25648 6934
rect 25596 6870 25648 6876
rect 25504 6792 25556 6798
rect 25332 6718 25452 6746
rect 25504 6734 25556 6740
rect 25320 5568 25372 5574
rect 25320 5510 25372 5516
rect 25332 4690 25360 5510
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25424 4622 25452 6718
rect 25516 5710 25544 6734
rect 25700 6662 25728 7346
rect 25976 7274 26004 7754
rect 26068 7342 26096 7822
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 25964 7268 26016 7274
rect 25964 7210 26016 7216
rect 26160 7206 26188 7686
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 25776 7100 26084 7120
rect 25776 7098 25782 7100
rect 25838 7098 25862 7100
rect 25918 7098 25942 7100
rect 25998 7098 26022 7100
rect 26078 7098 26084 7100
rect 25838 7046 25840 7098
rect 26020 7046 26022 7098
rect 25776 7044 25782 7046
rect 25838 7044 25862 7046
rect 25918 7044 25942 7046
rect 25998 7044 26022 7046
rect 26078 7044 26084 7046
rect 25776 7024 26084 7044
rect 26148 6928 26200 6934
rect 26148 6870 26200 6876
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25700 5794 25728 6598
rect 25776 6012 26084 6032
rect 25776 6010 25782 6012
rect 25838 6010 25862 6012
rect 25918 6010 25942 6012
rect 25998 6010 26022 6012
rect 26078 6010 26084 6012
rect 25838 5958 25840 6010
rect 26020 5958 26022 6010
rect 25776 5956 25782 5958
rect 25838 5956 25862 5958
rect 25918 5956 25942 5958
rect 25998 5956 26022 5958
rect 26078 5956 26084 5958
rect 25776 5936 26084 5956
rect 25596 5772 25648 5778
rect 25700 5766 25820 5794
rect 26160 5778 26188 6870
rect 25596 5714 25648 5720
rect 25504 5704 25556 5710
rect 25504 5646 25556 5652
rect 25516 5302 25544 5646
rect 25504 5296 25556 5302
rect 25504 5238 25556 5244
rect 25516 5166 25544 5238
rect 25608 5234 25636 5714
rect 25792 5710 25820 5766
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 26620 5710 26648 8350
rect 26804 7342 26832 10610
rect 26896 10538 26924 12038
rect 26884 10532 26936 10538
rect 26884 10474 26936 10480
rect 26988 7562 27016 29702
rect 27068 29640 27120 29646
rect 27264 29594 27292 31282
rect 27356 30025 27384 31470
rect 27342 30016 27398 30025
rect 27342 29951 27398 29960
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 27068 29582 27120 29588
rect 27080 19922 27108 29582
rect 27172 29566 27292 29594
rect 27172 27033 27200 29566
rect 27252 29504 27304 29510
rect 27252 29446 27304 29452
rect 27264 29238 27292 29446
rect 27252 29232 27304 29238
rect 27252 29174 27304 29180
rect 27252 29096 27304 29102
rect 27250 29064 27252 29073
rect 27304 29064 27306 29073
rect 27250 28999 27306 29008
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27264 28150 27292 28358
rect 27252 28144 27304 28150
rect 27252 28086 27304 28092
rect 27250 27976 27306 27985
rect 27250 27911 27306 27920
rect 27264 27062 27292 27911
rect 27356 27130 27384 29786
rect 27448 27470 27476 35974
rect 27540 35737 27568 37062
rect 27632 36786 27660 37198
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 27620 36576 27672 36582
rect 27620 36518 27672 36524
rect 27526 35728 27582 35737
rect 27632 35698 27660 36518
rect 27526 35663 27582 35672
rect 27620 35692 27672 35698
rect 27620 35634 27672 35640
rect 27620 35488 27672 35494
rect 27618 35456 27620 35465
rect 27672 35456 27674 35465
rect 27618 35391 27674 35400
rect 27620 34944 27672 34950
rect 27620 34886 27672 34892
rect 27632 34746 27660 34886
rect 27620 34740 27672 34746
rect 27620 34682 27672 34688
rect 27528 34468 27580 34474
rect 27528 34410 27580 34416
rect 27540 31414 27568 34410
rect 27632 32473 27660 34682
rect 27618 32464 27674 32473
rect 27618 32399 27674 32408
rect 27724 32337 27752 40967
rect 27816 40746 27844 41919
rect 27908 41274 27936 46906
rect 28000 44577 28028 49422
rect 27986 44568 28042 44577
rect 27986 44503 28042 44512
rect 27988 44396 28040 44402
rect 27988 44338 28040 44344
rect 28000 43217 28028 44338
rect 27986 43208 28042 43217
rect 27986 43143 28042 43152
rect 27988 43104 28040 43110
rect 27988 43046 28040 43052
rect 28000 42362 28028 43046
rect 27988 42356 28040 42362
rect 27988 42298 28040 42304
rect 27988 42016 28040 42022
rect 27988 41958 28040 41964
rect 28000 41818 28028 41958
rect 27988 41812 28040 41818
rect 27988 41754 28040 41760
rect 27988 41472 28040 41478
rect 28092 41449 28120 59463
rect 28184 57798 28212 63922
rect 28264 63844 28316 63850
rect 28264 63786 28316 63792
rect 28276 63510 28304 63786
rect 28264 63504 28316 63510
rect 28264 63446 28316 63452
rect 28368 63374 28396 63922
rect 28264 63368 28316 63374
rect 28264 63310 28316 63316
rect 28356 63368 28408 63374
rect 28356 63310 28408 63316
rect 28276 57974 28304 63310
rect 28354 63064 28410 63073
rect 28354 62999 28410 63008
rect 28368 62490 28396 62999
rect 28356 62484 28408 62490
rect 28356 62426 28408 62432
rect 28356 61804 28408 61810
rect 28356 61746 28408 61752
rect 28368 60602 28396 61746
rect 28460 61305 28488 65418
rect 28552 63578 28580 74506
rect 29012 69884 29040 76910
rect 29104 70038 29132 76978
rect 29276 76084 29328 76090
rect 29276 76026 29328 76032
rect 29288 75857 29316 76026
rect 29274 75848 29330 75857
rect 29274 75783 29330 75792
rect 29184 70508 29236 70514
rect 29184 70450 29236 70456
rect 29092 70032 29144 70038
rect 29196 70009 29224 70450
rect 29092 69974 29144 69980
rect 29182 70000 29238 70009
rect 29182 69935 29238 69944
rect 29012 69856 29132 69884
rect 29000 69760 29052 69766
rect 29000 69702 29052 69708
rect 28906 68776 28962 68785
rect 28906 68711 28962 68720
rect 28920 68678 28948 68711
rect 28908 68672 28960 68678
rect 28908 68614 28960 68620
rect 29012 67946 29040 69702
rect 28828 67918 29040 67946
rect 28828 66842 28856 67918
rect 28908 67856 28960 67862
rect 28908 67798 28960 67804
rect 28920 67425 28948 67798
rect 29000 67720 29052 67726
rect 29000 67662 29052 67668
rect 28906 67416 28962 67425
rect 28906 67351 28962 67360
rect 28908 67040 28960 67046
rect 28908 66982 28960 66988
rect 28816 66836 28868 66842
rect 28816 66778 28868 66784
rect 28816 66632 28868 66638
rect 28816 66574 28868 66580
rect 28632 66156 28684 66162
rect 28632 66098 28684 66104
rect 28724 66156 28776 66162
rect 28724 66098 28776 66104
rect 28644 64569 28672 66098
rect 28630 64560 28686 64569
rect 28630 64495 28686 64504
rect 28632 64320 28684 64326
rect 28632 64262 28684 64268
rect 28540 63572 28592 63578
rect 28540 63514 28592 63520
rect 28538 63472 28594 63481
rect 28538 63407 28540 63416
rect 28592 63407 28594 63416
rect 28540 63378 28592 63384
rect 28540 63300 28592 63306
rect 28540 63242 28592 63248
rect 28552 63073 28580 63242
rect 28538 63064 28594 63073
rect 28644 63034 28672 64262
rect 28538 62999 28594 63008
rect 28632 63028 28684 63034
rect 28632 62970 28684 62976
rect 28538 62928 28594 62937
rect 28538 62863 28540 62872
rect 28592 62863 28594 62872
rect 28540 62834 28592 62840
rect 28632 62824 28684 62830
rect 28632 62766 28684 62772
rect 28540 62756 28592 62762
rect 28540 62698 28592 62704
rect 28446 61296 28502 61305
rect 28446 61231 28502 61240
rect 28448 61192 28500 61198
rect 28448 61134 28500 61140
rect 28460 60738 28488 61134
rect 28552 61033 28580 62698
rect 28644 62354 28672 62766
rect 28632 62348 28684 62354
rect 28632 62290 28684 62296
rect 28632 62212 28684 62218
rect 28632 62154 28684 62160
rect 28644 61849 28672 62154
rect 28630 61840 28686 61849
rect 28736 61810 28764 66098
rect 28828 64161 28856 66574
rect 28920 66473 28948 66982
rect 28906 66464 28962 66473
rect 28906 66399 28962 66408
rect 28908 66088 28960 66094
rect 28908 66030 28960 66036
rect 28920 65006 28948 66030
rect 28908 65000 28960 65006
rect 28908 64942 28960 64948
rect 28908 64388 28960 64394
rect 28908 64330 28960 64336
rect 28814 64152 28870 64161
rect 28814 64087 28870 64096
rect 28816 63844 28868 63850
rect 28816 63786 28868 63792
rect 28630 61775 28686 61784
rect 28724 61804 28776 61810
rect 28724 61746 28776 61752
rect 28630 61704 28686 61713
rect 28630 61639 28686 61648
rect 28724 61668 28776 61674
rect 28644 61418 28672 61639
rect 28724 61610 28776 61616
rect 28736 61577 28764 61610
rect 28828 61606 28856 63786
rect 28920 62966 28948 64330
rect 28908 62960 28960 62966
rect 28908 62902 28960 62908
rect 28816 61600 28868 61606
rect 28722 61568 28778 61577
rect 28816 61542 28868 61548
rect 28722 61503 28778 61512
rect 28828 61441 28856 61542
rect 28814 61432 28870 61441
rect 28644 61390 28764 61418
rect 28632 61260 28684 61266
rect 28632 61202 28684 61208
rect 28538 61024 28594 61033
rect 28538 60959 28594 60968
rect 28644 60858 28672 61202
rect 28632 60852 28684 60858
rect 28632 60794 28684 60800
rect 28460 60710 28672 60738
rect 28368 60574 28488 60602
rect 28356 60512 28408 60518
rect 28356 60454 28408 60460
rect 28368 60110 28396 60454
rect 28460 60330 28488 60574
rect 28538 60344 28594 60353
rect 28460 60302 28538 60330
rect 28538 60279 28594 60288
rect 28356 60104 28408 60110
rect 28356 60046 28408 60052
rect 28644 59974 28672 60710
rect 28356 59968 28408 59974
rect 28356 59910 28408 59916
rect 28632 59968 28684 59974
rect 28632 59910 28684 59916
rect 28258 57946 28304 57974
rect 28258 57916 28286 57946
rect 28368 57934 28396 59910
rect 28736 59786 28764 61390
rect 28814 61367 28870 61376
rect 28816 61328 28868 61334
rect 28814 61296 28816 61305
rect 28868 61296 28870 61305
rect 28814 61231 28870 61240
rect 28816 61192 28868 61198
rect 28814 61160 28816 61169
rect 28868 61160 28870 61169
rect 28814 61095 28870 61104
rect 28920 61044 28948 62902
rect 28828 61016 28948 61044
rect 28828 60625 28856 61016
rect 28908 60716 28960 60722
rect 28908 60658 28960 60664
rect 28814 60616 28870 60625
rect 28814 60551 28870 60560
rect 28814 60072 28870 60081
rect 28814 60007 28870 60016
rect 28552 59758 28764 59786
rect 28356 57928 28408 57934
rect 28258 57888 28304 57916
rect 28172 57792 28224 57798
rect 28172 57734 28224 57740
rect 28172 57248 28224 57254
rect 28172 57190 28224 57196
rect 28184 57089 28212 57190
rect 28170 57080 28226 57089
rect 28170 57015 28226 57024
rect 28172 56704 28224 56710
rect 28170 56672 28172 56681
rect 28224 56672 28226 56681
rect 28170 56607 28226 56616
rect 28170 56536 28226 56545
rect 28170 56471 28226 56480
rect 28184 55146 28212 56471
rect 28172 55140 28224 55146
rect 28172 55082 28224 55088
rect 28184 54534 28212 55082
rect 28172 54528 28224 54534
rect 28172 54470 28224 54476
rect 28172 53440 28224 53446
rect 28172 53382 28224 53388
rect 28184 53242 28212 53382
rect 28172 53236 28224 53242
rect 28172 53178 28224 53184
rect 28184 51105 28212 53178
rect 28170 51096 28226 51105
rect 28170 51031 28226 51040
rect 28172 50448 28224 50454
rect 28172 50390 28224 50396
rect 28184 49298 28212 50390
rect 28172 49292 28224 49298
rect 28172 49234 28224 49240
rect 28172 49156 28224 49162
rect 28172 49098 28224 49104
rect 28184 41721 28212 49098
rect 28276 49042 28304 57888
rect 28356 57870 28408 57876
rect 28354 56808 28410 56817
rect 28354 56743 28410 56752
rect 28368 49162 28396 56743
rect 28448 55752 28500 55758
rect 28448 55694 28500 55700
rect 28460 55350 28488 55694
rect 28448 55344 28500 55350
rect 28448 55286 28500 55292
rect 28460 53174 28488 55286
rect 28448 53168 28500 53174
rect 28448 53110 28500 53116
rect 28460 52494 28488 53110
rect 28448 52488 28500 52494
rect 28448 52430 28500 52436
rect 28460 52086 28488 52430
rect 28448 52080 28500 52086
rect 28448 52022 28500 52028
rect 28446 51912 28502 51921
rect 28446 51847 28502 51856
rect 28356 49156 28408 49162
rect 28356 49098 28408 49104
rect 28276 49014 28396 49042
rect 28262 48920 28318 48929
rect 28262 48855 28264 48864
rect 28316 48855 28318 48864
rect 28264 48826 28316 48832
rect 28262 48784 28318 48793
rect 28262 48719 28264 48728
rect 28316 48719 28318 48728
rect 28264 48690 28316 48696
rect 28264 48544 28316 48550
rect 28264 48486 28316 48492
rect 28276 44878 28304 48486
rect 28368 48278 28396 49014
rect 28356 48272 28408 48278
rect 28356 48214 28408 48220
rect 28356 47456 28408 47462
rect 28356 47398 28408 47404
rect 28368 46918 28396 47398
rect 28356 46912 28408 46918
rect 28356 46854 28408 46860
rect 28356 45892 28408 45898
rect 28356 45834 28408 45840
rect 28368 45490 28396 45834
rect 28356 45484 28408 45490
rect 28356 45426 28408 45432
rect 28356 44940 28408 44946
rect 28356 44882 28408 44888
rect 28264 44872 28316 44878
rect 28264 44814 28316 44820
rect 28368 44470 28396 44882
rect 28356 44464 28408 44470
rect 28356 44406 28408 44412
rect 28264 44396 28316 44402
rect 28264 44338 28316 44344
rect 28276 43858 28304 44338
rect 28264 43852 28316 43858
rect 28264 43794 28316 43800
rect 28356 43784 28408 43790
rect 28356 43726 28408 43732
rect 28264 43716 28316 43722
rect 28264 43658 28316 43664
rect 28276 42906 28304 43658
rect 28264 42900 28316 42906
rect 28264 42842 28316 42848
rect 28264 42696 28316 42702
rect 28264 42638 28316 42644
rect 28276 42226 28304 42638
rect 28368 42634 28396 43726
rect 28356 42628 28408 42634
rect 28356 42570 28408 42576
rect 28368 42294 28396 42570
rect 28356 42288 28408 42294
rect 28356 42230 28408 42236
rect 28264 42220 28316 42226
rect 28264 42162 28316 42168
rect 28170 41712 28226 41721
rect 28170 41647 28226 41656
rect 28172 41608 28224 41614
rect 28276 41596 28304 42162
rect 28356 42084 28408 42090
rect 28356 42026 28408 42032
rect 28224 41568 28304 41596
rect 28172 41550 28224 41556
rect 27988 41414 28040 41420
rect 28078 41440 28134 41449
rect 27896 41268 27948 41274
rect 27896 41210 27948 41216
rect 28000 41041 28028 41414
rect 28078 41375 28134 41384
rect 28080 41268 28132 41274
rect 28080 41210 28132 41216
rect 28092 41052 28120 41210
rect 28184 41206 28212 41550
rect 28262 41440 28318 41449
rect 28262 41375 28318 41384
rect 28276 41206 28304 41375
rect 28172 41200 28224 41206
rect 28172 41142 28224 41148
rect 28264 41200 28316 41206
rect 28264 41142 28316 41148
rect 27986 41032 28042 41041
rect 28092 41024 28304 41052
rect 27986 40967 28042 40976
rect 28172 40928 28224 40934
rect 27986 40896 28042 40905
rect 28042 40854 28120 40882
rect 28172 40870 28224 40876
rect 27986 40831 28042 40840
rect 27816 40718 27936 40746
rect 27804 40656 27856 40662
rect 27804 40598 27856 40604
rect 27816 40225 27844 40598
rect 27802 40216 27858 40225
rect 27802 40151 27858 40160
rect 27802 40080 27858 40089
rect 27802 40015 27858 40024
rect 27710 32328 27766 32337
rect 27710 32263 27766 32272
rect 27712 32224 27764 32230
rect 27712 32166 27764 32172
rect 27724 32065 27752 32166
rect 27710 32056 27766 32065
rect 27710 31991 27766 32000
rect 27712 31884 27764 31890
rect 27712 31826 27764 31832
rect 27618 31784 27674 31793
rect 27618 31719 27674 31728
rect 27528 31408 27580 31414
rect 27528 31350 27580 31356
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27540 30977 27568 31214
rect 27526 30968 27582 30977
rect 27526 30903 27582 30912
rect 27526 30832 27582 30841
rect 27526 30767 27582 30776
rect 27540 29345 27568 30767
rect 27632 30326 27660 31719
rect 27724 31482 27752 31826
rect 27712 31476 27764 31482
rect 27712 31418 27764 31424
rect 27816 30682 27844 40015
rect 27724 30654 27844 30682
rect 27724 30394 27752 30654
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27620 30320 27672 30326
rect 27620 30262 27672 30268
rect 27724 29578 27752 30330
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27816 29850 27844 30194
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27908 29730 27936 40718
rect 28092 39896 28120 40854
rect 28184 40118 28212 40870
rect 28172 40112 28224 40118
rect 28172 40054 28224 40060
rect 28172 39976 28224 39982
rect 28000 39868 28120 39896
rect 28170 39944 28172 39953
rect 28224 39944 28226 39953
rect 28170 39879 28226 39888
rect 28000 39438 28028 39868
rect 28276 39828 28304 41024
rect 28368 40594 28396 42026
rect 28356 40588 28408 40594
rect 28356 40530 28408 40536
rect 28356 40452 28408 40458
rect 28356 40394 28408 40400
rect 28368 40050 28396 40394
rect 28356 40044 28408 40050
rect 28356 39986 28408 39992
rect 28092 39800 28304 39828
rect 27988 39432 28040 39438
rect 27988 39374 28040 39380
rect 27986 38448 28042 38457
rect 27986 38383 28042 38392
rect 28000 37369 28028 38383
rect 27986 37360 28042 37369
rect 27986 37295 28042 37304
rect 27988 37256 28040 37262
rect 27988 37198 28040 37204
rect 28000 36786 28028 37198
rect 27988 36780 28040 36786
rect 27988 36722 28040 36728
rect 27988 35828 28040 35834
rect 27988 35770 28040 35776
rect 28000 33998 28028 35770
rect 27988 33992 28040 33998
rect 27988 33934 28040 33940
rect 27988 33516 28040 33522
rect 27988 33458 28040 33464
rect 28000 32774 28028 33458
rect 27988 32768 28040 32774
rect 28092 32745 28120 39800
rect 28264 39636 28316 39642
rect 28264 39578 28316 39584
rect 28172 39296 28224 39302
rect 28170 39264 28172 39273
rect 28224 39264 28226 39273
rect 28170 39199 28226 39208
rect 28172 38480 28224 38486
rect 28172 38422 28224 38428
rect 28184 38321 28212 38422
rect 28170 38312 28226 38321
rect 28170 38247 28226 38256
rect 28276 38214 28304 39578
rect 28356 39092 28408 39098
rect 28356 39034 28408 39040
rect 28264 38208 28316 38214
rect 28264 38150 28316 38156
rect 28172 37936 28224 37942
rect 28172 37878 28224 37884
rect 28184 37194 28212 37878
rect 28276 37874 28304 38150
rect 28264 37868 28316 37874
rect 28264 37810 28316 37816
rect 28368 37670 28396 39034
rect 28356 37664 28408 37670
rect 28356 37606 28408 37612
rect 28262 37224 28318 37233
rect 28172 37188 28224 37194
rect 28262 37159 28318 37168
rect 28172 37130 28224 37136
rect 28184 36360 28212 37130
rect 28276 37126 28304 37159
rect 28264 37120 28316 37126
rect 28264 37062 28316 37068
rect 28262 36952 28318 36961
rect 28262 36887 28264 36896
rect 28316 36887 28318 36896
rect 28264 36858 28316 36864
rect 28356 36712 28408 36718
rect 28356 36654 28408 36660
rect 28184 36332 28304 36360
rect 28172 36236 28224 36242
rect 28172 36178 28224 36184
rect 28184 35086 28212 36178
rect 28276 36106 28304 36332
rect 28368 36174 28396 36654
rect 28356 36168 28408 36174
rect 28356 36110 28408 36116
rect 28264 36100 28316 36106
rect 28264 36042 28316 36048
rect 28356 36032 28408 36038
rect 28356 35974 28408 35980
rect 28262 35728 28318 35737
rect 28262 35663 28264 35672
rect 28316 35663 28318 35672
rect 28264 35634 28316 35640
rect 28172 35080 28224 35086
rect 28172 35022 28224 35028
rect 28264 35012 28316 35018
rect 28264 34954 28316 34960
rect 28170 34912 28226 34921
rect 28170 34847 28226 34856
rect 28184 34202 28212 34847
rect 28172 34196 28224 34202
rect 28172 34138 28224 34144
rect 28276 33538 28304 34954
rect 28184 33510 28304 33538
rect 27988 32710 28040 32716
rect 28078 32736 28134 32745
rect 28078 32671 28134 32680
rect 28078 32600 28134 32609
rect 28078 32535 28134 32544
rect 28092 32434 28120 32535
rect 28080 32428 28132 32434
rect 28080 32370 28132 32376
rect 28078 32328 28134 32337
rect 28184 32298 28212 33510
rect 28264 33448 28316 33454
rect 28264 33390 28316 33396
rect 28276 32484 28304 33390
rect 28368 32552 28396 35974
rect 28460 32774 28488 51847
rect 28552 50250 28580 59758
rect 28724 59560 28776 59566
rect 28724 59502 28776 59508
rect 28630 59256 28686 59265
rect 28630 59191 28632 59200
rect 28684 59191 28686 59200
rect 28632 59162 28684 59168
rect 28630 58984 28686 58993
rect 28630 58919 28632 58928
rect 28684 58919 28686 58928
rect 28632 58890 28684 58896
rect 28630 58712 28686 58721
rect 28630 58647 28632 58656
rect 28684 58647 28686 58656
rect 28632 58618 28684 58624
rect 28632 58540 28684 58546
rect 28632 58482 28684 58488
rect 28644 56137 28672 58482
rect 28736 57225 28764 59502
rect 28722 57216 28778 57225
rect 28722 57151 28778 57160
rect 28722 56944 28778 56953
rect 28722 56879 28778 56888
rect 28736 56846 28764 56879
rect 28724 56840 28776 56846
rect 28724 56782 28776 56788
rect 28724 56364 28776 56370
rect 28724 56306 28776 56312
rect 28630 56128 28686 56137
rect 28630 56063 28686 56072
rect 28632 55616 28684 55622
rect 28632 55558 28684 55564
rect 28644 55282 28672 55558
rect 28736 55457 28764 56306
rect 28828 55593 28856 60007
rect 28920 59401 28948 60658
rect 28906 59392 28962 59401
rect 28906 59327 28962 59336
rect 28906 58848 28962 58857
rect 28906 58783 28962 58792
rect 28920 55826 28948 58783
rect 28908 55820 28960 55826
rect 28908 55762 28960 55768
rect 28814 55584 28870 55593
rect 28814 55519 28870 55528
rect 28722 55448 28778 55457
rect 28722 55383 28778 55392
rect 28814 55312 28870 55321
rect 28632 55276 28684 55282
rect 28814 55247 28816 55256
rect 28632 55218 28684 55224
rect 28868 55247 28870 55256
rect 28816 55218 28868 55224
rect 28814 55176 28870 55185
rect 28814 55111 28870 55120
rect 28632 55072 28684 55078
rect 28632 55014 28684 55020
rect 28644 54874 28672 55014
rect 28632 54868 28684 54874
rect 28632 54810 28684 54816
rect 28632 54596 28684 54602
rect 28632 54538 28684 54544
rect 28644 54233 28672 54538
rect 28630 54224 28686 54233
rect 28630 54159 28686 54168
rect 28724 53576 28776 53582
rect 28724 53518 28776 53524
rect 28632 53100 28684 53106
rect 28632 53042 28684 53048
rect 28644 52902 28672 53042
rect 28632 52896 28684 52902
rect 28632 52838 28684 52844
rect 28630 52728 28686 52737
rect 28630 52663 28686 52672
rect 28644 52630 28672 52663
rect 28632 52624 28684 52630
rect 28632 52566 28684 52572
rect 28632 52488 28684 52494
rect 28632 52430 28684 52436
rect 28644 52193 28672 52430
rect 28736 52329 28764 53518
rect 28722 52320 28778 52329
rect 28722 52255 28778 52264
rect 28630 52184 28686 52193
rect 28630 52119 28686 52128
rect 28724 52148 28776 52154
rect 28644 51377 28672 52119
rect 28724 52090 28776 52096
rect 28736 52057 28764 52090
rect 28722 52048 28778 52057
rect 28722 51983 28778 51992
rect 28722 51912 28778 51921
rect 28722 51847 28778 51856
rect 28736 51406 28764 51847
rect 28724 51400 28776 51406
rect 28630 51368 28686 51377
rect 28724 51342 28776 51348
rect 28630 51303 28686 51312
rect 28828 51252 28856 55111
rect 29012 53224 29040 67662
rect 29104 67114 29132 69856
rect 29472 69714 29500 77266
rect 30012 76832 30064 76838
rect 30116 76809 30144 77318
rect 30012 76774 30064 76780
rect 30102 76800 30158 76809
rect 29736 76424 29788 76430
rect 30024 76401 30052 76774
rect 30102 76735 30158 76744
rect 29736 76366 29788 76372
rect 30010 76392 30066 76401
rect 29644 72684 29696 72690
rect 29644 72626 29696 72632
rect 29380 69686 29500 69714
rect 29184 69556 29236 69562
rect 29184 69498 29236 69504
rect 29092 67108 29144 67114
rect 29092 67050 29144 67056
rect 29092 66836 29144 66842
rect 29092 66778 29144 66784
rect 29104 64326 29132 66778
rect 29092 64320 29144 64326
rect 29092 64262 29144 64268
rect 29092 64048 29144 64054
rect 29092 63990 29144 63996
rect 29104 63374 29132 63990
rect 29092 63368 29144 63374
rect 29092 63310 29144 63316
rect 29196 63034 29224 69498
rect 29380 69476 29408 69686
rect 29552 69488 29604 69494
rect 29380 69448 29500 69476
rect 29368 69352 29420 69358
rect 29274 69320 29330 69329
rect 29368 69294 29420 69300
rect 29274 69255 29276 69264
rect 29328 69255 29330 69264
rect 29276 69226 29328 69232
rect 29276 68808 29328 68814
rect 29276 68750 29328 68756
rect 29288 63306 29316 68750
rect 29276 63300 29328 63306
rect 29276 63242 29328 63248
rect 29184 63028 29236 63034
rect 29380 63016 29408 69294
rect 29472 68474 29500 69448
rect 29552 69430 29604 69436
rect 29460 68468 29512 68474
rect 29460 68410 29512 68416
rect 29460 67720 29512 67726
rect 29460 67662 29512 67668
rect 29472 66298 29500 67662
rect 29460 66292 29512 66298
rect 29460 66234 29512 66240
rect 29564 66178 29592 69430
rect 29472 66150 29592 66178
rect 29472 64122 29500 66150
rect 29552 66020 29604 66026
rect 29552 65962 29604 65968
rect 29460 64116 29512 64122
rect 29460 64058 29512 64064
rect 29460 63980 29512 63986
rect 29460 63922 29512 63928
rect 29184 62970 29236 62976
rect 29288 62988 29408 63016
rect 29184 62824 29236 62830
rect 29184 62766 29236 62772
rect 29092 62280 29144 62286
rect 29092 62222 29144 62228
rect 29104 61334 29132 62222
rect 29196 61810 29224 62766
rect 29288 62354 29316 62988
rect 29368 62892 29420 62898
rect 29368 62834 29420 62840
rect 29276 62348 29328 62354
rect 29276 62290 29328 62296
rect 29184 61804 29236 61810
rect 29184 61746 29236 61752
rect 29092 61328 29144 61334
rect 29092 61270 29144 61276
rect 29092 61192 29144 61198
rect 29090 61160 29092 61169
rect 29144 61160 29146 61169
rect 29090 61095 29146 61104
rect 29092 61056 29144 61062
rect 29092 60998 29144 61004
rect 29104 60722 29132 60998
rect 29196 60874 29224 61746
rect 29380 61418 29408 62834
rect 29472 62490 29500 63922
rect 29564 63238 29592 65962
rect 29552 63232 29604 63238
rect 29552 63174 29604 63180
rect 29460 62484 29512 62490
rect 29460 62426 29512 62432
rect 29460 62348 29512 62354
rect 29460 62290 29512 62296
rect 29288 61390 29408 61418
rect 29288 61334 29316 61390
rect 29276 61328 29328 61334
rect 29276 61270 29328 61276
rect 29368 61328 29420 61334
rect 29368 61270 29420 61276
rect 29274 60888 29330 60897
rect 29196 60846 29274 60874
rect 29274 60823 29330 60832
rect 29182 60752 29238 60761
rect 29092 60716 29144 60722
rect 29380 60734 29408 61270
rect 29472 60874 29500 62290
rect 29564 61010 29592 63174
rect 29656 61169 29684 72626
rect 29748 69494 29776 76366
rect 30010 76327 30066 76336
rect 30196 76288 30248 76294
rect 30196 76230 30248 76236
rect 30104 76016 30156 76022
rect 30104 75958 30156 75964
rect 29828 75948 29880 75954
rect 29828 75890 29880 75896
rect 29840 69562 29868 75890
rect 30012 75744 30064 75750
rect 30012 75686 30064 75692
rect 29920 75336 29972 75342
rect 29920 75278 29972 75284
rect 29828 69556 29880 69562
rect 29828 69498 29880 69504
rect 29736 69488 29788 69494
rect 29736 69430 29788 69436
rect 29932 69306 29960 75278
rect 30024 74905 30052 75686
rect 30010 74896 30066 74905
rect 30010 74831 30066 74840
rect 30012 74656 30064 74662
rect 30012 74598 30064 74604
rect 30024 74089 30052 74598
rect 30010 74080 30066 74089
rect 30010 74015 30066 74024
rect 30012 73568 30064 73574
rect 30012 73510 30064 73516
rect 30024 73137 30052 73510
rect 30010 73128 30066 73137
rect 30010 73063 30066 73072
rect 30012 73024 30064 73030
rect 30012 72966 30064 72972
rect 30024 72593 30052 72966
rect 30010 72584 30066 72593
rect 30010 72519 30066 72528
rect 30012 72480 30064 72486
rect 30012 72422 30064 72428
rect 30024 72185 30052 72422
rect 30010 72176 30066 72185
rect 30010 72111 30066 72120
rect 30012 71936 30064 71942
rect 30012 71878 30064 71884
rect 30024 71641 30052 71878
rect 30010 71632 30066 71641
rect 30010 71567 30066 71576
rect 30012 71392 30064 71398
rect 30012 71334 30064 71340
rect 30024 71233 30052 71334
rect 30010 71224 30066 71233
rect 30010 71159 30066 71168
rect 30012 70848 30064 70854
rect 30012 70790 30064 70796
rect 30024 70689 30052 70790
rect 30010 70680 30066 70689
rect 30010 70615 30066 70624
rect 30012 70304 30064 70310
rect 30010 70272 30012 70281
rect 30064 70272 30066 70281
rect 30010 70207 30066 70216
rect 30012 69760 30064 69766
rect 30010 69728 30012 69737
rect 30064 69728 30066 69737
rect 30010 69663 30066 69672
rect 29748 69278 29960 69306
rect 29748 63458 29776 69278
rect 29920 69216 29972 69222
rect 29920 69158 29972 69164
rect 29932 68377 29960 69158
rect 30012 68672 30064 68678
rect 30012 68614 30064 68620
rect 29918 68368 29974 68377
rect 29918 68303 29974 68312
rect 29920 68128 29972 68134
rect 29920 68070 29972 68076
rect 29828 67040 29880 67046
rect 29932 67017 29960 68070
rect 30024 67969 30052 68614
rect 30010 67960 30066 67969
rect 30010 67895 30066 67904
rect 30012 67856 30064 67862
rect 30012 67798 30064 67804
rect 29828 66982 29880 66988
rect 29918 67008 29974 67017
rect 29840 65113 29868 66982
rect 29918 66943 29974 66952
rect 30024 66065 30052 67798
rect 30116 66230 30144 75958
rect 30208 75449 30236 76230
rect 30194 75440 30250 75449
rect 30194 75375 30250 75384
rect 30196 75200 30248 75206
rect 30196 75142 30248 75148
rect 30208 74497 30236 75142
rect 30194 74488 30250 74497
rect 30194 74423 30250 74432
rect 30196 74112 30248 74118
rect 30196 74054 30248 74060
rect 30208 73545 30236 74054
rect 30194 73536 30250 73545
rect 30194 73471 30250 73480
rect 30196 72072 30248 72078
rect 30196 72014 30248 72020
rect 30104 66224 30156 66230
rect 30104 66166 30156 66172
rect 30104 66088 30156 66094
rect 30010 66056 30066 66065
rect 30104 66030 30156 66036
rect 30010 65991 30066 66000
rect 29920 65952 29972 65958
rect 29920 65894 29972 65900
rect 29932 65686 29960 65894
rect 29920 65680 29972 65686
rect 29920 65622 29972 65628
rect 29920 65544 29972 65550
rect 29920 65486 29972 65492
rect 29826 65104 29882 65113
rect 29826 65039 29882 65048
rect 29828 65000 29880 65006
rect 29828 64942 29880 64948
rect 29840 64394 29868 64942
rect 29828 64388 29880 64394
rect 29828 64330 29880 64336
rect 29932 63617 29960 65486
rect 30012 65068 30064 65074
rect 30012 65010 30064 65016
rect 30024 63986 30052 65010
rect 30012 63980 30064 63986
rect 30012 63922 30064 63928
rect 29918 63608 29974 63617
rect 29918 63543 29974 63552
rect 29748 63430 29960 63458
rect 29828 63368 29880 63374
rect 29828 63310 29880 63316
rect 29736 63300 29788 63306
rect 29736 63242 29788 63248
rect 29748 61402 29776 63242
rect 29736 61396 29788 61402
rect 29736 61338 29788 61344
rect 29734 61296 29790 61305
rect 29734 61231 29790 61240
rect 29642 61160 29698 61169
rect 29642 61095 29698 61104
rect 29564 60982 29684 61010
rect 29472 60846 29592 60874
rect 29182 60687 29238 60696
rect 29288 60706 29408 60734
rect 29460 60784 29512 60790
rect 29460 60726 29512 60732
rect 29092 60658 29144 60664
rect 29090 60616 29146 60625
rect 29090 60551 29146 60560
rect 29104 58614 29132 60551
rect 29092 58608 29144 58614
rect 29092 58550 29144 58556
rect 29104 57934 29132 58550
rect 29092 57928 29144 57934
rect 29092 57870 29144 57876
rect 29196 57798 29224 60687
rect 29092 57792 29144 57798
rect 29092 57734 29144 57740
rect 29184 57792 29236 57798
rect 29184 57734 29236 57740
rect 29104 57050 29132 57734
rect 29196 57390 29224 57734
rect 29184 57384 29236 57390
rect 29184 57326 29236 57332
rect 29092 57044 29144 57050
rect 29092 56986 29144 56992
rect 29092 56908 29144 56914
rect 29092 56850 29144 56856
rect 29104 56438 29132 56850
rect 29196 56506 29224 57326
rect 29184 56500 29236 56506
rect 29184 56442 29236 56448
rect 29092 56432 29144 56438
rect 29144 56380 29224 56386
rect 29092 56374 29224 56380
rect 29104 56358 29224 56374
rect 29092 56296 29144 56302
rect 29092 56238 29144 56244
rect 29104 54058 29132 56238
rect 29196 55593 29224 56358
rect 29182 55584 29238 55593
rect 29182 55519 29238 55528
rect 29184 55412 29236 55418
rect 29184 55354 29236 55360
rect 29092 54052 29144 54058
rect 29092 53994 29144 54000
rect 29196 53553 29224 55354
rect 29182 53544 29238 53553
rect 29182 53479 29238 53488
rect 29092 53440 29144 53446
rect 29090 53408 29092 53417
rect 29144 53408 29146 53417
rect 29090 53343 29146 53352
rect 29288 53242 29316 60706
rect 29472 60654 29500 60726
rect 29368 60648 29420 60654
rect 29368 60590 29420 60596
rect 29460 60648 29512 60654
rect 29460 60590 29512 60596
rect 29380 60489 29408 60590
rect 29366 60480 29422 60489
rect 29366 60415 29422 60424
rect 29366 60208 29422 60217
rect 29366 60143 29422 60152
rect 29380 59022 29408 60143
rect 29460 59968 29512 59974
rect 29460 59910 29512 59916
rect 29368 59016 29420 59022
rect 29368 58958 29420 58964
rect 29368 58540 29420 58546
rect 29368 58482 29420 58488
rect 29380 58138 29408 58482
rect 29368 58132 29420 58138
rect 29368 58074 29420 58080
rect 29368 57928 29420 57934
rect 29368 57870 29420 57876
rect 29380 56681 29408 57870
rect 29366 56672 29422 56681
rect 29366 56607 29422 56616
rect 29380 55622 29408 56607
rect 29368 55616 29420 55622
rect 29368 55558 29420 55564
rect 29380 54330 29408 55558
rect 29472 54330 29500 59910
rect 29368 54324 29420 54330
rect 29368 54266 29420 54272
rect 29460 54324 29512 54330
rect 29460 54266 29512 54272
rect 29368 54188 29420 54194
rect 29368 54130 29420 54136
rect 28966 53196 29040 53224
rect 29276 53236 29328 53242
rect 28966 53088 28994 53196
rect 29276 53178 29328 53184
rect 29274 53136 29330 53145
rect 29196 53094 29274 53122
rect 28966 53060 29132 53088
rect 28906 53000 28962 53009
rect 28906 52935 28962 52944
rect 28920 52562 28948 52935
rect 28908 52556 28960 52562
rect 29000 52556 29052 52562
rect 28960 52516 29000 52544
rect 28908 52498 28960 52504
rect 29000 52498 29052 52504
rect 29000 52352 29052 52358
rect 29104 52340 29132 53060
rect 29196 52698 29224 53094
rect 29274 53071 29330 53080
rect 29276 52964 29328 52970
rect 29276 52906 29328 52912
rect 29288 52737 29316 52906
rect 29274 52728 29330 52737
rect 29184 52692 29236 52698
rect 29274 52663 29330 52672
rect 29184 52634 29236 52640
rect 29380 52601 29408 54130
rect 29458 54088 29514 54097
rect 29458 54023 29514 54032
rect 29472 52698 29500 54023
rect 29460 52692 29512 52698
rect 29460 52634 29512 52640
rect 29366 52592 29422 52601
rect 29276 52556 29328 52562
rect 29366 52527 29422 52536
rect 29276 52498 29328 52504
rect 29052 52312 29132 52340
rect 29000 52294 29052 52300
rect 29182 52184 29238 52193
rect 29012 52142 29182 52170
rect 28908 51944 28960 51950
rect 28908 51886 28960 51892
rect 28920 51270 28948 51886
rect 28644 51224 28856 51252
rect 28908 51264 28960 51270
rect 28906 51232 28908 51241
rect 28960 51232 28962 51241
rect 28540 50244 28592 50250
rect 28540 50186 28592 50192
rect 28540 49904 28592 49910
rect 28540 49846 28592 49852
rect 28552 45529 28580 49846
rect 28538 45520 28594 45529
rect 28538 45455 28594 45464
rect 28540 45416 28592 45422
rect 28540 45358 28592 45364
rect 28552 44402 28580 45358
rect 28540 44396 28592 44402
rect 28540 44338 28592 44344
rect 28644 44316 28672 51224
rect 28906 51167 28962 51176
rect 29012 51074 29040 52142
rect 29182 52119 29238 52128
rect 29090 52048 29146 52057
rect 29288 52034 29316 52498
rect 29458 52456 29514 52465
rect 29458 52391 29514 52400
rect 29368 52148 29420 52154
rect 29368 52090 29420 52096
rect 29196 52018 29316 52034
rect 29090 51983 29146 51992
rect 29184 52012 29316 52018
rect 29104 51814 29132 51983
rect 29236 52006 29316 52012
rect 29184 51954 29236 51960
rect 29276 51944 29328 51950
rect 29276 51886 29328 51892
rect 29092 51808 29144 51814
rect 29092 51750 29144 51756
rect 29092 51264 29144 51270
rect 29092 51206 29144 51212
rect 29182 51232 29238 51241
rect 29104 51105 29132 51206
rect 29182 51167 29238 51176
rect 28920 51046 29040 51074
rect 29090 51096 29146 51105
rect 28816 50924 28868 50930
rect 28816 50866 28868 50872
rect 28724 50244 28776 50250
rect 28724 50186 28776 50192
rect 28736 49881 28764 50186
rect 28722 49872 28778 49881
rect 28722 49807 28778 49816
rect 28724 49224 28776 49230
rect 28724 49166 28776 49172
rect 28736 48249 28764 49166
rect 28828 49065 28856 50866
rect 28814 49056 28870 49065
rect 28814 48991 28870 49000
rect 28814 48648 28870 48657
rect 28814 48583 28870 48592
rect 28722 48240 28778 48249
rect 28722 48175 28778 48184
rect 28722 48104 28778 48113
rect 28722 48039 28778 48048
rect 28736 47054 28764 48039
rect 28724 47048 28776 47054
rect 28724 46990 28776 46996
rect 28724 46708 28776 46714
rect 28724 46650 28776 46656
rect 28736 45082 28764 46650
rect 28828 46578 28856 48583
rect 28920 46714 28948 51046
rect 29090 51031 29146 51040
rect 29000 50856 29052 50862
rect 29000 50798 29052 50804
rect 29012 50425 29040 50798
rect 29092 50720 29144 50726
rect 29092 50662 29144 50668
rect 28998 50416 29054 50425
rect 28998 50351 29054 50360
rect 29000 50244 29052 50250
rect 29000 50186 29052 50192
rect 29012 49842 29040 50186
rect 29104 49910 29132 50662
rect 29092 49904 29144 49910
rect 29092 49846 29144 49852
rect 29000 49836 29052 49842
rect 29000 49778 29052 49784
rect 29000 48884 29052 48890
rect 29000 48826 29052 48832
rect 29012 48142 29040 48826
rect 29092 48748 29144 48754
rect 29092 48690 29144 48696
rect 29000 48136 29052 48142
rect 29000 48078 29052 48084
rect 29000 48000 29052 48006
rect 28998 47968 29000 47977
rect 29052 47968 29054 47977
rect 28998 47903 29054 47912
rect 29000 47728 29052 47734
rect 29000 47670 29052 47676
rect 28908 46708 28960 46714
rect 28908 46650 28960 46656
rect 28816 46572 28868 46578
rect 28816 46514 28868 46520
rect 28906 45928 28962 45937
rect 28906 45863 28962 45872
rect 28920 45626 28948 45863
rect 28908 45620 28960 45626
rect 28908 45562 28960 45568
rect 28908 45280 28960 45286
rect 28908 45222 28960 45228
rect 28724 45076 28776 45082
rect 28724 45018 28776 45024
rect 28920 44946 28948 45222
rect 28908 44940 28960 44946
rect 28908 44882 28960 44888
rect 28724 44872 28776 44878
rect 28724 44814 28776 44820
rect 28814 44840 28870 44849
rect 28736 44441 28764 44814
rect 28814 44775 28870 44784
rect 28722 44432 28778 44441
rect 28828 44402 28856 44775
rect 28908 44736 28960 44742
rect 28908 44678 28960 44684
rect 28722 44367 28778 44376
rect 28816 44396 28868 44402
rect 28816 44338 28868 44344
rect 28644 44288 28764 44316
rect 28920 44305 28948 44678
rect 28632 42900 28684 42906
rect 28632 42842 28684 42848
rect 28540 42220 28592 42226
rect 28540 42162 28592 42168
rect 28552 41614 28580 42162
rect 28644 42072 28672 42842
rect 28625 42044 28672 42072
rect 28625 41936 28653 42044
rect 28625 41908 28672 41936
rect 28540 41608 28592 41614
rect 28540 41550 28592 41556
rect 28552 41449 28580 41550
rect 28538 41440 28594 41449
rect 28538 41375 28594 41384
rect 28552 41177 28580 41375
rect 28538 41168 28594 41177
rect 28644 41154 28672 41908
rect 28736 41592 28764 44288
rect 28906 44296 28962 44305
rect 28906 44231 28962 44240
rect 28906 44160 28962 44169
rect 28906 44095 28962 44104
rect 28920 43194 28948 44095
rect 29012 43353 29040 47670
rect 29104 46374 29132 48690
rect 29092 46368 29144 46374
rect 29092 46310 29144 46316
rect 29104 45665 29132 46310
rect 29196 45966 29224 51167
rect 29184 45960 29236 45966
rect 29184 45902 29236 45908
rect 29184 45824 29236 45830
rect 29184 45766 29236 45772
rect 29090 45656 29146 45665
rect 29090 45591 29146 45600
rect 29090 45520 29146 45529
rect 29090 45455 29146 45464
rect 29104 45286 29132 45455
rect 29092 45280 29144 45286
rect 29092 45222 29144 45228
rect 29092 45008 29144 45014
rect 29092 44950 29144 44956
rect 28998 43344 29054 43353
rect 29104 43314 29132 44950
rect 28998 43279 29054 43288
rect 29092 43308 29144 43314
rect 29092 43250 29144 43256
rect 28920 43166 29132 43194
rect 29104 42786 29132 43166
rect 28908 42764 28960 42770
rect 28908 42706 28960 42712
rect 29012 42758 29132 42786
rect 28816 42560 28868 42566
rect 28816 42502 28868 42508
rect 28828 41818 28856 42502
rect 28920 42378 28948 42706
rect 29012 42566 29040 42758
rect 29000 42560 29052 42566
rect 29000 42502 29052 42508
rect 28920 42350 29132 42378
rect 28908 42288 28960 42294
rect 28908 42230 28960 42236
rect 28920 41970 28948 42230
rect 29104 42090 29132 42350
rect 29196 42265 29224 45766
rect 29288 45354 29316 51886
rect 29380 51474 29408 52090
rect 29472 51814 29500 52391
rect 29564 52358 29592 60846
rect 29656 53990 29684 60982
rect 29748 60790 29776 61231
rect 29840 60897 29868 63310
rect 29826 60888 29882 60897
rect 29826 60823 29882 60832
rect 29736 60784 29788 60790
rect 29736 60726 29788 60732
rect 29932 60734 29960 63430
rect 30024 62898 30052 63922
rect 30012 62892 30064 62898
rect 30012 62834 30064 62840
rect 30012 62280 30064 62286
rect 30012 62222 30064 62228
rect 30024 61198 30052 62222
rect 30012 61192 30064 61198
rect 30012 61134 30064 61140
rect 30024 61033 30052 61134
rect 30116 61062 30144 66030
rect 30104 61056 30156 61062
rect 30010 61024 30066 61033
rect 30104 60998 30156 61004
rect 30010 60959 30066 60968
rect 29932 60706 30052 60734
rect 29736 60512 29788 60518
rect 29736 60454 29788 60460
rect 29828 60512 29880 60518
rect 29828 60454 29880 60460
rect 29748 59226 29776 60454
rect 29840 59809 29868 60454
rect 29920 60104 29972 60110
rect 29920 60046 29972 60052
rect 29826 59800 29882 59809
rect 29826 59735 29882 59744
rect 29828 59628 29880 59634
rect 29828 59570 29880 59576
rect 29736 59220 29788 59226
rect 29736 59162 29788 59168
rect 29736 58948 29788 58954
rect 29736 58890 29788 58896
rect 29748 58041 29776 58890
rect 29840 58449 29868 59570
rect 29826 58440 29882 58449
rect 29826 58375 29882 58384
rect 29828 58336 29880 58342
rect 29828 58278 29880 58284
rect 29734 58032 29790 58041
rect 29734 57967 29790 57976
rect 29734 57896 29790 57905
rect 29734 57831 29790 57840
rect 29748 57594 29776 57831
rect 29736 57588 29788 57594
rect 29736 57530 29788 57536
rect 29734 57488 29790 57497
rect 29734 57423 29736 57432
rect 29788 57423 29790 57432
rect 29736 57394 29788 57400
rect 29736 57316 29788 57322
rect 29736 57258 29788 57264
rect 29748 57225 29776 57258
rect 29734 57216 29790 57225
rect 29734 57151 29790 57160
rect 29736 56840 29788 56846
rect 29736 56782 29788 56788
rect 29748 56506 29776 56782
rect 29736 56500 29788 56506
rect 29736 56442 29788 56448
rect 29736 55684 29788 55690
rect 29736 55626 29788 55632
rect 29748 55185 29776 55626
rect 29734 55176 29790 55185
rect 29734 55111 29790 55120
rect 29734 54768 29790 54777
rect 29734 54703 29790 54712
rect 29748 54670 29776 54703
rect 29736 54664 29788 54670
rect 29736 54606 29788 54612
rect 29644 53984 29696 53990
rect 29644 53926 29696 53932
rect 29734 53816 29790 53825
rect 29644 53780 29696 53786
rect 29734 53751 29790 53760
rect 29644 53722 29696 53728
rect 29656 53689 29684 53722
rect 29642 53680 29698 53689
rect 29642 53615 29698 53624
rect 29748 53582 29776 53751
rect 29736 53576 29788 53582
rect 29736 53518 29788 53524
rect 29736 53440 29788 53446
rect 29736 53382 29788 53388
rect 29644 53100 29696 53106
rect 29644 53042 29696 53048
rect 29656 53009 29684 53042
rect 29748 53038 29776 53382
rect 29840 53122 29868 58278
rect 29932 56681 29960 60046
rect 30024 58682 30052 60706
rect 30104 58948 30156 58954
rect 30104 58890 30156 58896
rect 30012 58676 30064 58682
rect 30012 58618 30064 58624
rect 30012 58540 30064 58546
rect 30012 58482 30064 58488
rect 30024 56778 30052 58482
rect 30116 58342 30144 58890
rect 30104 58336 30156 58342
rect 30104 58278 30156 58284
rect 30104 57792 30156 57798
rect 30104 57734 30156 57740
rect 30012 56772 30064 56778
rect 30012 56714 30064 56720
rect 29918 56672 29974 56681
rect 29918 56607 29974 56616
rect 29920 56500 29972 56506
rect 29920 56442 29972 56448
rect 29932 55321 29960 56442
rect 30024 56370 30052 56714
rect 30012 56364 30064 56370
rect 30012 56306 30064 56312
rect 29918 55312 29974 55321
rect 30024 55282 30052 56306
rect 29918 55247 29974 55256
rect 30012 55276 30064 55282
rect 30012 55218 30064 55224
rect 30024 55078 30052 55218
rect 30012 55072 30064 55078
rect 30012 55014 30064 55020
rect 30024 54194 30052 55014
rect 30012 54188 30064 54194
rect 30012 54130 30064 54136
rect 30010 53136 30066 53145
rect 29840 53094 29960 53122
rect 29736 53032 29788 53038
rect 29642 53000 29698 53009
rect 29736 52974 29788 52980
rect 29642 52935 29698 52944
rect 29552 52352 29604 52358
rect 29552 52294 29604 52300
rect 29656 52086 29684 52935
rect 29828 52896 29880 52902
rect 29828 52838 29880 52844
rect 29736 52420 29788 52426
rect 29736 52362 29788 52368
rect 29644 52080 29696 52086
rect 29644 52022 29696 52028
rect 29644 51944 29696 51950
rect 29644 51886 29696 51892
rect 29460 51808 29512 51814
rect 29460 51750 29512 51756
rect 29550 51776 29606 51785
rect 29550 51711 29606 51720
rect 29460 51536 29512 51542
rect 29460 51478 29512 51484
rect 29368 51468 29420 51474
rect 29368 51410 29420 51416
rect 29366 51368 29422 51377
rect 29366 51303 29422 51312
rect 29380 46170 29408 51303
rect 29368 46164 29420 46170
rect 29368 46106 29420 46112
rect 29368 45960 29420 45966
rect 29368 45902 29420 45908
rect 29276 45348 29328 45354
rect 29276 45290 29328 45296
rect 29276 45008 29328 45014
rect 29276 44950 29328 44956
rect 29288 43217 29316 44950
rect 29380 43353 29408 45902
rect 29366 43344 29422 43353
rect 29366 43279 29422 43288
rect 29274 43208 29330 43217
rect 29274 43143 29330 43152
rect 29276 43104 29328 43110
rect 29276 43046 29328 43052
rect 29288 42945 29316 43046
rect 29274 42936 29330 42945
rect 29274 42871 29330 42880
rect 29472 42786 29500 51478
rect 29564 51066 29592 51711
rect 29656 51610 29684 51886
rect 29644 51604 29696 51610
rect 29644 51546 29696 51552
rect 29748 51513 29776 52362
rect 29734 51504 29790 51513
rect 29734 51439 29790 51448
rect 29642 51368 29698 51377
rect 29642 51303 29698 51312
rect 29656 51074 29684 51303
rect 29552 51060 29604 51066
rect 29656 51046 29776 51074
rect 29552 51002 29604 51008
rect 29644 50992 29696 50998
rect 29644 50934 29696 50940
rect 29552 48816 29604 48822
rect 29552 48758 29604 48764
rect 29564 48385 29592 48758
rect 29550 48376 29606 48385
rect 29550 48311 29606 48320
rect 29550 48240 29606 48249
rect 29550 48175 29606 48184
rect 29564 45554 29592 48175
rect 29656 45665 29684 50934
rect 29748 50425 29776 51046
rect 29840 50998 29868 52838
rect 29932 51649 29960 53094
rect 30010 53071 30012 53080
rect 30064 53071 30066 53080
rect 30012 53042 30064 53048
rect 30012 52692 30064 52698
rect 30012 52634 30064 52640
rect 30024 52086 30052 52634
rect 30012 52080 30064 52086
rect 30012 52022 30064 52028
rect 29918 51640 29974 51649
rect 29918 51575 29974 51584
rect 29920 51332 29972 51338
rect 29920 51274 29972 51280
rect 29828 50992 29880 50998
rect 29828 50934 29880 50940
rect 29932 50833 29960 51274
rect 29918 50824 29974 50833
rect 30116 50794 30144 57734
rect 30208 54330 30236 72014
rect 30840 71596 30892 71602
rect 30840 71538 30892 71544
rect 30288 70984 30340 70990
rect 30288 70926 30340 70932
rect 30300 55418 30328 70926
rect 30656 69896 30708 69902
rect 30656 69838 30708 69844
rect 30472 68332 30524 68338
rect 30472 68274 30524 68280
rect 30380 66020 30432 66026
rect 30380 65962 30432 65968
rect 30392 65074 30420 65962
rect 30380 65068 30432 65074
rect 30380 65010 30432 65016
rect 30380 64388 30432 64394
rect 30380 64330 30432 64336
rect 30392 63306 30420 64330
rect 30380 63300 30432 63306
rect 30380 63242 30432 63248
rect 30380 59220 30432 59226
rect 30380 59162 30432 59168
rect 30392 58546 30420 59162
rect 30380 58540 30432 58546
rect 30380 58482 30432 58488
rect 30380 58404 30432 58410
rect 30380 58346 30432 58352
rect 30288 55412 30340 55418
rect 30288 55354 30340 55360
rect 30286 55312 30342 55321
rect 30286 55247 30342 55256
rect 30300 54602 30328 55247
rect 30392 54874 30420 58346
rect 30380 54868 30432 54874
rect 30380 54810 30432 54816
rect 30380 54664 30432 54670
rect 30380 54606 30432 54612
rect 30288 54596 30340 54602
rect 30288 54538 30340 54544
rect 30300 54505 30328 54538
rect 30286 54496 30342 54505
rect 30286 54431 30342 54440
rect 30196 54324 30248 54330
rect 30196 54266 30248 54272
rect 30288 54052 30340 54058
rect 30288 53994 30340 54000
rect 30196 53984 30248 53990
rect 30196 53926 30248 53932
rect 29918 50759 29974 50768
rect 30104 50788 30156 50794
rect 30104 50730 30156 50736
rect 29828 50720 29880 50726
rect 29826 50688 29828 50697
rect 29920 50720 29972 50726
rect 29880 50688 29882 50697
rect 29920 50662 29972 50668
rect 29826 50623 29882 50632
rect 29734 50416 29790 50425
rect 29734 50351 29790 50360
rect 29736 50244 29788 50250
rect 29736 50186 29788 50192
rect 29748 50017 29776 50186
rect 29828 50176 29880 50182
rect 29826 50144 29828 50153
rect 29880 50144 29882 50153
rect 29826 50079 29882 50088
rect 29734 50008 29790 50017
rect 29734 49943 29790 49952
rect 29828 49904 29880 49910
rect 29828 49846 29880 49852
rect 29736 49768 29788 49774
rect 29736 49710 29788 49716
rect 29748 49473 29776 49710
rect 29734 49464 29790 49473
rect 29734 49399 29790 49408
rect 29736 49156 29788 49162
rect 29736 49098 29788 49104
rect 29748 47161 29776 49098
rect 29734 47152 29790 47161
rect 29734 47087 29790 47096
rect 29736 46980 29788 46986
rect 29736 46922 29788 46928
rect 29748 46753 29776 46922
rect 29734 46744 29790 46753
rect 29734 46679 29790 46688
rect 29736 46572 29788 46578
rect 29736 46514 29788 46520
rect 29748 46209 29776 46514
rect 29734 46200 29790 46209
rect 29734 46135 29790 46144
rect 29734 46064 29790 46073
rect 29734 45999 29790 46008
rect 29748 45966 29776 45999
rect 29736 45960 29788 45966
rect 29736 45902 29788 45908
rect 29642 45656 29698 45665
rect 29642 45591 29698 45600
rect 29748 45558 29776 45902
rect 29564 45526 29684 45554
rect 29552 45484 29604 45490
rect 29552 45426 29604 45432
rect 29564 43382 29592 45426
rect 29656 45014 29684 45526
rect 29736 45552 29788 45558
rect 29736 45494 29788 45500
rect 29644 45008 29696 45014
rect 29644 44950 29696 44956
rect 29748 44878 29776 45494
rect 29736 44872 29788 44878
rect 29736 44814 29788 44820
rect 29644 44736 29696 44742
rect 29644 44678 29696 44684
rect 29552 43376 29604 43382
rect 29552 43318 29604 43324
rect 29552 43104 29604 43110
rect 29552 43046 29604 43052
rect 29288 42758 29500 42786
rect 29182 42256 29238 42265
rect 29182 42191 29238 42200
rect 29092 42084 29144 42090
rect 29144 42044 29224 42072
rect 29092 42026 29144 42032
rect 29090 41984 29146 41993
rect 28920 41942 28994 41970
rect 28966 41834 28994 41942
rect 29090 41919 29146 41928
rect 28816 41812 28868 41818
rect 28816 41754 28868 41760
rect 28920 41806 28994 41834
rect 28816 41608 28868 41614
rect 28724 41586 28776 41592
rect 28816 41550 28868 41556
rect 28724 41528 28776 41534
rect 28722 41440 28778 41449
rect 28722 41375 28778 41384
rect 28736 41274 28764 41375
rect 28724 41268 28776 41274
rect 28724 41210 28776 41216
rect 28538 41103 28594 41112
rect 28625 41126 28672 41154
rect 28625 41052 28653 41126
rect 28552 41024 28653 41052
rect 28828 41041 28856 41550
rect 28920 41460 28948 41806
rect 29104 41562 29132 41919
rect 29196 41682 29224 42044
rect 29184 41676 29236 41682
rect 29184 41618 29236 41624
rect 29104 41534 29224 41562
rect 29092 41472 29144 41478
rect 28920 41432 29040 41460
rect 28908 41268 28960 41274
rect 28908 41210 28960 41216
rect 28920 41177 28948 41210
rect 28906 41168 28962 41177
rect 28906 41103 28962 41112
rect 29012 41052 29040 41432
rect 29092 41414 29144 41420
rect 28814 41032 28870 41041
rect 28552 40118 28580 41024
rect 28814 40967 28870 40976
rect 28920 41024 29040 41052
rect 28816 40928 28868 40934
rect 28630 40896 28686 40905
rect 28630 40831 28686 40840
rect 28736 40888 28816 40916
rect 28540 40112 28592 40118
rect 28540 40054 28592 40060
rect 28538 39808 28594 39817
rect 28538 39743 28594 39752
rect 28448 32768 28500 32774
rect 28448 32710 28500 32716
rect 28368 32524 28488 32552
rect 28276 32456 28396 32484
rect 28078 32263 28134 32272
rect 28172 32292 28224 32298
rect 28092 31890 28120 32263
rect 28172 32234 28224 32240
rect 28080 31884 28132 31890
rect 28080 31826 28132 31832
rect 28078 31784 28134 31793
rect 28078 31719 28134 31728
rect 28092 31385 28120 31719
rect 28078 31376 28134 31385
rect 28078 31311 28134 31320
rect 28080 30388 28132 30394
rect 28080 30330 28132 30336
rect 28092 30054 28120 30330
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 28184 29782 28212 32234
rect 28264 31952 28316 31958
rect 28264 31894 28316 31900
rect 28276 30802 28304 31894
rect 28368 30938 28396 32456
rect 28460 32026 28488 32524
rect 28448 32020 28500 32026
rect 28448 31962 28500 31968
rect 28446 31512 28502 31521
rect 28446 31447 28502 31456
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 28264 30796 28316 30802
rect 28264 30738 28316 30744
rect 28356 30388 28408 30394
rect 28356 30330 28408 30336
rect 28264 30048 28316 30054
rect 28262 30016 28264 30025
rect 28316 30016 28318 30025
rect 28262 29951 28318 29960
rect 27816 29702 27936 29730
rect 28172 29776 28224 29782
rect 28368 29753 28396 30330
rect 28172 29718 28224 29724
rect 28354 29744 28410 29753
rect 28080 29708 28132 29714
rect 27712 29572 27764 29578
rect 27712 29514 27764 29520
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27526 29336 27582 29345
rect 27526 29271 27582 29280
rect 27528 29096 27580 29102
rect 27528 29038 27580 29044
rect 27540 28801 27568 29038
rect 27632 28966 27660 29446
rect 27712 29300 27764 29306
rect 27712 29242 27764 29248
rect 27724 29170 27752 29242
rect 27712 29164 27764 29170
rect 27712 29106 27764 29112
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 27526 28792 27582 28801
rect 27526 28727 27582 28736
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 27632 28642 27660 28698
rect 27540 28614 27660 28642
rect 27540 28370 27568 28614
rect 27620 28552 27672 28558
rect 27724 28540 27752 29106
rect 27672 28512 27752 28540
rect 27620 28494 27672 28500
rect 27540 28342 27660 28370
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27528 27328 27580 27334
rect 27528 27270 27580 27276
rect 27344 27124 27396 27130
rect 27344 27066 27396 27072
rect 27252 27056 27304 27062
rect 27158 27024 27214 27033
rect 27252 26998 27304 27004
rect 27436 27056 27488 27062
rect 27436 26998 27488 27004
rect 27158 26959 27214 26968
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27250 26888 27306 26897
rect 27068 19916 27120 19922
rect 27068 19858 27120 19864
rect 27066 19816 27122 19825
rect 27066 19751 27122 19760
rect 27080 17202 27108 19751
rect 27068 17196 27120 17202
rect 27068 17138 27120 17144
rect 27080 16182 27108 17138
rect 27068 16176 27120 16182
rect 27068 16118 27120 16124
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 27080 14550 27108 14962
rect 27068 14544 27120 14550
rect 27068 14486 27120 14492
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 27080 10062 27108 13126
rect 27172 11218 27200 26862
rect 27250 26823 27306 26832
rect 27264 21962 27292 26823
rect 27356 25974 27384 26930
rect 27448 26926 27476 26998
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27448 26761 27476 26862
rect 27434 26752 27490 26761
rect 27434 26687 27490 26696
rect 27434 26616 27490 26625
rect 27434 26551 27490 26560
rect 27448 26518 27476 26551
rect 27436 26512 27488 26518
rect 27436 26454 27488 26460
rect 27436 26308 27488 26314
rect 27436 26250 27488 26256
rect 27344 25968 27396 25974
rect 27344 25910 27396 25916
rect 27356 25498 27384 25910
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27344 25356 27396 25362
rect 27344 25298 27396 25304
rect 27356 24614 27384 25298
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 27344 24404 27396 24410
rect 27344 24346 27396 24352
rect 27252 21956 27304 21962
rect 27252 21898 27304 21904
rect 27250 21856 27306 21865
rect 27250 21791 27306 21800
rect 27264 19938 27292 21791
rect 27356 21622 27384 24346
rect 27448 22273 27476 26250
rect 27540 25158 27568 27270
rect 27632 25430 27660 28342
rect 27710 27976 27766 27985
rect 27710 27911 27712 27920
rect 27764 27911 27766 27920
rect 27712 27882 27764 27888
rect 27710 27568 27766 27577
rect 27710 27503 27712 27512
rect 27764 27503 27766 27512
rect 27712 27474 27764 27480
rect 27710 27432 27766 27441
rect 27710 27367 27766 27376
rect 27724 26382 27752 27367
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27816 26024 27844 29702
rect 28080 29650 28132 29656
rect 27894 29608 27950 29617
rect 28092 29594 28120 29650
rect 27950 29566 28120 29594
rect 27894 29543 27950 29552
rect 28000 29170 28028 29566
rect 28078 29472 28134 29481
rect 28078 29407 28134 29416
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 27894 28928 27950 28937
rect 27894 28863 27950 28872
rect 27724 25996 27844 26024
rect 27620 25424 27672 25430
rect 27620 25366 27672 25372
rect 27618 25256 27674 25265
rect 27618 25191 27620 25200
rect 27672 25191 27674 25200
rect 27620 25162 27672 25168
rect 27528 25152 27580 25158
rect 27528 25094 27580 25100
rect 27632 24970 27660 25162
rect 27540 24942 27660 24970
rect 27540 24410 27568 24942
rect 27620 24744 27672 24750
rect 27620 24686 27672 24692
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27632 23798 27660 24686
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27632 23186 27660 23734
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 27632 22710 27660 22986
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27632 22386 27660 22646
rect 27540 22358 27660 22386
rect 27724 22386 27752 25996
rect 27804 25900 27856 25906
rect 27804 25842 27856 25848
rect 27816 24886 27844 25842
rect 27804 24880 27856 24886
rect 27804 24822 27856 24828
rect 27816 24410 27844 24822
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27804 24064 27856 24070
rect 27802 24032 27804 24041
rect 27856 24032 27858 24041
rect 27802 23967 27858 23976
rect 27802 23760 27858 23769
rect 27802 23695 27858 23704
rect 27816 23662 27844 23695
rect 27804 23656 27856 23662
rect 27804 23598 27856 23604
rect 27724 22358 27844 22386
rect 27434 22264 27490 22273
rect 27540 22234 27568 22358
rect 27434 22199 27490 22208
rect 27528 22228 27580 22234
rect 27816 22216 27844 22358
rect 27528 22170 27580 22176
rect 27632 22188 27844 22216
rect 27436 22160 27488 22166
rect 27436 22102 27488 22108
rect 27526 22128 27582 22137
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 27448 21146 27476 22102
rect 27526 22063 27582 22072
rect 27436 21140 27488 21146
rect 27436 21082 27488 21088
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 27264 19910 27384 19938
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27264 13138 27292 19790
rect 27356 18329 27384 19910
rect 27448 19446 27476 20266
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 27342 18320 27398 18329
rect 27342 18255 27398 18264
rect 27344 18216 27396 18222
rect 27344 18158 27396 18164
rect 27356 16454 27384 18158
rect 27448 17270 27476 19382
rect 27540 18902 27568 22063
rect 27632 21570 27660 22188
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27724 21690 27752 22034
rect 27802 21992 27858 22001
rect 27802 21927 27804 21936
rect 27856 21927 27858 21936
rect 27804 21898 27856 21904
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27632 21542 27752 21570
rect 27618 21312 27674 21321
rect 27618 21247 27674 21256
rect 27632 20942 27660 21247
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27528 18896 27580 18902
rect 27528 18838 27580 18844
rect 27526 18728 27582 18737
rect 27526 18663 27582 18672
rect 27540 17338 27568 18663
rect 27724 18306 27752 21542
rect 27804 19780 27856 19786
rect 27804 19722 27856 19728
rect 27632 18278 27752 18306
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27436 17264 27488 17270
rect 27436 17206 27488 17212
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 27356 14550 27384 16118
rect 27448 16046 27476 17206
rect 27632 16794 27660 18278
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27436 15496 27488 15502
rect 27436 15438 27488 15444
rect 27448 15162 27476 15438
rect 27540 15366 27568 16594
rect 27632 16454 27660 16730
rect 27724 16522 27752 17070
rect 27712 16516 27764 16522
rect 27712 16458 27764 16464
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27618 16280 27674 16289
rect 27618 16215 27674 16224
rect 27632 16182 27660 16215
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27724 15570 27752 16458
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27618 15464 27674 15473
rect 27618 15399 27620 15408
rect 27672 15399 27674 15408
rect 27620 15370 27672 15376
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27540 15178 27568 15302
rect 27436 15156 27488 15162
rect 27540 15150 27752 15178
rect 27436 15098 27488 15104
rect 27620 15088 27672 15094
rect 27620 15030 27672 15036
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27344 14544 27396 14550
rect 27344 14486 27396 14492
rect 27448 14006 27476 14758
rect 27540 14482 27568 14894
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27436 13524 27488 13530
rect 27436 13466 27488 13472
rect 27448 13190 27476 13466
rect 27436 13184 27488 13190
rect 27264 13110 27384 13138
rect 27436 13126 27488 13132
rect 27252 12980 27304 12986
rect 27252 12922 27304 12928
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27264 11098 27292 12922
rect 27172 11070 27292 11098
rect 27068 10056 27120 10062
rect 27068 9998 27120 10004
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 27080 8634 27108 9522
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 27080 8498 27108 8570
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27080 8022 27108 8434
rect 27068 8016 27120 8022
rect 27068 7958 27120 7964
rect 26988 7534 27108 7562
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26988 6934 27016 7346
rect 26976 6928 27028 6934
rect 26976 6870 27028 6876
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25792 5166 25820 5646
rect 25504 5160 25556 5166
rect 25504 5102 25556 5108
rect 25780 5160 25832 5166
rect 25780 5102 25832 5108
rect 26148 5160 26200 5166
rect 26148 5102 26200 5108
rect 25776 4924 26084 4944
rect 25776 4922 25782 4924
rect 25838 4922 25862 4924
rect 25918 4922 25942 4924
rect 25998 4922 26022 4924
rect 26078 4922 26084 4924
rect 25838 4870 25840 4922
rect 26020 4870 26022 4922
rect 25776 4868 25782 4870
rect 25838 4868 25862 4870
rect 25918 4868 25942 4870
rect 25998 4868 26022 4870
rect 26078 4868 26084 4870
rect 25776 4848 26084 4868
rect 26160 4690 26188 5102
rect 26148 4684 26200 4690
rect 26148 4626 26200 4632
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25136 4480 25188 4486
rect 25136 4422 25188 4428
rect 25148 3534 25176 4422
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 25424 3398 25452 4558
rect 25776 3836 26084 3856
rect 25776 3834 25782 3836
rect 25838 3834 25862 3836
rect 25918 3834 25942 3836
rect 25998 3834 26022 3836
rect 26078 3834 26084 3836
rect 25838 3782 25840 3834
rect 26020 3782 26022 3834
rect 25776 3780 25782 3782
rect 25838 3780 25862 3782
rect 25918 3780 25942 3782
rect 25998 3780 26022 3782
rect 26078 3780 26084 3782
rect 25776 3760 26084 3780
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 26620 3126 26648 5646
rect 27080 5234 27108 7534
rect 27172 5574 27200 11070
rect 27252 10532 27304 10538
rect 27252 10474 27304 10480
rect 27264 8838 27292 10474
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27264 6662 27292 8774
rect 27356 8294 27384 13110
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27448 12442 27476 12786
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27540 12306 27568 14418
rect 27632 13841 27660 15030
rect 27618 13832 27674 13841
rect 27724 13802 27752 15150
rect 27816 14414 27844 19722
rect 27908 16289 27936 28863
rect 28000 28558 28028 29106
rect 28092 28558 28120 29407
rect 28184 29306 28212 29718
rect 28354 29679 28410 29688
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28368 29306 28396 29582
rect 28172 29300 28224 29306
rect 28172 29242 28224 29248
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28170 29200 28226 29209
rect 28170 29135 28226 29144
rect 28356 29164 28408 29170
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 28080 28552 28132 28558
rect 28080 28494 28132 28500
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 28000 25106 28028 28358
rect 28092 27606 28120 28494
rect 28080 27600 28132 27606
rect 28080 27542 28132 27548
rect 28080 27328 28132 27334
rect 28080 27270 28132 27276
rect 28092 27062 28120 27270
rect 28080 27056 28132 27062
rect 28080 26998 28132 27004
rect 28092 26518 28120 26998
rect 28080 26512 28132 26518
rect 28080 26454 28132 26460
rect 28092 26314 28120 26454
rect 28080 26308 28132 26314
rect 28080 26250 28132 26256
rect 28080 25900 28132 25906
rect 28080 25842 28132 25848
rect 28092 25294 28120 25842
rect 28184 25498 28212 29135
rect 28356 29106 28408 29112
rect 28264 27532 28316 27538
rect 28264 27474 28316 27480
rect 28172 25492 28224 25498
rect 28172 25434 28224 25440
rect 28080 25288 28132 25294
rect 28080 25230 28132 25236
rect 28000 25078 28120 25106
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 28000 23594 28028 24550
rect 27988 23588 28040 23594
rect 27988 23530 28040 23536
rect 28000 19854 28028 23530
rect 28092 21865 28120 25078
rect 28276 24698 28304 27474
rect 28368 25242 28396 29106
rect 28460 28422 28488 31447
rect 28448 28416 28500 28422
rect 28448 28358 28500 28364
rect 28448 28212 28500 28218
rect 28448 28154 28500 28160
rect 28460 28082 28488 28154
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28448 27464 28500 27470
rect 28446 27432 28448 27441
rect 28500 27432 28502 27441
rect 28446 27367 28502 27376
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28460 25906 28488 27270
rect 28448 25900 28500 25906
rect 28448 25842 28500 25848
rect 28368 25214 28488 25242
rect 28354 25120 28410 25129
rect 28354 25055 28410 25064
rect 28184 24670 28304 24698
rect 28078 21856 28134 21865
rect 28078 21791 28134 21800
rect 28184 21706 28212 24670
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28276 22030 28304 24550
rect 28368 24206 28396 25055
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28460 24052 28488 25214
rect 28368 24024 28488 24052
rect 28264 22024 28316 22030
rect 28264 21966 28316 21972
rect 28092 21678 28212 21706
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28000 18834 28028 19790
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 28000 18358 28028 18770
rect 27988 18352 28040 18358
rect 27988 18294 28040 18300
rect 27988 17332 28040 17338
rect 27988 17274 28040 17280
rect 27894 16280 27950 16289
rect 27894 16215 27950 16224
rect 28000 16096 28028 17274
rect 27908 16068 28028 16096
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 27618 13767 27674 13776
rect 27712 13796 27764 13802
rect 27712 13738 27764 13744
rect 27528 12300 27580 12306
rect 27528 12242 27580 12248
rect 27540 11626 27568 12242
rect 27816 11898 27844 14350
rect 27908 13954 27936 16068
rect 27988 15904 28040 15910
rect 27988 15846 28040 15852
rect 28000 15026 28028 15846
rect 28092 15026 28120 21678
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 28184 20534 28212 21490
rect 28264 20936 28316 20942
rect 28262 20904 28264 20913
rect 28316 20904 28318 20913
rect 28262 20839 28318 20848
rect 28172 20528 28224 20534
rect 28172 20470 28224 20476
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28184 19446 28212 20198
rect 28264 19916 28316 19922
rect 28264 19858 28316 19864
rect 28276 19514 28304 19858
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 28172 18896 28224 18902
rect 28172 18838 28224 18844
rect 28184 17270 28212 18838
rect 28368 18426 28396 24024
rect 28448 23792 28500 23798
rect 28448 23734 28500 23740
rect 28460 22234 28488 23734
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28446 22128 28502 22137
rect 28446 22063 28502 22072
rect 28460 21962 28488 22063
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28446 21856 28502 21865
rect 28446 21791 28502 21800
rect 28460 18902 28488 21791
rect 28448 18896 28500 18902
rect 28448 18838 28500 18844
rect 28448 18692 28500 18698
rect 28448 18634 28500 18640
rect 28356 18420 28408 18426
rect 28356 18362 28408 18368
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28172 17264 28224 17270
rect 28172 17206 28224 17212
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 27988 14544 28040 14550
rect 27986 14512 27988 14521
rect 28040 14512 28042 14521
rect 27986 14447 28042 14456
rect 28092 14074 28120 14962
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 27908 13926 28120 13954
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27804 11892 27856 11898
rect 27804 11834 27856 11840
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 27540 11354 27568 11562
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27436 11212 27488 11218
rect 27436 11154 27488 11160
rect 27448 9586 27476 11154
rect 27540 10606 27568 11290
rect 27632 10742 27660 11834
rect 28092 10810 28120 13926
rect 28184 13258 28212 17206
rect 28276 16590 28304 18226
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28368 17513 28396 17614
rect 28354 17504 28410 17513
rect 28354 17439 28410 17448
rect 28264 16584 28316 16590
rect 28264 16526 28316 16532
rect 28276 15706 28304 16526
rect 28356 16244 28408 16250
rect 28356 16186 28408 16192
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 28262 15192 28318 15201
rect 28262 15127 28264 15136
rect 28316 15127 28318 15136
rect 28264 15098 28316 15104
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28172 13252 28224 13258
rect 28172 13194 28224 13200
rect 28184 12434 28212 13194
rect 28276 12986 28304 14418
rect 28368 12986 28396 16186
rect 28460 16114 28488 18634
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28460 15910 28488 16050
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28552 15722 28580 39743
rect 28644 39098 28672 40831
rect 28632 39092 28684 39098
rect 28632 39034 28684 39040
rect 28632 38752 28684 38758
rect 28632 38694 28684 38700
rect 28644 38321 28672 38694
rect 28630 38312 28686 38321
rect 28630 38247 28686 38256
rect 28630 38040 28686 38049
rect 28630 37975 28686 37984
rect 28644 37398 28672 37975
rect 28736 37777 28764 40888
rect 28816 40870 28868 40876
rect 28816 40112 28868 40118
rect 28816 40054 28868 40060
rect 28828 38010 28856 40054
rect 28920 39642 28948 41024
rect 28998 40896 29054 40905
rect 28998 40831 29054 40840
rect 29012 40458 29040 40831
rect 29000 40452 29052 40458
rect 29000 40394 29052 40400
rect 28908 39636 28960 39642
rect 28908 39578 28960 39584
rect 28908 39296 28960 39302
rect 28908 39238 28960 39244
rect 28920 38729 28948 39238
rect 29000 39024 29052 39030
rect 29000 38966 29052 38972
rect 28906 38720 28962 38729
rect 28906 38655 28962 38664
rect 28908 38548 28960 38554
rect 28908 38490 28960 38496
rect 28816 38004 28868 38010
rect 28816 37946 28868 37952
rect 28920 37890 28948 38490
rect 28828 37862 28948 37890
rect 28722 37768 28778 37777
rect 28722 37703 28778 37712
rect 28724 37664 28776 37670
rect 28724 37606 28776 37612
rect 28632 37392 28684 37398
rect 28632 37334 28684 37340
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 28644 36786 28672 37198
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28736 36666 28764 37606
rect 28644 36638 28764 36666
rect 28644 36038 28672 36638
rect 28724 36576 28776 36582
rect 28724 36518 28776 36524
rect 28632 36032 28684 36038
rect 28632 35974 28684 35980
rect 28736 32910 28764 36518
rect 28828 35766 28856 37862
rect 29012 37754 29040 38966
rect 28920 37726 29040 37754
rect 28816 35760 28868 35766
rect 28816 35702 28868 35708
rect 28816 35624 28868 35630
rect 28816 35566 28868 35572
rect 28828 35290 28856 35566
rect 28816 35284 28868 35290
rect 28816 35226 28868 35232
rect 28920 34898 28948 37726
rect 29000 37664 29052 37670
rect 29000 37606 29052 37612
rect 29012 36786 29040 37606
rect 29104 37262 29132 41414
rect 29196 39302 29224 41534
rect 29184 39296 29236 39302
rect 29184 39238 29236 39244
rect 29184 38344 29236 38350
rect 29184 38286 29236 38292
rect 29196 37466 29224 38286
rect 29184 37460 29236 37466
rect 29184 37402 29236 37408
rect 29092 37256 29144 37262
rect 29092 37198 29144 37204
rect 29184 36848 29236 36854
rect 29184 36790 29236 36796
rect 29000 36780 29052 36786
rect 29000 36722 29052 36728
rect 29092 36780 29144 36786
rect 29092 36722 29144 36728
rect 29000 36644 29052 36650
rect 29000 36586 29052 36592
rect 28828 34870 28948 34898
rect 28828 34388 28856 34870
rect 28908 34740 28960 34746
rect 28908 34682 28960 34688
rect 28920 34513 28948 34682
rect 29012 34542 29040 36586
rect 29104 35630 29132 36722
rect 29196 36038 29224 36790
rect 29184 36032 29236 36038
rect 29184 35974 29236 35980
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 29104 34610 29132 35566
rect 29184 34740 29236 34746
rect 29184 34682 29236 34688
rect 29092 34604 29144 34610
rect 29092 34546 29144 34552
rect 29000 34536 29052 34542
rect 28906 34504 28962 34513
rect 29000 34478 29052 34484
rect 28906 34439 28962 34448
rect 28828 34360 29040 34388
rect 28816 33992 28868 33998
rect 28816 33934 28868 33940
rect 28724 32904 28776 32910
rect 28724 32846 28776 32852
rect 28632 32768 28684 32774
rect 28632 32710 28684 32716
rect 28722 32736 28778 32745
rect 28644 32314 28672 32710
rect 28722 32671 28778 32680
rect 28736 32434 28764 32671
rect 28828 32609 28856 33934
rect 28908 33856 28960 33862
rect 28908 33798 28960 33804
rect 28920 33561 28948 33798
rect 28906 33552 28962 33561
rect 28906 33487 28962 33496
rect 28908 32768 28960 32774
rect 28908 32710 28960 32716
rect 28814 32600 28870 32609
rect 28814 32535 28870 32544
rect 28724 32428 28776 32434
rect 28724 32370 28776 32376
rect 28644 32286 28856 32314
rect 28630 32056 28686 32065
rect 28630 31991 28686 32000
rect 28644 30734 28672 31991
rect 28724 31884 28776 31890
rect 28724 31826 28776 31832
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28736 30682 28764 31826
rect 28828 30841 28856 32286
rect 28920 32201 28948 32710
rect 29012 32609 29040 34360
rect 28998 32600 29054 32609
rect 28998 32535 29054 32544
rect 29196 32450 29224 34682
rect 29288 33402 29316 42758
rect 29564 42684 29592 43046
rect 29366 42664 29422 42673
rect 29366 42599 29422 42608
rect 29472 42656 29592 42684
rect 29656 42673 29684 44678
rect 29840 44554 29868 49846
rect 29748 44526 29868 44554
rect 29748 42684 29776 44526
rect 29828 44396 29880 44402
rect 29828 44338 29880 44344
rect 29840 43897 29868 44338
rect 29826 43888 29882 43897
rect 29826 43823 29882 43832
rect 29828 43784 29880 43790
rect 29828 43726 29880 43732
rect 29840 43489 29868 43726
rect 29932 43625 29960 50662
rect 30012 49768 30064 49774
rect 30012 49710 30064 49716
rect 30024 48686 30052 49710
rect 30012 48680 30064 48686
rect 30012 48622 30064 48628
rect 30024 47734 30052 48622
rect 30102 48376 30158 48385
rect 30102 48311 30158 48320
rect 30012 47728 30064 47734
rect 30012 47670 30064 47676
rect 30012 45960 30064 45966
rect 30012 45902 30064 45908
rect 30024 45422 30052 45902
rect 30012 45416 30064 45422
rect 30012 45358 30064 45364
rect 30024 44878 30052 45358
rect 30012 44872 30064 44878
rect 30012 44814 30064 44820
rect 30010 44568 30066 44577
rect 30010 44503 30012 44512
rect 30064 44503 30066 44512
rect 30012 44474 30064 44480
rect 30010 44296 30066 44305
rect 30010 44231 30012 44240
rect 30064 44231 30066 44240
rect 30012 44202 30064 44208
rect 30012 43648 30064 43654
rect 29918 43616 29974 43625
rect 30012 43590 30064 43596
rect 29918 43551 29974 43560
rect 29826 43480 29882 43489
rect 29826 43415 29882 43424
rect 29828 43376 29880 43382
rect 29828 43318 29880 43324
rect 29840 42906 29868 43318
rect 29920 43308 29972 43314
rect 29920 43250 29972 43256
rect 29828 42900 29880 42906
rect 29828 42842 29880 42848
rect 29642 42664 29698 42673
rect 29380 38842 29408 42599
rect 29472 42129 29500 42656
rect 29748 42656 29868 42684
rect 29642 42599 29698 42608
rect 29644 42560 29696 42566
rect 29644 42502 29696 42508
rect 29736 42560 29788 42566
rect 29736 42502 29788 42508
rect 29550 42392 29606 42401
rect 29656 42362 29684 42502
rect 29748 42362 29776 42502
rect 29550 42327 29606 42336
rect 29644 42356 29696 42362
rect 29458 42120 29514 42129
rect 29458 42055 29514 42064
rect 29460 42016 29512 42022
rect 29460 41958 29512 41964
rect 29472 39438 29500 41958
rect 29564 41177 29592 42327
rect 29644 42298 29696 42304
rect 29736 42356 29788 42362
rect 29736 42298 29788 42304
rect 29734 42256 29790 42265
rect 29734 42191 29790 42200
rect 29644 42084 29696 42090
rect 29644 42026 29696 42032
rect 29550 41168 29606 41177
rect 29550 41103 29606 41112
rect 29550 41032 29606 41041
rect 29550 40967 29606 40976
rect 29460 39432 29512 39438
rect 29460 39374 29512 39380
rect 29380 38814 29500 38842
rect 29368 38752 29420 38758
rect 29368 38694 29420 38700
rect 29380 37369 29408 38694
rect 29472 38185 29500 38814
rect 29458 38176 29514 38185
rect 29458 38111 29514 38120
rect 29460 37868 29512 37874
rect 29460 37810 29512 37816
rect 29366 37360 29422 37369
rect 29366 37295 29422 37304
rect 29472 37262 29500 37810
rect 29564 37466 29592 40967
rect 29656 40497 29684 42026
rect 29748 41449 29776 42191
rect 29840 41818 29868 42656
rect 29932 42537 29960 43250
rect 30024 42809 30052 43590
rect 30116 43382 30144 48311
rect 30104 43376 30156 43382
rect 30104 43318 30156 43324
rect 30104 43240 30156 43246
rect 30104 43182 30156 43188
rect 30010 42800 30066 42809
rect 30010 42735 30066 42744
rect 30116 42684 30144 43182
rect 30024 42656 30144 42684
rect 29918 42528 29974 42537
rect 29918 42463 29974 42472
rect 29920 42220 29972 42226
rect 29920 42162 29972 42168
rect 29932 42090 29960 42162
rect 30024 42129 30052 42656
rect 30104 42356 30156 42362
rect 30104 42298 30156 42304
rect 30010 42120 30066 42129
rect 29920 42084 29972 42090
rect 30010 42055 30066 42064
rect 29920 42026 29972 42032
rect 30012 42016 30064 42022
rect 30012 41958 30064 41964
rect 29828 41812 29880 41818
rect 29828 41754 29880 41760
rect 29920 41608 29972 41614
rect 30024 41596 30052 41958
rect 30116 41614 30144 42298
rect 29972 41568 30052 41596
rect 30104 41608 30156 41614
rect 29920 41550 29972 41556
rect 30104 41550 30156 41556
rect 30104 41472 30156 41478
rect 29734 41440 29790 41449
rect 29734 41375 29790 41384
rect 30010 41440 30066 41449
rect 30104 41414 30156 41420
rect 30010 41375 30066 41384
rect 29748 41138 29960 41154
rect 29748 41132 29972 41138
rect 29748 41126 29920 41132
rect 29642 40488 29698 40497
rect 29642 40423 29698 40432
rect 29644 39296 29696 39302
rect 29644 39238 29696 39244
rect 29552 37460 29604 37466
rect 29552 37402 29604 37408
rect 29552 37324 29604 37330
rect 29552 37266 29604 37272
rect 29460 37256 29512 37262
rect 29380 37216 29460 37244
rect 29380 36242 29408 37216
rect 29460 37198 29512 37204
rect 29460 37120 29512 37126
rect 29460 37062 29512 37068
rect 29368 36236 29420 36242
rect 29368 36178 29420 36184
rect 29368 36032 29420 36038
rect 29368 35974 29420 35980
rect 29380 33862 29408 35974
rect 29368 33856 29420 33862
rect 29368 33798 29420 33804
rect 29288 33374 29408 33402
rect 29276 33312 29328 33318
rect 29276 33254 29328 33260
rect 29288 33153 29316 33254
rect 29274 33144 29330 33153
rect 29274 33079 29330 33088
rect 29380 32450 29408 33374
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 29104 32422 29224 32450
rect 29288 32422 29408 32450
rect 28906 32192 28962 32201
rect 28906 32127 28962 32136
rect 29012 32065 29040 32370
rect 28998 32056 29054 32065
rect 28998 31991 29054 32000
rect 28998 31920 29054 31929
rect 28998 31855 29054 31864
rect 28814 30832 28870 30841
rect 28814 30767 28870 30776
rect 28644 29034 28672 30670
rect 28736 30654 28856 30682
rect 28724 30592 28776 30598
rect 28724 30534 28776 30540
rect 28632 29028 28684 29034
rect 28632 28970 28684 28976
rect 28644 28626 28672 28970
rect 28632 28620 28684 28626
rect 28632 28562 28684 28568
rect 28644 28218 28672 28562
rect 28632 28212 28684 28218
rect 28632 28154 28684 28160
rect 28630 27432 28686 27441
rect 28630 27367 28686 27376
rect 28644 26042 28672 27367
rect 28632 26036 28684 26042
rect 28632 25978 28684 25984
rect 28630 25936 28686 25945
rect 28630 25871 28686 25880
rect 28644 24410 28672 25871
rect 28736 24614 28764 30534
rect 28828 28762 28856 30654
rect 28906 30424 28962 30433
rect 28906 30359 28962 30368
rect 28920 30190 28948 30359
rect 28908 30184 28960 30190
rect 28908 30126 28960 30132
rect 28908 29504 28960 29510
rect 28908 29446 28960 29452
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 28920 28529 28948 29446
rect 28906 28520 28962 28529
rect 29012 28506 29040 31855
rect 29104 30734 29132 32422
rect 29182 32328 29238 32337
rect 29182 32263 29238 32272
rect 29092 30728 29144 30734
rect 29092 30670 29144 30676
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 29104 28626 29132 30534
rect 29092 28620 29144 28626
rect 29092 28562 29144 28568
rect 29012 28478 29132 28506
rect 28906 28455 28962 28464
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 29012 28234 29040 28358
rect 28920 28206 29040 28234
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28724 24608 28776 24614
rect 28724 24550 28776 24556
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28722 23896 28778 23905
rect 28722 23831 28778 23840
rect 28632 23724 28684 23730
rect 28632 23666 28684 23672
rect 28644 23633 28672 23666
rect 28630 23624 28686 23633
rect 28630 23559 28686 23568
rect 28736 23526 28764 23831
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 28632 22568 28684 22574
rect 28632 22510 28684 22516
rect 28644 22098 28672 22510
rect 28736 22438 28764 23462
rect 28724 22432 28776 22438
rect 28724 22374 28776 22380
rect 28632 22092 28684 22098
rect 28828 22094 28856 28018
rect 28920 27470 28948 28206
rect 28998 27840 29054 27849
rect 28998 27775 29054 27784
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28920 26625 28948 27270
rect 28906 26616 28962 26625
rect 28906 26551 28962 26560
rect 28908 26512 28960 26518
rect 28908 26454 28960 26460
rect 28920 26081 28948 26454
rect 28906 26072 28962 26081
rect 28906 26007 28962 26016
rect 28906 25936 28962 25945
rect 28906 25871 28962 25880
rect 28920 24954 28948 25871
rect 29012 25430 29040 27775
rect 29104 26042 29132 28478
rect 29196 27130 29224 32263
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 29184 26852 29236 26858
rect 29184 26794 29236 26800
rect 29092 26036 29144 26042
rect 29092 25978 29144 25984
rect 29090 25800 29146 25809
rect 29090 25735 29146 25744
rect 29000 25424 29052 25430
rect 29000 25366 29052 25372
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 28908 24948 28960 24954
rect 28908 24890 28960 24896
rect 29012 24585 29040 25230
rect 29104 24954 29132 25735
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29092 24744 29144 24750
rect 29092 24686 29144 24692
rect 28998 24576 29054 24585
rect 28998 24511 29054 24520
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 28908 24200 28960 24206
rect 28906 24168 28908 24177
rect 28960 24168 28962 24177
rect 28906 24103 28962 24112
rect 29012 23594 29040 24346
rect 29000 23588 29052 23594
rect 29000 23530 29052 23536
rect 28908 23112 28960 23118
rect 29104 23100 29132 24686
rect 29196 24410 29224 26794
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 29196 23225 29224 23666
rect 29182 23216 29238 23225
rect 29182 23151 29238 23160
rect 29104 23072 29224 23100
rect 28908 23054 28960 23060
rect 28920 22409 28948 23054
rect 29000 23044 29052 23050
rect 29000 22986 29052 22992
rect 29012 22642 29040 22986
rect 29092 22976 29144 22982
rect 29092 22918 29144 22924
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 28906 22400 28962 22409
rect 28906 22335 28962 22344
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 28632 22034 28684 22040
rect 28736 22066 28856 22094
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28644 18766 28672 21558
rect 28736 20058 28764 22066
rect 28816 21956 28868 21962
rect 28816 21898 28868 21904
rect 28828 21570 28856 21898
rect 28920 21865 28948 22170
rect 28906 21856 28962 21865
rect 28906 21791 28962 21800
rect 29012 21690 29040 22578
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 28828 21542 29040 21570
rect 28816 20868 28868 20874
rect 28816 20810 28868 20816
rect 28724 20052 28776 20058
rect 28724 19994 28776 20000
rect 28722 19816 28778 19825
rect 28722 19751 28778 19760
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28644 17882 28672 18702
rect 28632 17876 28684 17882
rect 28632 17818 28684 17824
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28460 15694 28580 15722
rect 28264 12980 28316 12986
rect 28264 12922 28316 12928
rect 28356 12980 28408 12986
rect 28356 12922 28408 12928
rect 28460 12918 28488 15694
rect 28538 14104 28594 14113
rect 28538 14039 28594 14048
rect 28552 14006 28580 14039
rect 28644 14006 28672 17682
rect 28736 17338 28764 19751
rect 28828 19417 28856 20810
rect 28906 20360 28962 20369
rect 28906 20295 28962 20304
rect 28814 19408 28870 19417
rect 28920 19378 28948 20295
rect 29012 20058 29040 21542
rect 29000 20052 29052 20058
rect 29000 19994 29052 20000
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 28814 19343 28870 19352
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28908 19236 28960 19242
rect 28908 19178 28960 19184
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28724 17332 28776 17338
rect 28724 17274 28776 17280
rect 28828 17105 28856 17614
rect 28920 17542 28948 19178
rect 29012 18834 29040 19382
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 29012 18290 29040 18770
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 28998 18184 29054 18193
rect 28998 18119 29054 18128
rect 28908 17536 28960 17542
rect 28908 17478 28960 17484
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 28814 17096 28870 17105
rect 28814 17031 28870 17040
rect 28920 16697 28948 17138
rect 28906 16688 28962 16697
rect 28816 16652 28868 16658
rect 28906 16623 28962 16632
rect 28816 16594 28868 16600
rect 28724 16516 28776 16522
rect 28724 16458 28776 16464
rect 28736 16182 28764 16458
rect 28724 16176 28776 16182
rect 28724 16118 28776 16124
rect 28724 14340 28776 14346
rect 28724 14282 28776 14288
rect 28540 14000 28592 14006
rect 28540 13942 28592 13948
rect 28632 14000 28684 14006
rect 28632 13942 28684 13948
rect 28448 12912 28500 12918
rect 28448 12854 28500 12860
rect 28184 12406 28304 12434
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28184 11937 28212 12174
rect 28170 11928 28226 11937
rect 28170 11863 28226 11872
rect 28276 11150 28304 12406
rect 28460 11354 28488 12854
rect 28448 11348 28500 11354
rect 28448 11290 28500 11296
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 28276 10062 28304 11086
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27448 6662 27476 8910
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27252 6656 27304 6662
rect 27252 6598 27304 6604
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27540 6474 27568 8434
rect 27896 8288 27948 8294
rect 27896 8230 27948 8236
rect 27710 7712 27766 7721
rect 27710 7647 27766 7656
rect 27618 7168 27674 7177
rect 27618 7103 27674 7112
rect 27632 6798 27660 7103
rect 27724 6866 27752 7647
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27448 6446 27568 6474
rect 27160 5568 27212 5574
rect 27160 5510 27212 5516
rect 27448 5522 27476 6446
rect 27448 5494 27568 5522
rect 27068 5228 27120 5234
rect 27068 5170 27120 5176
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 26884 4752 26936 4758
rect 26884 4694 26936 4700
rect 26608 3120 26660 3126
rect 26608 3062 26660 3068
rect 25776 2748 26084 2768
rect 25776 2746 25782 2748
rect 25838 2746 25862 2748
rect 25918 2746 25942 2748
rect 25998 2746 26022 2748
rect 26078 2746 26084 2748
rect 25838 2694 25840 2746
rect 26020 2694 26022 2746
rect 25776 2692 25782 2694
rect 25838 2692 25862 2694
rect 25918 2692 25942 2694
rect 25998 2692 26022 2694
rect 26078 2692 26084 2694
rect 25776 2672 26084 2692
rect 26896 2650 26924 4694
rect 27448 4146 27476 4966
rect 27436 4140 27488 4146
rect 27436 4082 27488 4088
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 27264 3602 27292 3878
rect 27252 3596 27304 3602
rect 27252 3538 27304 3544
rect 27540 3194 27568 5494
rect 27712 5024 27764 5030
rect 27712 4966 27764 4972
rect 27724 4690 27752 4966
rect 27712 4684 27764 4690
rect 27712 4626 27764 4632
rect 27804 4616 27856 4622
rect 27804 4558 27856 4564
rect 27712 4480 27764 4486
rect 27816 4457 27844 4558
rect 27712 4422 27764 4428
rect 27802 4448 27858 4457
rect 27724 4282 27752 4422
rect 27802 4383 27858 4392
rect 27712 4276 27764 4282
rect 27712 4218 27764 4224
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 27908 2582 27936 8230
rect 28276 7886 28304 8774
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 28356 7744 28408 7750
rect 28356 7686 28408 7692
rect 28368 7546 28396 7686
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28552 7002 28580 13942
rect 28736 13870 28764 14282
rect 28828 14278 28856 16594
rect 29012 15638 29040 18119
rect 29104 17218 29132 22918
rect 29196 22012 29224 23072
rect 29288 22982 29316 32422
rect 29366 32328 29422 32337
rect 29366 32263 29368 32272
rect 29420 32263 29422 32272
rect 29368 32234 29420 32240
rect 29368 31748 29420 31754
rect 29368 31690 29420 31696
rect 29380 31346 29408 31690
rect 29368 31340 29420 31346
rect 29368 31282 29420 31288
rect 29368 31204 29420 31210
rect 29368 31146 29420 31152
rect 29380 30734 29408 31146
rect 29368 30728 29420 30734
rect 29368 30670 29420 30676
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29380 28218 29408 30194
rect 29472 29730 29500 37062
rect 29564 36242 29592 37266
rect 29552 36236 29604 36242
rect 29552 36178 29604 36184
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 29564 34746 29592 35974
rect 29552 34740 29604 34746
rect 29552 34682 29604 34688
rect 29552 34536 29604 34542
rect 29552 34478 29604 34484
rect 29564 31385 29592 34478
rect 29550 31376 29606 31385
rect 29550 31311 29606 31320
rect 29552 31272 29604 31278
rect 29552 31214 29604 31220
rect 29564 30666 29592 31214
rect 29552 30660 29604 30666
rect 29552 30602 29604 30608
rect 29550 30560 29606 30569
rect 29550 30495 29606 30504
rect 29564 30190 29592 30495
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 29564 29889 29592 30126
rect 29550 29880 29606 29889
rect 29550 29815 29606 29824
rect 29472 29702 29592 29730
rect 29460 29164 29512 29170
rect 29460 29106 29512 29112
rect 29472 29073 29500 29106
rect 29458 29064 29514 29073
rect 29458 28999 29514 29008
rect 29460 28960 29512 28966
rect 29460 28902 29512 28908
rect 29472 28218 29500 28902
rect 29368 28212 29420 28218
rect 29368 28154 29420 28160
rect 29460 28212 29512 28218
rect 29460 28154 29512 28160
rect 29366 28112 29422 28121
rect 29564 28098 29592 29702
rect 29656 28694 29684 39238
rect 29748 39030 29776 41126
rect 29920 41074 29972 41080
rect 29918 41032 29974 41041
rect 29918 40967 29974 40976
rect 29828 40928 29880 40934
rect 29828 40870 29880 40876
rect 29736 39024 29788 39030
rect 29736 38966 29788 38972
rect 29840 38962 29868 40870
rect 29932 40526 29960 40967
rect 29920 40520 29972 40526
rect 29920 40462 29972 40468
rect 30024 39964 30052 41375
rect 30116 41138 30144 41414
rect 30104 41132 30156 41138
rect 30104 41074 30156 41080
rect 30024 39936 30144 39964
rect 29920 39908 29972 39914
rect 29920 39850 29972 39856
rect 29828 38956 29880 38962
rect 29828 38898 29880 38904
rect 29932 38842 29960 39850
rect 30012 39840 30064 39846
rect 30012 39782 30064 39788
rect 30116 39794 30144 39936
rect 30208 39914 30236 53926
rect 30300 51270 30328 53994
rect 30288 51264 30340 51270
rect 30288 51206 30340 51212
rect 30288 48000 30340 48006
rect 30288 47942 30340 47948
rect 30300 41585 30328 47942
rect 30286 41576 30342 41585
rect 30286 41511 30342 41520
rect 30288 41472 30340 41478
rect 30288 41414 30340 41420
rect 30196 39908 30248 39914
rect 30196 39850 30248 39856
rect 29748 38814 29960 38842
rect 29748 32978 29776 38814
rect 29920 38752 29972 38758
rect 29920 38694 29972 38700
rect 29828 38480 29880 38486
rect 29828 38422 29880 38428
rect 29840 38010 29868 38422
rect 29828 38004 29880 38010
rect 29828 37946 29880 37952
rect 29828 37868 29880 37874
rect 29828 37810 29880 37816
rect 29840 37330 29868 37810
rect 29828 37324 29880 37330
rect 29828 37266 29880 37272
rect 29826 36816 29882 36825
rect 29826 36751 29828 36760
rect 29880 36751 29882 36760
rect 29828 36722 29880 36728
rect 29932 36553 29960 38694
rect 30024 37777 30052 39782
rect 30116 39766 30236 39794
rect 30104 39296 30156 39302
rect 30104 39238 30156 39244
rect 30010 37768 30066 37777
rect 30010 37703 30066 37712
rect 30116 37618 30144 39238
rect 30208 38350 30236 39766
rect 30196 38344 30248 38350
rect 30196 38286 30248 38292
rect 30196 38208 30248 38214
rect 30196 38150 30248 38156
rect 30024 37590 30144 37618
rect 30024 36825 30052 37590
rect 30104 37188 30156 37194
rect 30104 37130 30156 37136
rect 30010 36816 30066 36825
rect 30116 36786 30144 37130
rect 30010 36751 30066 36760
rect 30104 36780 30156 36786
rect 30104 36722 30156 36728
rect 30010 36680 30066 36689
rect 30010 36615 30066 36624
rect 30104 36644 30156 36650
rect 29918 36544 29974 36553
rect 29918 36479 29974 36488
rect 29932 36310 29960 36341
rect 29920 36304 29972 36310
rect 29918 36272 29920 36281
rect 29972 36272 29974 36281
rect 29918 36207 29974 36216
rect 29932 36174 29960 36207
rect 29920 36168 29972 36174
rect 29920 36110 29972 36116
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 29828 34400 29880 34406
rect 29828 34342 29880 34348
rect 29840 33998 29868 34342
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29828 33856 29880 33862
rect 29828 33798 29880 33804
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29736 32836 29788 32842
rect 29736 32778 29788 32784
rect 29748 31958 29776 32778
rect 29840 32586 29868 33798
rect 29932 32745 29960 35634
rect 30024 35086 30052 36615
rect 30104 36586 30156 36592
rect 30012 35080 30064 35086
rect 30012 35022 30064 35028
rect 30012 34944 30064 34950
rect 30012 34886 30064 34892
rect 30024 34105 30052 34886
rect 30116 34241 30144 36586
rect 30208 35873 30236 38150
rect 30194 35864 30250 35873
rect 30300 35834 30328 41414
rect 30392 38554 30420 54606
rect 30484 52193 30512 68274
rect 30564 65408 30616 65414
rect 30564 65350 30616 65356
rect 30576 63442 30604 65350
rect 30564 63436 30616 63442
rect 30564 63378 30616 63384
rect 30564 63300 30616 63306
rect 30564 63242 30616 63248
rect 30576 57050 30604 63242
rect 30668 61878 30696 69838
rect 30748 64864 30800 64870
rect 30748 64806 30800 64812
rect 30760 63918 30788 64806
rect 30748 63912 30800 63918
rect 30748 63854 30800 63860
rect 30656 61872 30708 61878
rect 30656 61814 30708 61820
rect 30748 59492 30800 59498
rect 30748 59434 30800 59440
rect 30656 59152 30708 59158
rect 30656 59094 30708 59100
rect 30668 58614 30696 59094
rect 30656 58608 30708 58614
rect 30656 58550 30708 58556
rect 30656 57248 30708 57254
rect 30654 57216 30656 57225
rect 30708 57216 30710 57225
rect 30654 57151 30710 57160
rect 30564 57044 30616 57050
rect 30564 56986 30616 56992
rect 30760 56234 30788 59434
rect 30748 56228 30800 56234
rect 30748 56170 30800 56176
rect 30748 55956 30800 55962
rect 30748 55898 30800 55904
rect 30564 55888 30616 55894
rect 30564 55830 30616 55836
rect 30470 52184 30526 52193
rect 30470 52119 30526 52128
rect 30472 52080 30524 52086
rect 30472 52022 30524 52028
rect 30484 51542 30512 52022
rect 30472 51536 30524 51542
rect 30472 51478 30524 51484
rect 30472 51264 30524 51270
rect 30472 51206 30524 51212
rect 30484 50969 30512 51206
rect 30470 50960 30526 50969
rect 30470 50895 30526 50904
rect 30470 50688 30526 50697
rect 30470 50623 30526 50632
rect 30484 42226 30512 50623
rect 30576 42265 30604 55830
rect 30656 55820 30708 55826
rect 30656 55762 30708 55768
rect 30668 44169 30696 55762
rect 30760 47122 30788 55898
rect 30852 55146 30880 71538
rect 31852 65680 31904 65686
rect 31852 65622 31904 65628
rect 31300 64660 31352 64666
rect 31300 64602 31352 64608
rect 31116 64456 31168 64462
rect 31116 64398 31168 64404
rect 30932 60648 30984 60654
rect 30932 60590 30984 60596
rect 30944 55690 30972 60590
rect 31024 59696 31076 59702
rect 31024 59638 31076 59644
rect 30932 55684 30984 55690
rect 30932 55626 30984 55632
rect 30932 55344 30984 55350
rect 30932 55286 30984 55292
rect 30840 55140 30892 55146
rect 30840 55082 30892 55088
rect 30944 55049 30972 55286
rect 30930 55040 30986 55049
rect 30930 54975 30986 54984
rect 30932 54732 30984 54738
rect 30932 54674 30984 54680
rect 30944 53666 30972 54674
rect 31036 53786 31064 59638
rect 31024 53780 31076 53786
rect 31024 53722 31076 53728
rect 30944 53638 31064 53666
rect 30932 53032 30984 53038
rect 30932 52974 30984 52980
rect 30840 52624 30892 52630
rect 30840 52566 30892 52572
rect 30852 51066 30880 52566
rect 30944 51241 30972 52974
rect 30930 51232 30986 51241
rect 30930 51167 30986 51176
rect 30840 51060 30892 51066
rect 30840 51002 30892 51008
rect 30930 50960 30986 50969
rect 30852 50918 30930 50946
rect 30748 47116 30800 47122
rect 30748 47058 30800 47064
rect 30748 46980 30800 46986
rect 30748 46922 30800 46928
rect 30654 44160 30710 44169
rect 30654 44095 30710 44104
rect 30654 43344 30710 43353
rect 30654 43279 30710 43288
rect 30668 42294 30696 43279
rect 30656 42288 30708 42294
rect 30562 42256 30618 42265
rect 30472 42220 30524 42226
rect 30656 42230 30708 42236
rect 30562 42191 30618 42200
rect 30472 42162 30524 42168
rect 30760 42140 30788 46922
rect 30668 42112 30788 42140
rect 30564 41812 30616 41818
rect 30564 41754 30616 41760
rect 30472 41472 30524 41478
rect 30472 41414 30524 41420
rect 30380 38548 30432 38554
rect 30380 38490 30432 38496
rect 30380 38344 30432 38350
rect 30380 38286 30432 38292
rect 30194 35799 30250 35808
rect 30288 35828 30340 35834
rect 30288 35770 30340 35776
rect 30392 35714 30420 38286
rect 30208 35686 30420 35714
rect 30102 34232 30158 34241
rect 30102 34167 30158 34176
rect 30010 34096 30066 34105
rect 30208 34082 30236 35686
rect 30288 35624 30340 35630
rect 30288 35566 30340 35572
rect 30010 34031 30066 34040
rect 30116 34054 30236 34082
rect 30012 33856 30064 33862
rect 30012 33798 30064 33804
rect 29918 32736 29974 32745
rect 29918 32671 29974 32680
rect 30024 32609 30052 33798
rect 30010 32600 30066 32609
rect 29840 32558 29960 32586
rect 29932 32450 29960 32558
rect 30010 32535 30066 32544
rect 29932 32422 30052 32450
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 29736 31952 29788 31958
rect 29736 31894 29788 31900
rect 29734 31784 29790 31793
rect 29734 31719 29790 31728
rect 29644 28688 29696 28694
rect 29644 28630 29696 28636
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 29366 28047 29422 28056
rect 29472 28070 29592 28098
rect 29380 28014 29408 28047
rect 29368 28008 29420 28014
rect 29368 27950 29420 27956
rect 29472 27606 29500 28070
rect 29552 28008 29604 28014
rect 29552 27950 29604 27956
rect 29460 27600 29512 27606
rect 29460 27542 29512 27548
rect 29368 27396 29420 27402
rect 29368 27338 29420 27344
rect 29380 25838 29408 27338
rect 29460 27124 29512 27130
rect 29460 27066 29512 27072
rect 29472 26994 29500 27066
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 29472 26586 29500 26726
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 29460 25968 29512 25974
rect 29460 25910 29512 25916
rect 29368 25832 29420 25838
rect 29368 25774 29420 25780
rect 29368 25424 29420 25430
rect 29368 25366 29420 25372
rect 29380 23322 29408 25366
rect 29472 24818 29500 25910
rect 29460 24812 29512 24818
rect 29460 24754 29512 24760
rect 29460 24608 29512 24614
rect 29460 24550 29512 24556
rect 29472 24342 29500 24550
rect 29460 24336 29512 24342
rect 29460 24278 29512 24284
rect 29368 23316 29420 23322
rect 29368 23258 29420 23264
rect 29368 23180 29420 23186
rect 29368 23122 29420 23128
rect 29276 22976 29328 22982
rect 29276 22918 29328 22924
rect 29380 22710 29408 23122
rect 29368 22704 29420 22710
rect 29368 22646 29420 22652
rect 29380 22030 29408 22646
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29368 22024 29420 22030
rect 29196 21984 29316 22012
rect 29184 21888 29236 21894
rect 29288 21876 29316 21984
rect 29368 21966 29420 21972
rect 29288 21848 29408 21876
rect 29184 21830 29236 21836
rect 29196 21146 29224 21830
rect 29276 21548 29328 21554
rect 29276 21490 29328 21496
rect 29184 21140 29236 21146
rect 29184 21082 29236 21088
rect 29184 20868 29236 20874
rect 29184 20810 29236 20816
rect 29196 20466 29224 20810
rect 29184 20460 29236 20466
rect 29184 20402 29236 20408
rect 29196 19802 29224 20402
rect 29288 19961 29316 21490
rect 29380 21486 29408 21848
rect 29368 21480 29420 21486
rect 29368 21422 29420 21428
rect 29472 20074 29500 22578
rect 29380 20046 29500 20074
rect 29274 19952 29330 19961
rect 29274 19887 29330 19896
rect 29196 19774 29316 19802
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 29196 19514 29224 19654
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29196 17338 29224 19314
rect 29288 17814 29316 19774
rect 29380 18358 29408 20046
rect 29460 19984 29512 19990
rect 29460 19926 29512 19932
rect 29472 19242 29500 19926
rect 29460 19236 29512 19242
rect 29460 19178 29512 19184
rect 29564 18970 29592 27950
rect 29656 22137 29684 28494
rect 29642 22128 29698 22137
rect 29642 22063 29698 22072
rect 29644 21956 29696 21962
rect 29644 21898 29696 21904
rect 29656 19378 29684 21898
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29368 18352 29420 18358
rect 29368 18294 29420 18300
rect 29380 18086 29408 18294
rect 29368 18080 29420 18086
rect 29368 18022 29420 18028
rect 29276 17808 29328 17814
rect 29276 17750 29328 17756
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 29104 17190 29684 17218
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29000 15632 29052 15638
rect 29000 15574 29052 15580
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 28908 14952 28960 14958
rect 28908 14894 28960 14900
rect 28816 14272 28868 14278
rect 28920 14249 28948 14894
rect 28816 14214 28868 14220
rect 28906 14240 28962 14249
rect 28906 14175 28962 14184
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28908 13864 28960 13870
rect 28908 13806 28960 13812
rect 28736 13530 28764 13806
rect 28724 13524 28776 13530
rect 28724 13466 28776 13472
rect 28736 13394 28764 13466
rect 28724 13388 28776 13394
rect 28724 13330 28776 13336
rect 28736 12918 28764 13330
rect 28724 12912 28776 12918
rect 28724 12854 28776 12860
rect 28814 12880 28870 12889
rect 28814 12815 28870 12824
rect 28828 11762 28856 12815
rect 28920 12345 28948 13806
rect 29012 13297 29040 15438
rect 28998 13288 29054 13297
rect 28998 13223 29054 13232
rect 28906 12336 28962 12345
rect 28906 12271 28962 12280
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28736 9625 28764 11086
rect 28816 9920 28868 9926
rect 28816 9862 28868 9868
rect 28722 9616 28778 9625
rect 28632 9580 28684 9586
rect 28722 9551 28778 9560
rect 28632 9522 28684 9528
rect 28644 8974 28672 9522
rect 28724 9104 28776 9110
rect 28724 9046 28776 9052
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28736 7886 28764 9046
rect 28828 9042 28856 9862
rect 28920 9081 28948 11086
rect 29196 10606 29224 17070
rect 29368 12776 29420 12782
rect 29368 12718 29420 12724
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29276 11688 29328 11694
rect 29276 11630 29328 11636
rect 29288 10985 29316 11630
rect 29380 11529 29408 12718
rect 29564 12434 29592 12718
rect 29472 12406 29592 12434
rect 29472 11762 29500 12406
rect 29656 12170 29684 17190
rect 29644 12164 29696 12170
rect 29644 12106 29696 12112
rect 29748 11830 29776 31719
rect 29840 22778 29868 32302
rect 30024 31754 30052 32422
rect 30116 31929 30144 34054
rect 30196 32768 30248 32774
rect 30196 32710 30248 32716
rect 30102 31920 30158 31929
rect 30102 31855 30158 31864
rect 30104 31816 30156 31822
rect 30104 31758 30156 31764
rect 29932 31726 30052 31754
rect 29932 26586 29960 31726
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 30024 31414 30052 31622
rect 30012 31408 30064 31414
rect 30012 31350 30064 31356
rect 30012 31272 30064 31278
rect 30012 31214 30064 31220
rect 30024 30394 30052 31214
rect 30116 30938 30144 31758
rect 30208 31686 30236 32710
rect 30196 31680 30248 31686
rect 30196 31622 30248 31628
rect 30300 31226 30328 35566
rect 30380 35080 30432 35086
rect 30380 35022 30432 35028
rect 30392 32026 30420 35022
rect 30380 32020 30432 32026
rect 30380 31962 30432 31968
rect 30380 31884 30432 31890
rect 30380 31826 30432 31832
rect 30208 31198 30328 31226
rect 30104 30932 30156 30938
rect 30104 30874 30156 30880
rect 30102 30696 30158 30705
rect 30102 30631 30158 30640
rect 30012 30388 30064 30394
rect 30012 30330 30064 30336
rect 30010 30288 30066 30297
rect 30010 30223 30066 30232
rect 30024 29850 30052 30223
rect 30012 29844 30064 29850
rect 30012 29786 30064 29792
rect 30116 29306 30144 30631
rect 30104 29300 30156 29306
rect 30104 29242 30156 29248
rect 30012 29164 30064 29170
rect 30012 29106 30064 29112
rect 30024 28801 30052 29106
rect 30010 28792 30066 28801
rect 30010 28727 30066 28736
rect 30104 28688 30156 28694
rect 30104 28630 30156 28636
rect 30012 28416 30064 28422
rect 30012 28358 30064 28364
rect 30024 27033 30052 28358
rect 30010 27024 30066 27033
rect 30010 26959 30066 26968
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 29920 26580 29972 26586
rect 29920 26522 29972 26528
rect 30024 25974 30052 26862
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 30010 25528 30066 25537
rect 30010 25463 30012 25472
rect 30064 25463 30066 25472
rect 30012 25434 30064 25440
rect 30116 25378 30144 28630
rect 30024 25350 30144 25378
rect 29920 24132 29972 24138
rect 29920 24074 29972 24080
rect 29932 22817 29960 24074
rect 29918 22808 29974 22817
rect 29828 22772 29880 22778
rect 29918 22743 29974 22752
rect 29828 22714 29880 22720
rect 30024 22094 30052 25350
rect 30102 24848 30158 24857
rect 30102 24783 30158 24792
rect 30116 22250 30144 24783
rect 30208 22386 30236 31198
rect 30286 31104 30342 31113
rect 30286 31039 30342 31048
rect 30300 22545 30328 31039
rect 30392 30841 30420 31826
rect 30378 30832 30434 30841
rect 30378 30767 30434 30776
rect 30380 30660 30432 30666
rect 30380 30602 30432 30608
rect 30392 26858 30420 30602
rect 30380 26852 30432 26858
rect 30380 26794 30432 26800
rect 30380 26376 30432 26382
rect 30380 26318 30432 26324
rect 30392 24750 30420 26318
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 30286 22536 30342 22545
rect 30286 22471 30342 22480
rect 30208 22358 30328 22386
rect 30116 22222 30236 22250
rect 29840 22066 30052 22094
rect 30102 22128 30158 22137
rect 29840 19990 29868 22066
rect 30102 22063 30158 22072
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29932 21622 29960 21966
rect 30012 21956 30064 21962
rect 30012 21898 30064 21904
rect 29920 21616 29972 21622
rect 29920 21558 29972 21564
rect 29932 20942 29960 21558
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 30024 20482 30052 21898
rect 30116 21146 30144 22063
rect 30208 21690 30236 22222
rect 30300 22098 30328 22358
rect 30288 22092 30340 22098
rect 30288 22034 30340 22040
rect 30196 21684 30248 21690
rect 30196 21626 30248 21632
rect 30196 21480 30248 21486
rect 30196 21422 30248 21428
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30208 21026 30236 21422
rect 29932 20454 30052 20482
rect 30116 20998 30236 21026
rect 29828 19984 29880 19990
rect 29828 19926 29880 19932
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29840 18465 29868 19790
rect 29826 18456 29882 18465
rect 29826 18391 29882 18400
rect 29932 18154 29960 20454
rect 30012 20392 30064 20398
rect 30012 20334 30064 20340
rect 30024 19446 30052 20334
rect 30012 19440 30064 19446
rect 30012 19382 30064 19388
rect 30010 19000 30066 19009
rect 30010 18935 30066 18944
rect 29920 18148 29972 18154
rect 29920 18090 29972 18096
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29918 18048 29974 18057
rect 29840 16454 29868 18022
rect 29918 17983 29974 17992
rect 29932 17678 29960 17983
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 30024 17270 30052 18935
rect 30012 17264 30064 17270
rect 30012 17206 30064 17212
rect 30116 17134 30144 20998
rect 30288 20052 30340 20058
rect 30288 19994 30340 20000
rect 30196 19984 30248 19990
rect 30196 19926 30248 19932
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 30104 16584 30156 16590
rect 30104 16526 30156 16532
rect 29828 16448 29880 16454
rect 29828 16390 29880 16396
rect 30116 16153 30144 16526
rect 30102 16144 30158 16153
rect 29920 16108 29972 16114
rect 30102 16079 30158 16088
rect 29920 16050 29972 16056
rect 29932 15745 29960 16050
rect 30208 15960 30236 19926
rect 30300 19334 30328 19994
rect 30392 19786 30420 24686
rect 30380 19780 30432 19786
rect 30380 19722 30432 19728
rect 30300 19306 30420 19334
rect 30288 18148 30340 18154
rect 30288 18090 30340 18096
rect 30024 15932 30236 15960
rect 29918 15736 29974 15745
rect 29918 15671 29974 15680
rect 29920 15428 29972 15434
rect 29920 15370 29972 15376
rect 29932 15201 29960 15370
rect 29918 15192 29974 15201
rect 29918 15127 29974 15136
rect 29826 14784 29882 14793
rect 29826 14719 29882 14728
rect 29840 14414 29868 14719
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 30024 13326 30052 15932
rect 30300 15858 30328 18090
rect 30116 15830 30328 15858
rect 30116 14482 30144 15830
rect 30392 14498 30420 19306
rect 30104 14476 30156 14482
rect 30104 14418 30156 14424
rect 30208 14470 30420 14498
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 29736 11824 29788 11830
rect 29736 11766 29788 11772
rect 29460 11756 29512 11762
rect 29460 11698 29512 11704
rect 29366 11520 29422 11529
rect 29366 11455 29422 11464
rect 29274 10976 29330 10985
rect 29274 10911 29330 10920
rect 29368 10804 29420 10810
rect 29368 10746 29420 10752
rect 29184 10600 29236 10606
rect 29184 10542 29236 10548
rect 29196 9518 29224 10542
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 28906 9072 28962 9081
rect 28816 9036 28868 9042
rect 28906 9007 28962 9016
rect 28816 8978 28868 8984
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 28828 7698 28856 8978
rect 28906 8664 28962 8673
rect 28906 8599 28962 8608
rect 28736 7670 28856 7698
rect 28540 6996 28592 7002
rect 28540 6938 28592 6944
rect 28736 6866 28764 7670
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28080 6656 28132 6662
rect 28080 6598 28132 6604
rect 28092 6390 28120 6598
rect 28080 6384 28132 6390
rect 28080 6326 28132 6332
rect 28736 6254 28764 6802
rect 28920 6798 28948 8599
rect 29196 8430 29224 9454
rect 29380 8838 29408 10746
rect 29932 10577 29960 12106
rect 29918 10568 29974 10577
rect 29918 10503 29974 10512
rect 29734 10024 29790 10033
rect 29734 9959 29736 9968
rect 29788 9959 29790 9968
rect 29736 9930 29788 9936
rect 30024 9178 30052 13262
rect 30116 11354 30144 14418
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 30012 9172 30064 9178
rect 30012 9114 30064 9120
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29368 8832 29420 8838
rect 29368 8774 29420 8780
rect 29368 8628 29420 8634
rect 29368 8570 29420 8576
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 28908 6792 28960 6798
rect 28814 6760 28870 6769
rect 28908 6734 28960 6740
rect 29012 6730 29040 7346
rect 28814 6695 28870 6704
rect 29000 6724 29052 6730
rect 28724 6248 28776 6254
rect 28724 6190 28776 6196
rect 27988 6112 28040 6118
rect 27988 6054 28040 6060
rect 28000 5710 28028 6054
rect 28828 5710 28856 6695
rect 29000 6666 29052 6672
rect 29012 5914 29040 6666
rect 29104 6662 29132 7482
rect 29196 7342 29224 8366
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29092 6656 29144 6662
rect 29092 6598 29144 6604
rect 29288 6458 29316 8434
rect 29276 6452 29328 6458
rect 29276 6394 29328 6400
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29000 5908 29052 5914
rect 29000 5850 29052 5856
rect 27988 5704 28040 5710
rect 27988 5646 28040 5652
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 29104 5370 29132 6258
rect 29288 5914 29316 6394
rect 29380 6390 29408 8570
rect 29840 8129 29868 8910
rect 29826 8120 29882 8129
rect 29826 8055 29882 8064
rect 30208 6866 30236 14470
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30392 8906 30420 9590
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30484 7546 30512 41414
rect 30576 36310 30604 41754
rect 30668 41478 30696 42112
rect 30746 41712 30802 41721
rect 30746 41647 30802 41656
rect 30656 41472 30708 41478
rect 30656 41414 30708 41420
rect 30654 40760 30710 40769
rect 30654 40695 30710 40704
rect 30564 36304 30616 36310
rect 30564 36246 30616 36252
rect 30668 36156 30696 40695
rect 30576 36128 30696 36156
rect 30576 32842 30604 36128
rect 30760 36088 30788 41647
rect 30852 41585 30880 50918
rect 30930 50895 30986 50904
rect 30932 50856 30984 50862
rect 30932 50798 30984 50804
rect 30944 50561 30972 50798
rect 30930 50552 30986 50561
rect 30930 50487 30986 50496
rect 30932 49972 30984 49978
rect 30932 49914 30984 49920
rect 30944 49337 30972 49914
rect 30930 49328 30986 49337
rect 30930 49263 30986 49272
rect 30932 49156 30984 49162
rect 30932 49098 30984 49104
rect 30944 47297 30972 49098
rect 30930 47288 30986 47297
rect 30930 47223 30986 47232
rect 30932 47116 30984 47122
rect 30932 47058 30984 47064
rect 30944 46306 30972 47058
rect 30932 46300 30984 46306
rect 30932 46242 30984 46248
rect 31036 46186 31064 53638
rect 31128 48278 31156 64398
rect 31208 58608 31260 58614
rect 31208 58550 31260 58556
rect 31220 55706 31248 58550
rect 31312 55894 31340 64602
rect 31668 63912 31720 63918
rect 31390 63880 31446 63889
rect 31668 63854 31720 63860
rect 31390 63815 31446 63824
rect 31404 55962 31432 63815
rect 31484 58472 31536 58478
rect 31484 58414 31536 58420
rect 31392 55956 31444 55962
rect 31392 55898 31444 55904
rect 31300 55888 31352 55894
rect 31300 55830 31352 55836
rect 31220 55678 31340 55706
rect 31208 54868 31260 54874
rect 31208 54810 31260 54816
rect 31116 48272 31168 48278
rect 31116 48214 31168 48220
rect 31116 48136 31168 48142
rect 31116 48078 31168 48084
rect 31128 46481 31156 48078
rect 31114 46472 31170 46481
rect 31114 46407 31170 46416
rect 31116 46368 31168 46374
rect 31116 46310 31168 46316
rect 30944 46158 31064 46186
rect 30838 41576 30894 41585
rect 30838 41511 30894 41520
rect 30840 41472 30892 41478
rect 30840 41414 30892 41420
rect 30668 36060 30788 36088
rect 30564 32836 30616 32842
rect 30564 32778 30616 32784
rect 30668 32178 30696 36060
rect 30852 35986 30880 41414
rect 30576 32150 30696 32178
rect 30760 35958 30880 35986
rect 30576 31754 30604 32150
rect 30576 31726 30696 31754
rect 30564 31680 30616 31686
rect 30564 31622 30616 31628
rect 30576 31249 30604 31622
rect 30562 31240 30618 31249
rect 30562 31175 30618 31184
rect 30562 30968 30618 30977
rect 30562 30903 30618 30912
rect 30576 26926 30604 30903
rect 30564 26920 30616 26926
rect 30564 26862 30616 26868
rect 30564 25764 30616 25770
rect 30564 25706 30616 25712
rect 30576 21894 30604 25706
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30668 10810 30696 31726
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30760 8634 30788 35958
rect 30840 35828 30892 35834
rect 30840 35770 30892 35776
rect 30852 34746 30880 35770
rect 30840 34740 30892 34746
rect 30840 34682 30892 34688
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30852 32065 30880 33254
rect 30838 32056 30894 32065
rect 30838 31991 30894 32000
rect 30840 31952 30892 31958
rect 30840 31894 30892 31900
rect 30852 27130 30880 31894
rect 30944 27316 30972 46158
rect 31024 46096 31076 46102
rect 31024 46038 31076 46044
rect 31036 27470 31064 46038
rect 31128 41546 31156 46310
rect 31116 41540 31168 41546
rect 31116 41482 31168 41488
rect 31116 41404 31168 41410
rect 31116 41346 31168 41352
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 30944 27288 31064 27316
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30852 14618 30880 25230
rect 30944 17746 30972 26862
rect 31036 18222 31064 27288
rect 31024 18216 31076 18222
rect 31024 18158 31076 18164
rect 30932 17740 30984 17746
rect 30932 17682 30984 17688
rect 31128 16250 31156 41346
rect 31220 19514 31248 54810
rect 31312 54670 31340 55678
rect 31300 54664 31352 54670
rect 31300 54606 31352 54612
rect 31300 54528 31352 54534
rect 31300 54470 31352 54476
rect 31312 51241 31340 54470
rect 31392 54120 31444 54126
rect 31392 54062 31444 54068
rect 31298 51232 31354 51241
rect 31298 51167 31354 51176
rect 31298 50280 31354 50289
rect 31298 50215 31354 50224
rect 31312 36650 31340 50215
rect 31404 46481 31432 54062
rect 31390 46472 31446 46481
rect 31390 46407 31446 46416
rect 31392 46300 31444 46306
rect 31392 46242 31444 46248
rect 31404 42362 31432 46242
rect 31392 42356 31444 42362
rect 31392 42298 31444 42304
rect 31392 41812 31444 41818
rect 31392 41754 31444 41760
rect 31404 37097 31432 41754
rect 31390 37088 31446 37097
rect 31390 37023 31446 37032
rect 31300 36644 31352 36650
rect 31300 36586 31352 36592
rect 31392 36304 31444 36310
rect 31392 36246 31444 36252
rect 31298 36136 31354 36145
rect 31298 36071 31354 36080
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 31312 16658 31340 36071
rect 31404 29102 31432 36246
rect 31496 31074 31524 58414
rect 31576 56228 31628 56234
rect 31576 56170 31628 56176
rect 31484 31068 31536 31074
rect 31484 31010 31536 31016
rect 31482 30968 31538 30977
rect 31482 30903 31538 30912
rect 31392 29096 31444 29102
rect 31392 29038 31444 29044
rect 31496 27878 31524 30903
rect 31484 27872 31536 27878
rect 31484 27814 31536 27820
rect 31484 27600 31536 27606
rect 31484 27542 31536 27548
rect 31392 26512 31444 26518
rect 31392 26454 31444 26460
rect 31300 16652 31352 16658
rect 31300 16594 31352 16600
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 30840 14612 30892 14618
rect 30840 14554 30892 14560
rect 31404 13462 31432 26454
rect 31496 22574 31524 27542
rect 31484 22568 31536 22574
rect 31484 22510 31536 22516
rect 31588 20602 31616 56170
rect 31680 55826 31708 63854
rect 31864 57974 31892 65622
rect 31772 57946 31892 57974
rect 31772 56896 31800 57946
rect 31772 56868 31892 56896
rect 31668 55820 31720 55826
rect 31668 55762 31720 55768
rect 31760 55684 31812 55690
rect 31760 55626 31812 55632
rect 31668 55208 31720 55214
rect 31668 55150 31720 55156
rect 31680 52902 31708 55150
rect 31668 52896 31720 52902
rect 31668 52838 31720 52844
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 31576 19100 31628 19106
rect 31576 19042 31628 19048
rect 31588 14498 31616 19042
rect 31680 18426 31708 52838
rect 31772 46170 31800 55626
rect 31864 50980 31892 56868
rect 31864 50952 31984 50980
rect 31852 50856 31904 50862
rect 31852 50798 31904 50804
rect 31760 46164 31812 46170
rect 31760 46106 31812 46112
rect 31864 46102 31892 50798
rect 31852 46096 31904 46102
rect 31852 46038 31904 46044
rect 31956 45778 31984 50952
rect 31864 45762 31984 45778
rect 31852 45756 31984 45762
rect 31904 45750 31984 45756
rect 31852 45698 31904 45704
rect 31760 45280 31812 45286
rect 31760 45222 31812 45228
rect 31772 31929 31800 45222
rect 31864 45206 31984 45234
rect 31864 45121 31892 45206
rect 31850 45112 31906 45121
rect 31850 45047 31906 45056
rect 31852 45008 31904 45014
rect 31852 44950 31904 44956
rect 31864 41274 31892 44950
rect 31852 41268 31904 41274
rect 31852 41210 31904 41216
rect 31850 38040 31906 38049
rect 31850 37975 31906 37984
rect 31758 31920 31814 31929
rect 31758 31855 31814 31864
rect 31760 30660 31812 30666
rect 31760 30602 31812 30608
rect 31772 27606 31800 30602
rect 31760 27600 31812 27606
rect 31760 27542 31812 27548
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31772 19922 31800 27406
rect 31760 19916 31812 19922
rect 31760 19858 31812 19864
rect 31864 19334 31892 37975
rect 31772 19306 31892 19334
rect 31772 19106 31800 19306
rect 31760 19100 31812 19106
rect 31760 19042 31812 19048
rect 31956 18816 31984 45206
rect 31772 18788 31984 18816
rect 31772 18630 31800 18788
rect 31760 18624 31812 18630
rect 31760 18566 31812 18572
rect 31668 18420 31720 18426
rect 31668 18362 31720 18368
rect 31588 14470 31892 14498
rect 31392 13456 31444 13462
rect 31392 13398 31444 13404
rect 31864 9654 31892 14470
rect 31852 9648 31904 9654
rect 31852 9590 31904 9596
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 29826 6488 29882 6497
rect 29826 6423 29828 6432
rect 29880 6423 29882 6432
rect 29828 6394 29880 6400
rect 29368 6384 29420 6390
rect 29368 6326 29420 6332
rect 30102 6216 30158 6225
rect 30102 6151 30158 6160
rect 29368 6112 29420 6118
rect 29368 6054 29420 6060
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 29380 5302 29408 6054
rect 30116 5710 30144 6151
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 29826 5400 29882 5409
rect 29826 5335 29828 5344
rect 29880 5335 29882 5344
rect 29828 5306 29880 5312
rect 29368 5296 29420 5302
rect 29368 5238 29420 5244
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 29092 5228 29144 5234
rect 29092 5170 29144 5176
rect 28184 4865 28212 5170
rect 28170 4856 28226 4865
rect 28170 4791 28226 4800
rect 28722 4720 28778 4729
rect 29012 4690 29040 5170
rect 28722 4655 28724 4664
rect 28776 4655 28778 4664
rect 29000 4684 29052 4690
rect 28724 4626 28776 4632
rect 29000 4626 29052 4632
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28184 3913 28212 4082
rect 29104 4010 29132 5170
rect 29920 5160 29972 5166
rect 29920 5102 29972 5108
rect 29368 5024 29420 5030
rect 29368 4966 29420 4972
rect 29092 4004 29144 4010
rect 29092 3946 29144 3952
rect 28632 3936 28684 3942
rect 28170 3904 28226 3913
rect 28632 3878 28684 3884
rect 28170 3839 28226 3848
rect 28644 3738 28672 3878
rect 28632 3732 28684 3738
rect 28632 3674 28684 3680
rect 29380 3534 29408 4966
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29748 3670 29776 4082
rect 29932 4078 29960 5102
rect 29828 4072 29880 4078
rect 29826 4040 29828 4049
rect 29920 4072 29972 4078
rect 29880 4040 29882 4049
rect 29920 4014 29972 4020
rect 29826 3975 29882 3984
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 28264 3528 28316 3534
rect 28262 3496 28264 3505
rect 29368 3528 29420 3534
rect 28316 3496 28318 3505
rect 29368 3470 29420 3476
rect 28262 3431 28318 3440
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 27896 2576 27948 2582
rect 27896 2518 27948 2524
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 25044 2372 25096 2378
rect 25044 2314 25096 2320
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 2870 368 2926 377
rect 2870 303 2926 312
rect 28276 241 28304 2382
rect 28736 2009 28764 2382
rect 28722 2000 28778 2009
rect 28722 1935 28778 1944
rect 28828 1601 28856 2994
rect 28920 2961 28948 3334
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 28906 2952 28962 2961
rect 28906 2887 28962 2896
rect 29748 2553 29776 2994
rect 29734 2544 29790 2553
rect 29734 2479 29790 2488
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28814 1592 28870 1601
rect 28814 1527 28870 1536
rect 28724 1352 28776 1358
rect 28724 1294 28776 1300
rect 28736 649 28764 1294
rect 29656 1057 29684 2382
rect 29642 1048 29698 1057
rect 29642 983 29698 992
rect 28722 640 28778 649
rect 28722 575 28778 584
rect 28262 232 28318 241
rect 28262 167 28318 176
<< via2 >>
rect 3790 79600 3846 79656
rect 27894 79600 27950 79656
rect 2778 78920 2834 78976
rect 1306 78240 1362 78296
rect 1398 77580 1454 77616
rect 1398 77560 1400 77580
rect 1400 77560 1452 77580
rect 1452 77560 1454 77580
rect 5921 77818 5977 77820
rect 6001 77818 6057 77820
rect 6081 77818 6137 77820
rect 6161 77818 6217 77820
rect 5921 77766 5967 77818
rect 5967 77766 5977 77818
rect 6001 77766 6031 77818
rect 6031 77766 6043 77818
rect 6043 77766 6057 77818
rect 6081 77766 6095 77818
rect 6095 77766 6107 77818
rect 6107 77766 6137 77818
rect 6161 77766 6171 77818
rect 6171 77766 6217 77818
rect 5921 77764 5977 77766
rect 6001 77764 6057 77766
rect 6081 77764 6137 77766
rect 6161 77764 6217 77766
rect 15852 77818 15908 77820
rect 15932 77818 15988 77820
rect 16012 77818 16068 77820
rect 16092 77818 16148 77820
rect 15852 77766 15898 77818
rect 15898 77766 15908 77818
rect 15932 77766 15962 77818
rect 15962 77766 15974 77818
rect 15974 77766 15988 77818
rect 16012 77766 16026 77818
rect 16026 77766 16038 77818
rect 16038 77766 16068 77818
rect 16092 77766 16102 77818
rect 16102 77766 16148 77818
rect 15852 77764 15908 77766
rect 15932 77764 15988 77766
rect 16012 77764 16068 77766
rect 16092 77764 16148 77766
rect 25782 77818 25838 77820
rect 25862 77818 25918 77820
rect 25942 77818 25998 77820
rect 26022 77818 26078 77820
rect 25782 77766 25828 77818
rect 25828 77766 25838 77818
rect 25862 77766 25892 77818
rect 25892 77766 25904 77818
rect 25904 77766 25918 77818
rect 25942 77766 25956 77818
rect 25956 77766 25968 77818
rect 25968 77766 25998 77818
rect 26022 77766 26032 77818
rect 26032 77766 26078 77818
rect 25782 77764 25838 77766
rect 25862 77764 25918 77766
rect 25942 77764 25998 77766
rect 26022 77764 26078 77766
rect 28814 79192 28870 79248
rect 28538 78648 28594 78704
rect 28170 78240 28226 78296
rect 10886 77274 10942 77276
rect 10966 77274 11022 77276
rect 11046 77274 11102 77276
rect 11126 77274 11182 77276
rect 10886 77222 10932 77274
rect 10932 77222 10942 77274
rect 10966 77222 10996 77274
rect 10996 77222 11008 77274
rect 11008 77222 11022 77274
rect 11046 77222 11060 77274
rect 11060 77222 11072 77274
rect 11072 77222 11102 77274
rect 11126 77222 11136 77274
rect 11136 77222 11182 77274
rect 10886 77220 10942 77222
rect 10966 77220 11022 77222
rect 11046 77220 11102 77222
rect 11126 77220 11182 77222
rect 1398 76916 1400 76936
rect 1400 76916 1452 76936
rect 1452 76916 1454 76936
rect 1398 76880 1454 76916
rect 5921 76730 5977 76732
rect 6001 76730 6057 76732
rect 6081 76730 6137 76732
rect 6161 76730 6217 76732
rect 5921 76678 5967 76730
rect 5967 76678 5977 76730
rect 6001 76678 6031 76730
rect 6031 76678 6043 76730
rect 6043 76678 6057 76730
rect 6081 76678 6095 76730
rect 6095 76678 6107 76730
rect 6107 76678 6137 76730
rect 6161 76678 6171 76730
rect 6171 76678 6217 76730
rect 5921 76676 5977 76678
rect 6001 76676 6057 76678
rect 6081 76676 6137 76678
rect 6161 76676 6217 76678
rect 2870 76200 2926 76256
rect 5921 75642 5977 75644
rect 6001 75642 6057 75644
rect 6081 75642 6137 75644
rect 6161 75642 6217 75644
rect 5921 75590 5967 75642
rect 5967 75590 5977 75642
rect 6001 75590 6031 75642
rect 6031 75590 6043 75642
rect 6043 75590 6057 75642
rect 6081 75590 6095 75642
rect 6095 75590 6107 75642
rect 6107 75590 6137 75642
rect 6161 75590 6171 75642
rect 6171 75590 6217 75642
rect 5921 75588 5977 75590
rect 6001 75588 6057 75590
rect 6081 75588 6137 75590
rect 6161 75588 6217 75590
rect 1582 75520 1638 75576
rect 1582 74976 1638 75032
rect 5921 74554 5977 74556
rect 6001 74554 6057 74556
rect 6081 74554 6137 74556
rect 6161 74554 6217 74556
rect 5921 74502 5967 74554
rect 5967 74502 5977 74554
rect 6001 74502 6031 74554
rect 6031 74502 6043 74554
rect 6043 74502 6057 74554
rect 6081 74502 6095 74554
rect 6095 74502 6107 74554
rect 6107 74502 6137 74554
rect 6161 74502 6171 74554
rect 6171 74502 6217 74554
rect 5921 74500 5977 74502
rect 6001 74500 6057 74502
rect 6081 74500 6137 74502
rect 6161 74500 6217 74502
rect 1582 74296 1638 74352
rect 1582 73616 1638 73672
rect 5921 73466 5977 73468
rect 6001 73466 6057 73468
rect 6081 73466 6137 73468
rect 6161 73466 6217 73468
rect 5921 73414 5967 73466
rect 5967 73414 5977 73466
rect 6001 73414 6031 73466
rect 6031 73414 6043 73466
rect 6043 73414 6057 73466
rect 6081 73414 6095 73466
rect 6095 73414 6107 73466
rect 6107 73414 6137 73466
rect 6161 73414 6171 73466
rect 6171 73414 6217 73466
rect 5921 73412 5977 73414
rect 6001 73412 6057 73414
rect 6081 73412 6137 73414
rect 6161 73412 6217 73414
rect 1582 72936 1638 72992
rect 5921 72378 5977 72380
rect 6001 72378 6057 72380
rect 6081 72378 6137 72380
rect 6161 72378 6217 72380
rect 5921 72326 5967 72378
rect 5967 72326 5977 72378
rect 6001 72326 6031 72378
rect 6031 72326 6043 72378
rect 6043 72326 6057 72378
rect 6081 72326 6095 72378
rect 6095 72326 6107 72378
rect 6107 72326 6137 72378
rect 6161 72326 6171 72378
rect 6171 72326 6217 72378
rect 5921 72324 5977 72326
rect 6001 72324 6057 72326
rect 6081 72324 6137 72326
rect 6161 72324 6217 72326
rect 1582 72256 1638 72312
rect 1582 71576 1638 71632
rect 5921 71290 5977 71292
rect 6001 71290 6057 71292
rect 6081 71290 6137 71292
rect 6161 71290 6217 71292
rect 5921 71238 5967 71290
rect 5967 71238 5977 71290
rect 6001 71238 6031 71290
rect 6031 71238 6043 71290
rect 6043 71238 6057 71290
rect 6081 71238 6095 71290
rect 6095 71238 6107 71290
rect 6107 71238 6137 71290
rect 6161 71238 6171 71290
rect 6171 71238 6217 71290
rect 5921 71236 5977 71238
rect 6001 71236 6057 71238
rect 6081 71236 6137 71238
rect 6161 71236 6217 71238
rect 1398 70932 1400 70952
rect 1400 70932 1452 70952
rect 1452 70932 1454 70952
rect 1398 70896 1454 70932
rect 1582 70352 1638 70408
rect 5921 70202 5977 70204
rect 6001 70202 6057 70204
rect 6081 70202 6137 70204
rect 6161 70202 6217 70204
rect 5921 70150 5967 70202
rect 5967 70150 5977 70202
rect 6001 70150 6031 70202
rect 6031 70150 6043 70202
rect 6043 70150 6057 70202
rect 6081 70150 6095 70202
rect 6095 70150 6107 70202
rect 6107 70150 6137 70202
rect 6161 70150 6171 70202
rect 6171 70150 6217 70202
rect 5921 70148 5977 70150
rect 6001 70148 6057 70150
rect 6081 70148 6137 70150
rect 6161 70148 6217 70150
rect 10886 76186 10942 76188
rect 10966 76186 11022 76188
rect 11046 76186 11102 76188
rect 11126 76186 11182 76188
rect 10886 76134 10932 76186
rect 10932 76134 10942 76186
rect 10966 76134 10996 76186
rect 10996 76134 11008 76186
rect 11008 76134 11022 76186
rect 11046 76134 11060 76186
rect 11060 76134 11072 76186
rect 11072 76134 11102 76186
rect 11126 76134 11136 76186
rect 11136 76134 11182 76186
rect 10886 76132 10942 76134
rect 10966 76132 11022 76134
rect 11046 76132 11102 76134
rect 11126 76132 11182 76134
rect 10886 75098 10942 75100
rect 10966 75098 11022 75100
rect 11046 75098 11102 75100
rect 11126 75098 11182 75100
rect 10886 75046 10932 75098
rect 10932 75046 10942 75098
rect 10966 75046 10996 75098
rect 10996 75046 11008 75098
rect 11008 75046 11022 75098
rect 11046 75046 11060 75098
rect 11060 75046 11072 75098
rect 11072 75046 11102 75098
rect 11126 75046 11136 75098
rect 11136 75046 11182 75098
rect 10886 75044 10942 75046
rect 10966 75044 11022 75046
rect 11046 75044 11102 75046
rect 11126 75044 11182 75046
rect 10886 74010 10942 74012
rect 10966 74010 11022 74012
rect 11046 74010 11102 74012
rect 11126 74010 11182 74012
rect 10886 73958 10932 74010
rect 10932 73958 10942 74010
rect 10966 73958 10996 74010
rect 10996 73958 11008 74010
rect 11008 73958 11022 74010
rect 11046 73958 11060 74010
rect 11060 73958 11072 74010
rect 11072 73958 11102 74010
rect 11126 73958 11136 74010
rect 11136 73958 11182 74010
rect 10886 73956 10942 73958
rect 10966 73956 11022 73958
rect 11046 73956 11102 73958
rect 11126 73956 11182 73958
rect 10886 72922 10942 72924
rect 10966 72922 11022 72924
rect 11046 72922 11102 72924
rect 11126 72922 11182 72924
rect 10886 72870 10932 72922
rect 10932 72870 10942 72922
rect 10966 72870 10996 72922
rect 10996 72870 11008 72922
rect 11008 72870 11022 72922
rect 11046 72870 11060 72922
rect 11060 72870 11072 72922
rect 11072 72870 11102 72922
rect 11126 72870 11136 72922
rect 11136 72870 11182 72922
rect 10886 72868 10942 72870
rect 10966 72868 11022 72870
rect 11046 72868 11102 72870
rect 11126 72868 11182 72870
rect 10886 71834 10942 71836
rect 10966 71834 11022 71836
rect 11046 71834 11102 71836
rect 11126 71834 11182 71836
rect 10886 71782 10932 71834
rect 10932 71782 10942 71834
rect 10966 71782 10996 71834
rect 10996 71782 11008 71834
rect 11008 71782 11022 71834
rect 11046 71782 11060 71834
rect 11060 71782 11072 71834
rect 11072 71782 11102 71834
rect 11126 71782 11136 71834
rect 11136 71782 11182 71834
rect 10886 71780 10942 71782
rect 10966 71780 11022 71782
rect 11046 71780 11102 71782
rect 11126 71780 11182 71782
rect 10886 70746 10942 70748
rect 10966 70746 11022 70748
rect 11046 70746 11102 70748
rect 11126 70746 11182 70748
rect 10886 70694 10932 70746
rect 10932 70694 10942 70746
rect 10966 70694 10996 70746
rect 10996 70694 11008 70746
rect 11008 70694 11022 70746
rect 11046 70694 11060 70746
rect 11060 70694 11072 70746
rect 11072 70694 11102 70746
rect 11126 70694 11136 70746
rect 11136 70694 11182 70746
rect 10886 70692 10942 70694
rect 10966 70692 11022 70694
rect 11046 70692 11102 70694
rect 11126 70692 11182 70694
rect 20817 77274 20873 77276
rect 20897 77274 20953 77276
rect 20977 77274 21033 77276
rect 21057 77274 21113 77276
rect 20817 77222 20863 77274
rect 20863 77222 20873 77274
rect 20897 77222 20927 77274
rect 20927 77222 20939 77274
rect 20939 77222 20953 77274
rect 20977 77222 20991 77274
rect 20991 77222 21003 77274
rect 21003 77222 21033 77274
rect 21057 77222 21067 77274
rect 21067 77222 21113 77274
rect 20817 77220 20873 77222
rect 20897 77220 20953 77222
rect 20977 77220 21033 77222
rect 21057 77220 21113 77222
rect 15852 76730 15908 76732
rect 15932 76730 15988 76732
rect 16012 76730 16068 76732
rect 16092 76730 16148 76732
rect 15852 76678 15898 76730
rect 15898 76678 15908 76730
rect 15932 76678 15962 76730
rect 15962 76678 15974 76730
rect 15974 76678 15988 76730
rect 16012 76678 16026 76730
rect 16026 76678 16038 76730
rect 16038 76678 16068 76730
rect 16092 76678 16102 76730
rect 16102 76678 16148 76730
rect 15852 76676 15908 76678
rect 15932 76676 15988 76678
rect 16012 76676 16068 76678
rect 16092 76676 16148 76678
rect 25782 76730 25838 76732
rect 25862 76730 25918 76732
rect 25942 76730 25998 76732
rect 26022 76730 26078 76732
rect 25782 76678 25828 76730
rect 25828 76678 25838 76730
rect 25862 76678 25892 76730
rect 25892 76678 25904 76730
rect 25904 76678 25918 76730
rect 25942 76678 25956 76730
rect 25956 76678 25968 76730
rect 25968 76678 25998 76730
rect 26022 76678 26032 76730
rect 26032 76678 26078 76730
rect 25782 76676 25838 76678
rect 25862 76676 25918 76678
rect 25942 76676 25998 76678
rect 26022 76676 26078 76678
rect 20817 76186 20873 76188
rect 20897 76186 20953 76188
rect 20977 76186 21033 76188
rect 21057 76186 21113 76188
rect 20817 76134 20863 76186
rect 20863 76134 20873 76186
rect 20897 76134 20927 76186
rect 20927 76134 20939 76186
rect 20939 76134 20953 76186
rect 20977 76134 20991 76186
rect 20991 76134 21003 76186
rect 21003 76134 21033 76186
rect 21057 76134 21067 76186
rect 21067 76134 21113 76186
rect 20817 76132 20873 76134
rect 20897 76132 20953 76134
rect 20977 76132 21033 76134
rect 21057 76132 21113 76134
rect 15852 75642 15908 75644
rect 15932 75642 15988 75644
rect 16012 75642 16068 75644
rect 16092 75642 16148 75644
rect 15852 75590 15898 75642
rect 15898 75590 15908 75642
rect 15932 75590 15962 75642
rect 15962 75590 15974 75642
rect 15974 75590 15988 75642
rect 16012 75590 16026 75642
rect 16026 75590 16038 75642
rect 16038 75590 16068 75642
rect 16092 75590 16102 75642
rect 16102 75590 16148 75642
rect 15852 75588 15908 75590
rect 15932 75588 15988 75590
rect 16012 75588 16068 75590
rect 16092 75588 16148 75590
rect 15852 74554 15908 74556
rect 15932 74554 15988 74556
rect 16012 74554 16068 74556
rect 16092 74554 16148 74556
rect 15852 74502 15898 74554
rect 15898 74502 15908 74554
rect 15932 74502 15962 74554
rect 15962 74502 15974 74554
rect 15974 74502 15988 74554
rect 16012 74502 16026 74554
rect 16026 74502 16038 74554
rect 16038 74502 16068 74554
rect 16092 74502 16102 74554
rect 16102 74502 16148 74554
rect 15852 74500 15908 74502
rect 15932 74500 15988 74502
rect 16012 74500 16068 74502
rect 16092 74500 16148 74502
rect 15852 73466 15908 73468
rect 15932 73466 15988 73468
rect 16012 73466 16068 73468
rect 16092 73466 16148 73468
rect 15852 73414 15898 73466
rect 15898 73414 15908 73466
rect 15932 73414 15962 73466
rect 15962 73414 15974 73466
rect 15974 73414 15988 73466
rect 16012 73414 16026 73466
rect 16026 73414 16038 73466
rect 16038 73414 16068 73466
rect 16092 73414 16102 73466
rect 16102 73414 16148 73466
rect 15852 73412 15908 73414
rect 15932 73412 15988 73414
rect 16012 73412 16068 73414
rect 16092 73412 16148 73414
rect 15842 73108 15844 73128
rect 15844 73108 15896 73128
rect 15896 73108 15898 73128
rect 15842 73072 15898 73108
rect 15852 72378 15908 72380
rect 15932 72378 15988 72380
rect 16012 72378 16068 72380
rect 16092 72378 16148 72380
rect 15852 72326 15898 72378
rect 15898 72326 15908 72378
rect 15932 72326 15962 72378
rect 15962 72326 15974 72378
rect 15974 72326 15988 72378
rect 16012 72326 16026 72378
rect 16026 72326 16038 72378
rect 16038 72326 16068 72378
rect 16092 72326 16102 72378
rect 16102 72326 16148 72378
rect 15852 72324 15908 72326
rect 15932 72324 15988 72326
rect 16012 72324 16068 72326
rect 16092 72324 16148 72326
rect 15852 71290 15908 71292
rect 15932 71290 15988 71292
rect 16012 71290 16068 71292
rect 16092 71290 16148 71292
rect 15852 71238 15898 71290
rect 15898 71238 15908 71290
rect 15932 71238 15962 71290
rect 15962 71238 15974 71290
rect 15974 71238 15988 71290
rect 16012 71238 16026 71290
rect 16026 71238 16038 71290
rect 16038 71238 16068 71290
rect 16092 71238 16102 71290
rect 16102 71238 16148 71290
rect 15852 71236 15908 71238
rect 15932 71236 15988 71238
rect 16012 71236 16068 71238
rect 16092 71236 16148 71238
rect 1582 69672 1638 69728
rect 10886 69658 10942 69660
rect 10966 69658 11022 69660
rect 11046 69658 11102 69660
rect 11126 69658 11182 69660
rect 10886 69606 10932 69658
rect 10932 69606 10942 69658
rect 10966 69606 10996 69658
rect 10996 69606 11008 69658
rect 11008 69606 11022 69658
rect 11046 69606 11060 69658
rect 11060 69606 11072 69658
rect 11072 69606 11102 69658
rect 11126 69606 11136 69658
rect 11136 69606 11182 69658
rect 10886 69604 10942 69606
rect 10966 69604 11022 69606
rect 11046 69604 11102 69606
rect 11126 69604 11182 69606
rect 5921 69114 5977 69116
rect 6001 69114 6057 69116
rect 6081 69114 6137 69116
rect 6161 69114 6217 69116
rect 5921 69062 5967 69114
rect 5967 69062 5977 69114
rect 6001 69062 6031 69114
rect 6031 69062 6043 69114
rect 6043 69062 6057 69114
rect 6081 69062 6095 69114
rect 6095 69062 6107 69114
rect 6107 69062 6137 69114
rect 6161 69062 6171 69114
rect 6171 69062 6217 69114
rect 5921 69060 5977 69062
rect 6001 69060 6057 69062
rect 6081 69060 6137 69062
rect 6161 69060 6217 69062
rect 1582 68992 1638 69048
rect 10886 68570 10942 68572
rect 10966 68570 11022 68572
rect 11046 68570 11102 68572
rect 11126 68570 11182 68572
rect 10886 68518 10932 68570
rect 10932 68518 10942 68570
rect 10966 68518 10996 68570
rect 10996 68518 11008 68570
rect 11008 68518 11022 68570
rect 11046 68518 11060 68570
rect 11060 68518 11072 68570
rect 11072 68518 11102 68570
rect 11126 68518 11136 68570
rect 11136 68518 11182 68570
rect 10886 68516 10942 68518
rect 10966 68516 11022 68518
rect 11046 68516 11102 68518
rect 11126 68516 11182 68518
rect 1582 68312 1638 68368
rect 5921 68026 5977 68028
rect 6001 68026 6057 68028
rect 6081 68026 6137 68028
rect 6161 68026 6217 68028
rect 5921 67974 5967 68026
rect 5967 67974 5977 68026
rect 6001 67974 6031 68026
rect 6031 67974 6043 68026
rect 6043 67974 6057 68026
rect 6081 67974 6095 68026
rect 6095 67974 6107 68026
rect 6107 67974 6137 68026
rect 6161 67974 6171 68026
rect 6171 67974 6217 68026
rect 5921 67972 5977 67974
rect 6001 67972 6057 67974
rect 6081 67972 6137 67974
rect 6161 67972 6217 67974
rect 1582 67668 1584 67688
rect 1584 67668 1636 67688
rect 1636 67668 1638 67688
rect 1582 67632 1638 67668
rect 10886 67482 10942 67484
rect 10966 67482 11022 67484
rect 11046 67482 11102 67484
rect 11126 67482 11182 67484
rect 10886 67430 10932 67482
rect 10932 67430 10942 67482
rect 10966 67430 10996 67482
rect 10996 67430 11008 67482
rect 11008 67430 11022 67482
rect 11046 67430 11060 67482
rect 11060 67430 11072 67482
rect 11072 67430 11102 67482
rect 11126 67430 11136 67482
rect 11136 67430 11182 67482
rect 10886 67428 10942 67430
rect 10966 67428 11022 67430
rect 11046 67428 11102 67430
rect 11126 67428 11182 67430
rect 1582 66952 1638 67008
rect 5921 66938 5977 66940
rect 6001 66938 6057 66940
rect 6081 66938 6137 66940
rect 6161 66938 6217 66940
rect 5921 66886 5967 66938
rect 5967 66886 5977 66938
rect 6001 66886 6031 66938
rect 6031 66886 6043 66938
rect 6043 66886 6057 66938
rect 6081 66886 6095 66938
rect 6095 66886 6107 66938
rect 6107 66886 6137 66938
rect 6161 66886 6171 66938
rect 6171 66886 6217 66938
rect 5921 66884 5977 66886
rect 6001 66884 6057 66886
rect 6081 66884 6137 66886
rect 6161 66884 6217 66886
rect 10886 66394 10942 66396
rect 10966 66394 11022 66396
rect 11046 66394 11102 66396
rect 11126 66394 11182 66396
rect 10886 66342 10932 66394
rect 10932 66342 10942 66394
rect 10966 66342 10996 66394
rect 10996 66342 11008 66394
rect 11008 66342 11022 66394
rect 11046 66342 11060 66394
rect 11060 66342 11072 66394
rect 11072 66342 11102 66394
rect 11126 66342 11136 66394
rect 11136 66342 11182 66394
rect 10886 66340 10942 66342
rect 10966 66340 11022 66342
rect 11046 66340 11102 66342
rect 11126 66340 11182 66342
rect 1582 66272 1638 66328
rect 5921 65850 5977 65852
rect 6001 65850 6057 65852
rect 6081 65850 6137 65852
rect 6161 65850 6217 65852
rect 5921 65798 5967 65850
rect 5967 65798 5977 65850
rect 6001 65798 6031 65850
rect 6031 65798 6043 65850
rect 6043 65798 6057 65850
rect 6081 65798 6095 65850
rect 6095 65798 6107 65850
rect 6107 65798 6137 65850
rect 6161 65798 6171 65850
rect 6171 65798 6217 65850
rect 5921 65796 5977 65798
rect 6001 65796 6057 65798
rect 6081 65796 6137 65798
rect 6161 65796 6217 65798
rect 1582 65728 1638 65784
rect 10886 65306 10942 65308
rect 10966 65306 11022 65308
rect 11046 65306 11102 65308
rect 11126 65306 11182 65308
rect 10886 65254 10932 65306
rect 10932 65254 10942 65306
rect 10966 65254 10996 65306
rect 10996 65254 11008 65306
rect 11008 65254 11022 65306
rect 11046 65254 11060 65306
rect 11060 65254 11072 65306
rect 11072 65254 11102 65306
rect 11126 65254 11136 65306
rect 11136 65254 11182 65306
rect 10886 65252 10942 65254
rect 10966 65252 11022 65254
rect 11046 65252 11102 65254
rect 11126 65252 11182 65254
rect 1582 65048 1638 65104
rect 5921 64762 5977 64764
rect 6001 64762 6057 64764
rect 6081 64762 6137 64764
rect 6161 64762 6217 64764
rect 5921 64710 5967 64762
rect 5967 64710 5977 64762
rect 6001 64710 6031 64762
rect 6031 64710 6043 64762
rect 6043 64710 6057 64762
rect 6081 64710 6095 64762
rect 6095 64710 6107 64762
rect 6107 64710 6137 64762
rect 6161 64710 6171 64762
rect 6171 64710 6217 64762
rect 5921 64708 5977 64710
rect 6001 64708 6057 64710
rect 6081 64708 6137 64710
rect 6161 64708 6217 64710
rect 1582 64404 1584 64424
rect 1584 64404 1636 64424
rect 1636 64404 1638 64424
rect 1582 64368 1638 64404
rect 10886 64218 10942 64220
rect 10966 64218 11022 64220
rect 11046 64218 11102 64220
rect 11126 64218 11182 64220
rect 10886 64166 10932 64218
rect 10932 64166 10942 64218
rect 10966 64166 10996 64218
rect 10996 64166 11008 64218
rect 11008 64166 11022 64218
rect 11046 64166 11060 64218
rect 11060 64166 11072 64218
rect 11072 64166 11102 64218
rect 11126 64166 11136 64218
rect 11136 64166 11182 64218
rect 10886 64164 10942 64166
rect 10966 64164 11022 64166
rect 11046 64164 11102 64166
rect 11126 64164 11182 64166
rect 1582 63688 1638 63744
rect 5921 63674 5977 63676
rect 6001 63674 6057 63676
rect 6081 63674 6137 63676
rect 6161 63674 6217 63676
rect 5921 63622 5967 63674
rect 5967 63622 5977 63674
rect 6001 63622 6031 63674
rect 6031 63622 6043 63674
rect 6043 63622 6057 63674
rect 6081 63622 6095 63674
rect 6095 63622 6107 63674
rect 6107 63622 6137 63674
rect 6161 63622 6171 63674
rect 6171 63622 6217 63674
rect 5921 63620 5977 63622
rect 6001 63620 6057 63622
rect 6081 63620 6137 63622
rect 6161 63620 6217 63622
rect 10886 63130 10942 63132
rect 10966 63130 11022 63132
rect 11046 63130 11102 63132
rect 11126 63130 11182 63132
rect 10886 63078 10932 63130
rect 10932 63078 10942 63130
rect 10966 63078 10996 63130
rect 10996 63078 11008 63130
rect 11008 63078 11022 63130
rect 11046 63078 11060 63130
rect 11060 63078 11072 63130
rect 11072 63078 11102 63130
rect 11126 63078 11136 63130
rect 11136 63078 11182 63130
rect 10886 63076 10942 63078
rect 10966 63076 11022 63078
rect 11046 63076 11102 63078
rect 11126 63076 11182 63078
rect 1582 63008 1638 63064
rect 5921 62586 5977 62588
rect 6001 62586 6057 62588
rect 6081 62586 6137 62588
rect 6161 62586 6217 62588
rect 5921 62534 5967 62586
rect 5967 62534 5977 62586
rect 6001 62534 6031 62586
rect 6031 62534 6043 62586
rect 6043 62534 6057 62586
rect 6081 62534 6095 62586
rect 6095 62534 6107 62586
rect 6107 62534 6137 62586
rect 6161 62534 6171 62586
rect 6171 62534 6217 62586
rect 5921 62532 5977 62534
rect 6001 62532 6057 62534
rect 6081 62532 6137 62534
rect 6161 62532 6217 62534
rect 1582 62328 1638 62384
rect 10886 62042 10942 62044
rect 10966 62042 11022 62044
rect 11046 62042 11102 62044
rect 11126 62042 11182 62044
rect 10886 61990 10932 62042
rect 10932 61990 10942 62042
rect 10966 61990 10996 62042
rect 10996 61990 11008 62042
rect 11008 61990 11022 62042
rect 11046 61990 11060 62042
rect 11060 61990 11072 62042
rect 11072 61990 11102 62042
rect 11126 61990 11136 62042
rect 11136 61990 11182 62042
rect 10886 61988 10942 61990
rect 10966 61988 11022 61990
rect 11046 61988 11102 61990
rect 11126 61988 11182 61990
rect 1582 61648 1638 61704
rect 5921 61498 5977 61500
rect 6001 61498 6057 61500
rect 6081 61498 6137 61500
rect 6161 61498 6217 61500
rect 5921 61446 5967 61498
rect 5967 61446 5977 61498
rect 6001 61446 6031 61498
rect 6031 61446 6043 61498
rect 6043 61446 6057 61498
rect 6081 61446 6095 61498
rect 6095 61446 6107 61498
rect 6107 61446 6137 61498
rect 6161 61446 6171 61498
rect 6171 61446 6217 61498
rect 5921 61444 5977 61446
rect 6001 61444 6057 61446
rect 6081 61444 6137 61446
rect 6161 61444 6217 61446
rect 1582 61140 1584 61160
rect 1584 61140 1636 61160
rect 1636 61140 1638 61160
rect 1582 61104 1638 61140
rect 10886 60954 10942 60956
rect 10966 60954 11022 60956
rect 11046 60954 11102 60956
rect 11126 60954 11182 60956
rect 10886 60902 10932 60954
rect 10932 60902 10942 60954
rect 10966 60902 10996 60954
rect 10996 60902 11008 60954
rect 11008 60902 11022 60954
rect 11046 60902 11060 60954
rect 11060 60902 11072 60954
rect 11072 60902 11102 60954
rect 11126 60902 11136 60954
rect 11136 60902 11182 60954
rect 10886 60900 10942 60902
rect 10966 60900 11022 60902
rect 11046 60900 11102 60902
rect 11126 60900 11182 60902
rect 1582 60424 1638 60480
rect 5921 60410 5977 60412
rect 6001 60410 6057 60412
rect 6081 60410 6137 60412
rect 6161 60410 6217 60412
rect 5921 60358 5967 60410
rect 5967 60358 5977 60410
rect 6001 60358 6031 60410
rect 6031 60358 6043 60410
rect 6043 60358 6057 60410
rect 6081 60358 6095 60410
rect 6095 60358 6107 60410
rect 6107 60358 6137 60410
rect 6161 60358 6171 60410
rect 6171 60358 6217 60410
rect 5921 60356 5977 60358
rect 6001 60356 6057 60358
rect 6081 60356 6137 60358
rect 6161 60356 6217 60358
rect 10886 59866 10942 59868
rect 10966 59866 11022 59868
rect 11046 59866 11102 59868
rect 11126 59866 11182 59868
rect 10886 59814 10932 59866
rect 10932 59814 10942 59866
rect 10966 59814 10996 59866
rect 10996 59814 11008 59866
rect 11008 59814 11022 59866
rect 11046 59814 11060 59866
rect 11060 59814 11072 59866
rect 11072 59814 11102 59866
rect 11126 59814 11136 59866
rect 11136 59814 11182 59866
rect 10886 59812 10942 59814
rect 10966 59812 11022 59814
rect 11046 59812 11102 59814
rect 11126 59812 11182 59814
rect 1582 59744 1638 59800
rect 5921 59322 5977 59324
rect 6001 59322 6057 59324
rect 6081 59322 6137 59324
rect 6161 59322 6217 59324
rect 5921 59270 5967 59322
rect 5967 59270 5977 59322
rect 6001 59270 6031 59322
rect 6031 59270 6043 59322
rect 6043 59270 6057 59322
rect 6081 59270 6095 59322
rect 6095 59270 6107 59322
rect 6107 59270 6137 59322
rect 6161 59270 6171 59322
rect 6171 59270 6217 59322
rect 5921 59268 5977 59270
rect 6001 59268 6057 59270
rect 6081 59268 6137 59270
rect 6161 59268 6217 59270
rect 1582 59064 1638 59120
rect 10886 58778 10942 58780
rect 10966 58778 11022 58780
rect 11046 58778 11102 58780
rect 11126 58778 11182 58780
rect 10886 58726 10932 58778
rect 10932 58726 10942 58778
rect 10966 58726 10996 58778
rect 10996 58726 11008 58778
rect 11008 58726 11022 58778
rect 11046 58726 11060 58778
rect 11060 58726 11072 58778
rect 11072 58726 11102 58778
rect 11126 58726 11136 58778
rect 11136 58726 11182 58778
rect 10886 58724 10942 58726
rect 10966 58724 11022 58726
rect 11046 58724 11102 58726
rect 11126 58724 11182 58726
rect 1582 58404 1638 58440
rect 1582 58384 1584 58404
rect 1584 58384 1636 58404
rect 1636 58384 1638 58404
rect 5921 58234 5977 58236
rect 6001 58234 6057 58236
rect 6081 58234 6137 58236
rect 6161 58234 6217 58236
rect 5921 58182 5967 58234
rect 5967 58182 5977 58234
rect 6001 58182 6031 58234
rect 6031 58182 6043 58234
rect 6043 58182 6057 58234
rect 6081 58182 6095 58234
rect 6095 58182 6107 58234
rect 6107 58182 6137 58234
rect 6161 58182 6171 58234
rect 6171 58182 6217 58234
rect 5921 58180 5977 58182
rect 6001 58180 6057 58182
rect 6081 58180 6137 58182
rect 6161 58180 6217 58182
rect 1582 57740 1584 57760
rect 1584 57740 1636 57760
rect 1636 57740 1638 57760
rect 1582 57704 1638 57740
rect 1582 57024 1638 57080
rect 1582 56480 1638 56536
rect 10886 57690 10942 57692
rect 10966 57690 11022 57692
rect 11046 57690 11102 57692
rect 11126 57690 11182 57692
rect 10886 57638 10932 57690
rect 10932 57638 10942 57690
rect 10966 57638 10996 57690
rect 10996 57638 11008 57690
rect 11008 57638 11022 57690
rect 11046 57638 11060 57690
rect 11060 57638 11072 57690
rect 11072 57638 11102 57690
rect 11126 57638 11136 57690
rect 11136 57638 11182 57690
rect 10886 57636 10942 57638
rect 10966 57636 11022 57638
rect 11046 57636 11102 57638
rect 11126 57636 11182 57638
rect 1582 55800 1638 55856
rect 1582 55140 1638 55176
rect 1582 55120 1584 55140
rect 1584 55120 1636 55140
rect 1636 55120 1638 55140
rect 1582 54476 1584 54496
rect 1584 54476 1636 54496
rect 1636 54476 1638 54496
rect 1582 54440 1638 54476
rect 1582 53760 1638 53816
rect 1582 53080 1638 53136
rect 1398 50496 1454 50552
rect 1582 51856 1638 51912
rect 1582 49816 1638 49872
rect 5921 57146 5977 57148
rect 6001 57146 6057 57148
rect 6081 57146 6137 57148
rect 6161 57146 6217 57148
rect 5921 57094 5967 57146
rect 5967 57094 5977 57146
rect 6001 57094 6031 57146
rect 6031 57094 6043 57146
rect 6043 57094 6057 57146
rect 6081 57094 6095 57146
rect 6095 57094 6107 57146
rect 6107 57094 6137 57146
rect 6161 57094 6171 57146
rect 6171 57094 6217 57146
rect 5921 57092 5977 57094
rect 6001 57092 6057 57094
rect 6081 57092 6137 57094
rect 6161 57092 6217 57094
rect 10886 56602 10942 56604
rect 10966 56602 11022 56604
rect 11046 56602 11102 56604
rect 11126 56602 11182 56604
rect 10886 56550 10932 56602
rect 10932 56550 10942 56602
rect 10966 56550 10996 56602
rect 10996 56550 11008 56602
rect 11008 56550 11022 56602
rect 11046 56550 11060 56602
rect 11060 56550 11072 56602
rect 11072 56550 11102 56602
rect 11126 56550 11136 56602
rect 11136 56550 11182 56602
rect 10886 56548 10942 56550
rect 10966 56548 11022 56550
rect 11046 56548 11102 56550
rect 11126 56548 11182 56550
rect 5921 56058 5977 56060
rect 6001 56058 6057 56060
rect 6081 56058 6137 56060
rect 6161 56058 6217 56060
rect 5921 56006 5967 56058
rect 5967 56006 5977 56058
rect 6001 56006 6031 56058
rect 6031 56006 6043 56058
rect 6043 56006 6057 56058
rect 6081 56006 6095 56058
rect 6095 56006 6107 56058
rect 6107 56006 6137 56058
rect 6161 56006 6171 56058
rect 6171 56006 6217 56058
rect 5921 56004 5977 56006
rect 6001 56004 6057 56006
rect 6081 56004 6137 56006
rect 6161 56004 6217 56006
rect 10886 55514 10942 55516
rect 10966 55514 11022 55516
rect 11046 55514 11102 55516
rect 11126 55514 11182 55516
rect 10886 55462 10932 55514
rect 10932 55462 10942 55514
rect 10966 55462 10996 55514
rect 10996 55462 11008 55514
rect 11008 55462 11022 55514
rect 11046 55462 11060 55514
rect 11060 55462 11072 55514
rect 11072 55462 11102 55514
rect 11126 55462 11136 55514
rect 11136 55462 11182 55514
rect 10886 55460 10942 55462
rect 10966 55460 11022 55462
rect 11046 55460 11102 55462
rect 11126 55460 11182 55462
rect 9494 55256 9550 55312
rect 1582 47232 1638 47288
rect 1582 46552 1638 46608
rect 1398 45872 1454 45928
rect 1490 45192 1546 45248
rect 1582 44512 1638 44568
rect 1582 42644 1584 42664
rect 1584 42644 1636 42664
rect 1636 42644 1638 42664
rect 1582 42608 1638 42644
rect 1582 41928 1638 41984
rect 1582 41248 1638 41304
rect 2042 52400 2098 52456
rect 2226 51176 2282 51232
rect 1582 40568 1638 40624
rect 1582 39888 1638 39944
rect 1582 39208 1638 39264
rect 1582 38528 1638 38584
rect 1582 37848 1638 37904
rect 1398 37304 1454 37360
rect 1582 36624 1638 36680
rect 1582 35944 1638 36000
rect 2226 47776 2282 47832
rect 2778 49136 2834 49192
rect 3422 48456 3478 48512
rect 2778 43832 2834 43888
rect 2226 43152 2282 43208
rect 1582 35264 1638 35320
rect 1582 34584 1638 34640
rect 1398 33904 1454 33960
rect 1582 33224 1638 33280
rect 1398 32680 1454 32736
rect 1490 32000 1546 32056
rect 1858 31864 1914 31920
rect 1582 31320 1638 31376
rect 1582 30640 1638 30696
rect 1582 29996 1584 30016
rect 1584 29996 1636 30016
rect 1636 29996 1638 30016
rect 1582 29960 1638 29996
rect 1582 29280 1638 29336
rect 1582 28600 1638 28656
rect 1582 28056 1638 28112
rect 1582 27376 1638 27432
rect 1582 26732 1584 26752
rect 1584 26732 1636 26752
rect 1636 26732 1638 26752
rect 1582 26696 1638 26732
rect 1582 26016 1638 26072
rect 1582 25336 1638 25392
rect 1582 24676 1638 24712
rect 1582 24656 1584 24676
rect 1584 24656 1636 24676
rect 1636 24656 1638 24676
rect 1582 24012 1584 24032
rect 1584 24012 1636 24032
rect 1636 24012 1638 24032
rect 1582 23976 1638 24012
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 1582 22752 1638 22808
rect 1582 22072 1638 22128
rect 1582 21412 1638 21448
rect 1582 21392 1584 21412
rect 1584 21392 1636 21412
rect 1636 21392 1638 21412
rect 1582 20748 1584 20768
rect 1584 20748 1636 20768
rect 1636 20748 1638 20768
rect 1582 20712 1638 20748
rect 1582 20032 1638 20088
rect 1582 19352 1638 19408
rect 1582 18808 1638 18864
rect 1582 18148 1638 18184
rect 1582 18128 1584 18148
rect 1584 18128 1636 18148
rect 1636 18128 1638 18148
rect 1582 17484 1584 17504
rect 1584 17484 1636 17504
rect 1636 17484 1638 17504
rect 1582 17448 1638 17484
rect 1582 16768 1638 16824
rect 1582 16088 1638 16144
rect 1582 15408 1638 15464
rect 1582 14764 1584 14784
rect 1584 14764 1636 14784
rect 1636 14764 1638 14784
rect 1582 14728 1638 14764
rect 1582 14220 1584 14240
rect 1584 14220 1636 14240
rect 1636 14220 1638 14240
rect 1582 14184 1638 14220
rect 1582 13504 1638 13560
rect 1582 12824 1638 12880
rect 1582 12144 1638 12200
rect 1582 11500 1584 11520
rect 1584 11500 1636 11520
rect 1636 11500 1638 11520
rect 1582 11464 1638 11500
rect 1582 10784 1638 10840
rect 1582 10104 1638 10160
rect 5921 54970 5977 54972
rect 6001 54970 6057 54972
rect 6081 54970 6137 54972
rect 6161 54970 6217 54972
rect 5921 54918 5967 54970
rect 5967 54918 5977 54970
rect 6001 54918 6031 54970
rect 6031 54918 6043 54970
rect 6043 54918 6057 54970
rect 6081 54918 6095 54970
rect 6095 54918 6107 54970
rect 6107 54918 6137 54970
rect 6161 54918 6171 54970
rect 6171 54918 6217 54970
rect 5921 54916 5977 54918
rect 6001 54916 6057 54918
rect 6081 54916 6137 54918
rect 6161 54916 6217 54918
rect 5921 53882 5977 53884
rect 6001 53882 6057 53884
rect 6081 53882 6137 53884
rect 6161 53882 6217 53884
rect 5921 53830 5967 53882
rect 5967 53830 5977 53882
rect 6001 53830 6031 53882
rect 6031 53830 6043 53882
rect 6043 53830 6057 53882
rect 6081 53830 6095 53882
rect 6095 53830 6107 53882
rect 6107 53830 6137 53882
rect 6161 53830 6171 53882
rect 6171 53830 6217 53882
rect 5921 53828 5977 53830
rect 6001 53828 6057 53830
rect 6081 53828 6137 53830
rect 6161 53828 6217 53830
rect 5921 52794 5977 52796
rect 6001 52794 6057 52796
rect 6081 52794 6137 52796
rect 6161 52794 6217 52796
rect 5921 52742 5967 52794
rect 5967 52742 5977 52794
rect 6001 52742 6031 52794
rect 6031 52742 6043 52794
rect 6043 52742 6057 52794
rect 6081 52742 6095 52794
rect 6095 52742 6107 52794
rect 6107 52742 6137 52794
rect 6161 52742 6171 52794
rect 6171 52742 6217 52794
rect 5921 52740 5977 52742
rect 6001 52740 6057 52742
rect 6081 52740 6137 52742
rect 6161 52740 6217 52742
rect 5921 51706 5977 51708
rect 6001 51706 6057 51708
rect 6081 51706 6137 51708
rect 6161 51706 6217 51708
rect 5921 51654 5967 51706
rect 5967 51654 5977 51706
rect 6001 51654 6031 51706
rect 6031 51654 6043 51706
rect 6043 51654 6057 51706
rect 6081 51654 6095 51706
rect 6095 51654 6107 51706
rect 6107 51654 6137 51706
rect 6161 51654 6171 51706
rect 6171 51654 6217 51706
rect 5921 51652 5977 51654
rect 6001 51652 6057 51654
rect 6081 51652 6137 51654
rect 6161 51652 6217 51654
rect 5921 50618 5977 50620
rect 6001 50618 6057 50620
rect 6081 50618 6137 50620
rect 6161 50618 6217 50620
rect 5921 50566 5967 50618
rect 5967 50566 5977 50618
rect 6001 50566 6031 50618
rect 6031 50566 6043 50618
rect 6043 50566 6057 50618
rect 6081 50566 6095 50618
rect 6095 50566 6107 50618
rect 6107 50566 6137 50618
rect 6161 50566 6171 50618
rect 6171 50566 6217 50618
rect 5921 50564 5977 50566
rect 6001 50564 6057 50566
rect 6081 50564 6137 50566
rect 6161 50564 6217 50566
rect 5921 49530 5977 49532
rect 6001 49530 6057 49532
rect 6081 49530 6137 49532
rect 6161 49530 6217 49532
rect 5921 49478 5967 49530
rect 5967 49478 5977 49530
rect 6001 49478 6031 49530
rect 6031 49478 6043 49530
rect 6043 49478 6057 49530
rect 6081 49478 6095 49530
rect 6095 49478 6107 49530
rect 6107 49478 6137 49530
rect 6161 49478 6171 49530
rect 6171 49478 6217 49530
rect 5921 49476 5977 49478
rect 6001 49476 6057 49478
rect 6081 49476 6137 49478
rect 6161 49476 6217 49478
rect 5921 48442 5977 48444
rect 6001 48442 6057 48444
rect 6081 48442 6137 48444
rect 6161 48442 6217 48444
rect 5921 48390 5967 48442
rect 5967 48390 5977 48442
rect 6001 48390 6031 48442
rect 6031 48390 6043 48442
rect 6043 48390 6057 48442
rect 6081 48390 6095 48442
rect 6095 48390 6107 48442
rect 6107 48390 6137 48442
rect 6161 48390 6171 48442
rect 6171 48390 6217 48442
rect 5921 48388 5977 48390
rect 6001 48388 6057 48390
rect 6081 48388 6137 48390
rect 6161 48388 6217 48390
rect 5921 47354 5977 47356
rect 6001 47354 6057 47356
rect 6081 47354 6137 47356
rect 6161 47354 6217 47356
rect 5921 47302 5967 47354
rect 5967 47302 5977 47354
rect 6001 47302 6031 47354
rect 6031 47302 6043 47354
rect 6043 47302 6057 47354
rect 6081 47302 6095 47354
rect 6095 47302 6107 47354
rect 6107 47302 6137 47354
rect 6161 47302 6171 47354
rect 6171 47302 6217 47354
rect 5921 47300 5977 47302
rect 6001 47300 6057 47302
rect 6081 47300 6137 47302
rect 6161 47300 6217 47302
rect 5921 46266 5977 46268
rect 6001 46266 6057 46268
rect 6081 46266 6137 46268
rect 6161 46266 6217 46268
rect 5921 46214 5967 46266
rect 5967 46214 5977 46266
rect 6001 46214 6031 46266
rect 6031 46214 6043 46266
rect 6043 46214 6057 46266
rect 6081 46214 6095 46266
rect 6095 46214 6107 46266
rect 6107 46214 6137 46266
rect 6161 46214 6171 46266
rect 6171 46214 6217 46266
rect 5921 46212 5977 46214
rect 6001 46212 6057 46214
rect 6081 46212 6137 46214
rect 6161 46212 6217 46214
rect 5921 45178 5977 45180
rect 6001 45178 6057 45180
rect 6081 45178 6137 45180
rect 6161 45178 6217 45180
rect 5921 45126 5967 45178
rect 5967 45126 5977 45178
rect 6001 45126 6031 45178
rect 6031 45126 6043 45178
rect 6043 45126 6057 45178
rect 6081 45126 6095 45178
rect 6095 45126 6107 45178
rect 6107 45126 6137 45178
rect 6161 45126 6171 45178
rect 6171 45126 6217 45178
rect 5921 45124 5977 45126
rect 6001 45124 6057 45126
rect 6081 45124 6137 45126
rect 6161 45124 6217 45126
rect 5921 44090 5977 44092
rect 6001 44090 6057 44092
rect 6081 44090 6137 44092
rect 6161 44090 6217 44092
rect 5921 44038 5967 44090
rect 5967 44038 5977 44090
rect 6001 44038 6031 44090
rect 6031 44038 6043 44090
rect 6043 44038 6057 44090
rect 6081 44038 6095 44090
rect 6095 44038 6107 44090
rect 6107 44038 6137 44090
rect 6161 44038 6171 44090
rect 6171 44038 6217 44090
rect 5921 44036 5977 44038
rect 6001 44036 6057 44038
rect 6081 44036 6137 44038
rect 6161 44036 6217 44038
rect 5921 43002 5977 43004
rect 6001 43002 6057 43004
rect 6081 43002 6137 43004
rect 6161 43002 6217 43004
rect 5921 42950 5967 43002
rect 5967 42950 5977 43002
rect 6001 42950 6031 43002
rect 6031 42950 6043 43002
rect 6043 42950 6057 43002
rect 6081 42950 6095 43002
rect 6095 42950 6107 43002
rect 6107 42950 6137 43002
rect 6161 42950 6171 43002
rect 6171 42950 6217 43002
rect 5921 42948 5977 42950
rect 6001 42948 6057 42950
rect 6081 42948 6137 42950
rect 6161 42948 6217 42950
rect 5921 41914 5977 41916
rect 6001 41914 6057 41916
rect 6081 41914 6137 41916
rect 6161 41914 6217 41916
rect 5921 41862 5967 41914
rect 5967 41862 5977 41914
rect 6001 41862 6031 41914
rect 6031 41862 6043 41914
rect 6043 41862 6057 41914
rect 6081 41862 6095 41914
rect 6095 41862 6107 41914
rect 6107 41862 6137 41914
rect 6161 41862 6171 41914
rect 6171 41862 6217 41914
rect 5921 41860 5977 41862
rect 6001 41860 6057 41862
rect 6081 41860 6137 41862
rect 6161 41860 6217 41862
rect 5921 40826 5977 40828
rect 6001 40826 6057 40828
rect 6081 40826 6137 40828
rect 6161 40826 6217 40828
rect 5921 40774 5967 40826
rect 5967 40774 5977 40826
rect 6001 40774 6031 40826
rect 6031 40774 6043 40826
rect 6043 40774 6057 40826
rect 6081 40774 6095 40826
rect 6095 40774 6107 40826
rect 6107 40774 6137 40826
rect 6161 40774 6171 40826
rect 6171 40774 6217 40826
rect 5921 40772 5977 40774
rect 6001 40772 6057 40774
rect 6081 40772 6137 40774
rect 6161 40772 6217 40774
rect 5921 39738 5977 39740
rect 6001 39738 6057 39740
rect 6081 39738 6137 39740
rect 6161 39738 6217 39740
rect 5921 39686 5967 39738
rect 5967 39686 5977 39738
rect 6001 39686 6031 39738
rect 6031 39686 6043 39738
rect 6043 39686 6057 39738
rect 6081 39686 6095 39738
rect 6095 39686 6107 39738
rect 6107 39686 6137 39738
rect 6161 39686 6171 39738
rect 6171 39686 6217 39738
rect 5921 39684 5977 39686
rect 6001 39684 6057 39686
rect 6081 39684 6137 39686
rect 6161 39684 6217 39686
rect 5921 38650 5977 38652
rect 6001 38650 6057 38652
rect 6081 38650 6137 38652
rect 6161 38650 6217 38652
rect 5921 38598 5967 38650
rect 5967 38598 5977 38650
rect 6001 38598 6031 38650
rect 6031 38598 6043 38650
rect 6043 38598 6057 38650
rect 6081 38598 6095 38650
rect 6095 38598 6107 38650
rect 6107 38598 6137 38650
rect 6161 38598 6171 38650
rect 6171 38598 6217 38650
rect 5921 38596 5977 38598
rect 6001 38596 6057 38598
rect 6081 38596 6137 38598
rect 6161 38596 6217 38598
rect 5921 37562 5977 37564
rect 6001 37562 6057 37564
rect 6081 37562 6137 37564
rect 6161 37562 6217 37564
rect 5921 37510 5967 37562
rect 5967 37510 5977 37562
rect 6001 37510 6031 37562
rect 6031 37510 6043 37562
rect 6043 37510 6057 37562
rect 6081 37510 6095 37562
rect 6095 37510 6107 37562
rect 6107 37510 6137 37562
rect 6161 37510 6171 37562
rect 6171 37510 6217 37562
rect 5921 37508 5977 37510
rect 6001 37508 6057 37510
rect 6081 37508 6137 37510
rect 6161 37508 6217 37510
rect 5921 36474 5977 36476
rect 6001 36474 6057 36476
rect 6081 36474 6137 36476
rect 6161 36474 6217 36476
rect 5921 36422 5967 36474
rect 5967 36422 5977 36474
rect 6001 36422 6031 36474
rect 6031 36422 6043 36474
rect 6043 36422 6057 36474
rect 6081 36422 6095 36474
rect 6095 36422 6107 36474
rect 6107 36422 6137 36474
rect 6161 36422 6171 36474
rect 6171 36422 6217 36474
rect 5921 36420 5977 36422
rect 6001 36420 6057 36422
rect 6081 36420 6137 36422
rect 6161 36420 6217 36422
rect 5921 35386 5977 35388
rect 6001 35386 6057 35388
rect 6081 35386 6137 35388
rect 6161 35386 6217 35388
rect 5921 35334 5967 35386
rect 5967 35334 5977 35386
rect 6001 35334 6031 35386
rect 6031 35334 6043 35386
rect 6043 35334 6057 35386
rect 6081 35334 6095 35386
rect 6095 35334 6107 35386
rect 6107 35334 6137 35386
rect 6161 35334 6171 35386
rect 6171 35334 6217 35386
rect 5921 35332 5977 35334
rect 6001 35332 6057 35334
rect 6081 35332 6137 35334
rect 6161 35332 6217 35334
rect 5921 34298 5977 34300
rect 6001 34298 6057 34300
rect 6081 34298 6137 34300
rect 6161 34298 6217 34300
rect 5921 34246 5967 34298
rect 5967 34246 5977 34298
rect 6001 34246 6031 34298
rect 6031 34246 6043 34298
rect 6043 34246 6057 34298
rect 6081 34246 6095 34298
rect 6095 34246 6107 34298
rect 6107 34246 6137 34298
rect 6161 34246 6171 34298
rect 6171 34246 6217 34298
rect 5921 34244 5977 34246
rect 6001 34244 6057 34246
rect 6081 34244 6137 34246
rect 6161 34244 6217 34246
rect 5921 33210 5977 33212
rect 6001 33210 6057 33212
rect 6081 33210 6137 33212
rect 6161 33210 6217 33212
rect 5921 33158 5967 33210
rect 5967 33158 5977 33210
rect 6001 33158 6031 33210
rect 6031 33158 6043 33210
rect 6043 33158 6057 33210
rect 6081 33158 6095 33210
rect 6095 33158 6107 33210
rect 6107 33158 6137 33210
rect 6161 33158 6171 33210
rect 6171 33158 6217 33210
rect 5921 33156 5977 33158
rect 6001 33156 6057 33158
rect 6081 33156 6137 33158
rect 6161 33156 6217 33158
rect 5921 32122 5977 32124
rect 6001 32122 6057 32124
rect 6081 32122 6137 32124
rect 6161 32122 6217 32124
rect 5921 32070 5967 32122
rect 5967 32070 5977 32122
rect 6001 32070 6031 32122
rect 6031 32070 6043 32122
rect 6043 32070 6057 32122
rect 6081 32070 6095 32122
rect 6095 32070 6107 32122
rect 6107 32070 6137 32122
rect 6161 32070 6171 32122
rect 6171 32070 6217 32122
rect 5921 32068 5977 32070
rect 6001 32068 6057 32070
rect 6081 32068 6137 32070
rect 6161 32068 6217 32070
rect 5921 31034 5977 31036
rect 6001 31034 6057 31036
rect 6081 31034 6137 31036
rect 6161 31034 6217 31036
rect 5921 30982 5967 31034
rect 5967 30982 5977 31034
rect 6001 30982 6031 31034
rect 6031 30982 6043 31034
rect 6043 30982 6057 31034
rect 6081 30982 6095 31034
rect 6095 30982 6107 31034
rect 6107 30982 6137 31034
rect 6161 30982 6171 31034
rect 6171 30982 6217 31034
rect 5921 30980 5977 30982
rect 6001 30980 6057 30982
rect 6081 30980 6137 30982
rect 6161 30980 6217 30982
rect 5921 29946 5977 29948
rect 6001 29946 6057 29948
rect 6081 29946 6137 29948
rect 6161 29946 6217 29948
rect 5921 29894 5967 29946
rect 5967 29894 5977 29946
rect 6001 29894 6031 29946
rect 6031 29894 6043 29946
rect 6043 29894 6057 29946
rect 6081 29894 6095 29946
rect 6095 29894 6107 29946
rect 6107 29894 6137 29946
rect 6161 29894 6171 29946
rect 6171 29894 6217 29946
rect 5921 29892 5977 29894
rect 6001 29892 6057 29894
rect 6081 29892 6137 29894
rect 6161 29892 6217 29894
rect 5921 28858 5977 28860
rect 6001 28858 6057 28860
rect 6081 28858 6137 28860
rect 6161 28858 6217 28860
rect 5921 28806 5967 28858
rect 5967 28806 5977 28858
rect 6001 28806 6031 28858
rect 6031 28806 6043 28858
rect 6043 28806 6057 28858
rect 6081 28806 6095 28858
rect 6095 28806 6107 28858
rect 6107 28806 6137 28858
rect 6161 28806 6171 28858
rect 6171 28806 6217 28858
rect 5921 28804 5977 28806
rect 6001 28804 6057 28806
rect 6081 28804 6137 28806
rect 6161 28804 6217 28806
rect 5921 27770 5977 27772
rect 6001 27770 6057 27772
rect 6081 27770 6137 27772
rect 6161 27770 6217 27772
rect 5921 27718 5967 27770
rect 5967 27718 5977 27770
rect 6001 27718 6031 27770
rect 6031 27718 6043 27770
rect 6043 27718 6057 27770
rect 6081 27718 6095 27770
rect 6095 27718 6107 27770
rect 6107 27718 6137 27770
rect 6161 27718 6171 27770
rect 6171 27718 6217 27770
rect 5921 27716 5977 27718
rect 6001 27716 6057 27718
rect 6081 27716 6137 27718
rect 6161 27716 6217 27718
rect 5921 26682 5977 26684
rect 6001 26682 6057 26684
rect 6081 26682 6137 26684
rect 6161 26682 6217 26684
rect 5921 26630 5967 26682
rect 5967 26630 5977 26682
rect 6001 26630 6031 26682
rect 6031 26630 6043 26682
rect 6043 26630 6057 26682
rect 6081 26630 6095 26682
rect 6095 26630 6107 26682
rect 6107 26630 6137 26682
rect 6161 26630 6171 26682
rect 6171 26630 6217 26682
rect 5921 26628 5977 26630
rect 6001 26628 6057 26630
rect 6081 26628 6137 26630
rect 6161 26628 6217 26630
rect 5921 25594 5977 25596
rect 6001 25594 6057 25596
rect 6081 25594 6137 25596
rect 6161 25594 6217 25596
rect 5921 25542 5967 25594
rect 5967 25542 5977 25594
rect 6001 25542 6031 25594
rect 6031 25542 6043 25594
rect 6043 25542 6057 25594
rect 6081 25542 6095 25594
rect 6095 25542 6107 25594
rect 6107 25542 6137 25594
rect 6161 25542 6171 25594
rect 6171 25542 6217 25594
rect 5921 25540 5977 25542
rect 6001 25540 6057 25542
rect 6081 25540 6137 25542
rect 6161 25540 6217 25542
rect 5921 24506 5977 24508
rect 6001 24506 6057 24508
rect 6081 24506 6137 24508
rect 6161 24506 6217 24508
rect 5921 24454 5967 24506
rect 5967 24454 5977 24506
rect 6001 24454 6031 24506
rect 6031 24454 6043 24506
rect 6043 24454 6057 24506
rect 6081 24454 6095 24506
rect 6095 24454 6107 24506
rect 6107 24454 6137 24506
rect 6161 24454 6171 24506
rect 6171 24454 6217 24506
rect 5921 24452 5977 24454
rect 6001 24452 6057 24454
rect 6081 24452 6137 24454
rect 6161 24452 6217 24454
rect 5921 23418 5977 23420
rect 6001 23418 6057 23420
rect 6081 23418 6137 23420
rect 6161 23418 6217 23420
rect 5921 23366 5967 23418
rect 5967 23366 5977 23418
rect 6001 23366 6031 23418
rect 6031 23366 6043 23418
rect 6043 23366 6057 23418
rect 6081 23366 6095 23418
rect 6095 23366 6107 23418
rect 6107 23366 6137 23418
rect 6161 23366 6171 23418
rect 6171 23366 6217 23418
rect 5921 23364 5977 23366
rect 6001 23364 6057 23366
rect 6081 23364 6137 23366
rect 6161 23364 6217 23366
rect 5921 22330 5977 22332
rect 6001 22330 6057 22332
rect 6081 22330 6137 22332
rect 6161 22330 6217 22332
rect 5921 22278 5967 22330
rect 5967 22278 5977 22330
rect 6001 22278 6031 22330
rect 6031 22278 6043 22330
rect 6043 22278 6057 22330
rect 6081 22278 6095 22330
rect 6095 22278 6107 22330
rect 6107 22278 6137 22330
rect 6161 22278 6171 22330
rect 6171 22278 6217 22330
rect 5921 22276 5977 22278
rect 6001 22276 6057 22278
rect 6081 22276 6137 22278
rect 6161 22276 6217 22278
rect 5921 21242 5977 21244
rect 6001 21242 6057 21244
rect 6081 21242 6137 21244
rect 6161 21242 6217 21244
rect 5921 21190 5967 21242
rect 5967 21190 5977 21242
rect 6001 21190 6031 21242
rect 6031 21190 6043 21242
rect 6043 21190 6057 21242
rect 6081 21190 6095 21242
rect 6095 21190 6107 21242
rect 6107 21190 6137 21242
rect 6161 21190 6171 21242
rect 6171 21190 6217 21242
rect 5921 21188 5977 21190
rect 6001 21188 6057 21190
rect 6081 21188 6137 21190
rect 6161 21188 6217 21190
rect 5921 20154 5977 20156
rect 6001 20154 6057 20156
rect 6081 20154 6137 20156
rect 6161 20154 6217 20156
rect 5921 20102 5967 20154
rect 5967 20102 5977 20154
rect 6001 20102 6031 20154
rect 6031 20102 6043 20154
rect 6043 20102 6057 20154
rect 6081 20102 6095 20154
rect 6095 20102 6107 20154
rect 6107 20102 6137 20154
rect 6161 20102 6171 20154
rect 6171 20102 6217 20154
rect 5921 20100 5977 20102
rect 6001 20100 6057 20102
rect 6081 20100 6137 20102
rect 6161 20100 6217 20102
rect 5921 19066 5977 19068
rect 6001 19066 6057 19068
rect 6081 19066 6137 19068
rect 6161 19066 6217 19068
rect 5921 19014 5967 19066
rect 5967 19014 5977 19066
rect 6001 19014 6031 19066
rect 6031 19014 6043 19066
rect 6043 19014 6057 19066
rect 6081 19014 6095 19066
rect 6095 19014 6107 19066
rect 6107 19014 6137 19066
rect 6161 19014 6171 19066
rect 6171 19014 6217 19066
rect 5921 19012 5977 19014
rect 6001 19012 6057 19014
rect 6081 19012 6137 19014
rect 6161 19012 6217 19014
rect 5921 17978 5977 17980
rect 6001 17978 6057 17980
rect 6081 17978 6137 17980
rect 6161 17978 6217 17980
rect 5921 17926 5967 17978
rect 5967 17926 5977 17978
rect 6001 17926 6031 17978
rect 6031 17926 6043 17978
rect 6043 17926 6057 17978
rect 6081 17926 6095 17978
rect 6095 17926 6107 17978
rect 6107 17926 6137 17978
rect 6161 17926 6171 17978
rect 6171 17926 6217 17978
rect 5921 17924 5977 17926
rect 6001 17924 6057 17926
rect 6081 17924 6137 17926
rect 6161 17924 6217 17926
rect 5921 16890 5977 16892
rect 6001 16890 6057 16892
rect 6081 16890 6137 16892
rect 6161 16890 6217 16892
rect 5921 16838 5967 16890
rect 5967 16838 5977 16890
rect 6001 16838 6031 16890
rect 6031 16838 6043 16890
rect 6043 16838 6057 16890
rect 6081 16838 6095 16890
rect 6095 16838 6107 16890
rect 6107 16838 6137 16890
rect 6161 16838 6171 16890
rect 6171 16838 6217 16890
rect 5921 16836 5977 16838
rect 6001 16836 6057 16838
rect 6081 16836 6137 16838
rect 6161 16836 6217 16838
rect 5921 15802 5977 15804
rect 6001 15802 6057 15804
rect 6081 15802 6137 15804
rect 6161 15802 6217 15804
rect 5921 15750 5967 15802
rect 5967 15750 5977 15802
rect 6001 15750 6031 15802
rect 6031 15750 6043 15802
rect 6043 15750 6057 15802
rect 6081 15750 6095 15802
rect 6095 15750 6107 15802
rect 6107 15750 6137 15802
rect 6161 15750 6171 15802
rect 6171 15750 6217 15802
rect 5921 15748 5977 15750
rect 6001 15748 6057 15750
rect 6081 15748 6137 15750
rect 6161 15748 6217 15750
rect 5921 14714 5977 14716
rect 6001 14714 6057 14716
rect 6081 14714 6137 14716
rect 6161 14714 6217 14716
rect 5921 14662 5967 14714
rect 5967 14662 5977 14714
rect 6001 14662 6031 14714
rect 6031 14662 6043 14714
rect 6043 14662 6057 14714
rect 6081 14662 6095 14714
rect 6095 14662 6107 14714
rect 6107 14662 6137 14714
rect 6161 14662 6171 14714
rect 6171 14662 6217 14714
rect 5921 14660 5977 14662
rect 6001 14660 6057 14662
rect 6081 14660 6137 14662
rect 6161 14660 6217 14662
rect 5921 13626 5977 13628
rect 6001 13626 6057 13628
rect 6081 13626 6137 13628
rect 6161 13626 6217 13628
rect 5921 13574 5967 13626
rect 5967 13574 5977 13626
rect 6001 13574 6031 13626
rect 6031 13574 6043 13626
rect 6043 13574 6057 13626
rect 6081 13574 6095 13626
rect 6095 13574 6107 13626
rect 6107 13574 6137 13626
rect 6161 13574 6171 13626
rect 6171 13574 6217 13626
rect 5921 13572 5977 13574
rect 6001 13572 6057 13574
rect 6081 13572 6137 13574
rect 6161 13572 6217 13574
rect 5921 12538 5977 12540
rect 6001 12538 6057 12540
rect 6081 12538 6137 12540
rect 6161 12538 6217 12540
rect 5921 12486 5967 12538
rect 5967 12486 5977 12538
rect 6001 12486 6031 12538
rect 6031 12486 6043 12538
rect 6043 12486 6057 12538
rect 6081 12486 6095 12538
rect 6095 12486 6107 12538
rect 6107 12486 6137 12538
rect 6161 12486 6171 12538
rect 6171 12486 6217 12538
rect 5921 12484 5977 12486
rect 6001 12484 6057 12486
rect 6081 12484 6137 12486
rect 6161 12484 6217 12486
rect 5921 11450 5977 11452
rect 6001 11450 6057 11452
rect 6081 11450 6137 11452
rect 6161 11450 6217 11452
rect 5921 11398 5967 11450
rect 5967 11398 5977 11450
rect 6001 11398 6031 11450
rect 6031 11398 6043 11450
rect 6043 11398 6057 11450
rect 6081 11398 6095 11450
rect 6095 11398 6107 11450
rect 6107 11398 6137 11450
rect 6161 11398 6171 11450
rect 6171 11398 6217 11450
rect 5921 11396 5977 11398
rect 6001 11396 6057 11398
rect 6081 11396 6137 11398
rect 6161 11396 6217 11398
rect 5921 10362 5977 10364
rect 6001 10362 6057 10364
rect 6081 10362 6137 10364
rect 6161 10362 6217 10364
rect 5921 10310 5967 10362
rect 5967 10310 5977 10362
rect 6001 10310 6031 10362
rect 6031 10310 6043 10362
rect 6043 10310 6057 10362
rect 6081 10310 6095 10362
rect 6095 10310 6107 10362
rect 6107 10310 6137 10362
rect 6161 10310 6171 10362
rect 6171 10310 6217 10362
rect 5921 10308 5977 10310
rect 6001 10308 6057 10310
rect 6081 10308 6137 10310
rect 6161 10308 6217 10310
rect 1582 9560 1638 9616
rect 5921 9274 5977 9276
rect 6001 9274 6057 9276
rect 6081 9274 6137 9276
rect 6161 9274 6217 9276
rect 5921 9222 5967 9274
rect 5967 9222 5977 9274
rect 6001 9222 6031 9274
rect 6031 9222 6043 9274
rect 6043 9222 6057 9274
rect 6081 9222 6095 9274
rect 6095 9222 6107 9274
rect 6107 9222 6137 9274
rect 6161 9222 6171 9274
rect 6171 9222 6217 9274
rect 5921 9220 5977 9222
rect 6001 9220 6057 9222
rect 6081 9220 6137 9222
rect 6161 9220 6217 9222
rect 1582 8880 1638 8936
rect 1582 8200 1638 8256
rect 5921 8186 5977 8188
rect 6001 8186 6057 8188
rect 6081 8186 6137 8188
rect 6161 8186 6217 8188
rect 5921 8134 5967 8186
rect 5967 8134 5977 8186
rect 6001 8134 6031 8186
rect 6031 8134 6043 8186
rect 6043 8134 6057 8186
rect 6081 8134 6095 8186
rect 6095 8134 6107 8186
rect 6107 8134 6137 8186
rect 6161 8134 6171 8186
rect 6171 8134 6217 8186
rect 5921 8132 5977 8134
rect 6001 8132 6057 8134
rect 6081 8132 6137 8134
rect 6161 8132 6217 8134
rect 1582 7520 1638 7576
rect 1582 6840 1638 6896
rect 9402 43696 9458 43752
rect 10886 54426 10942 54428
rect 10966 54426 11022 54428
rect 11046 54426 11102 54428
rect 11126 54426 11182 54428
rect 10886 54374 10932 54426
rect 10932 54374 10942 54426
rect 10966 54374 10996 54426
rect 10996 54374 11008 54426
rect 11008 54374 11022 54426
rect 11046 54374 11060 54426
rect 11060 54374 11072 54426
rect 11072 54374 11102 54426
rect 11126 54374 11136 54426
rect 11136 54374 11182 54426
rect 10886 54372 10942 54374
rect 10966 54372 11022 54374
rect 11046 54372 11102 54374
rect 11126 54372 11182 54374
rect 10886 53338 10942 53340
rect 10966 53338 11022 53340
rect 11046 53338 11102 53340
rect 11126 53338 11182 53340
rect 10886 53286 10932 53338
rect 10932 53286 10942 53338
rect 10966 53286 10996 53338
rect 10996 53286 11008 53338
rect 11008 53286 11022 53338
rect 11046 53286 11060 53338
rect 11060 53286 11072 53338
rect 11072 53286 11102 53338
rect 11126 53286 11136 53338
rect 11136 53286 11182 53338
rect 10886 53284 10942 53286
rect 10966 53284 11022 53286
rect 11046 53284 11102 53286
rect 11126 53284 11182 53286
rect 10886 52250 10942 52252
rect 10966 52250 11022 52252
rect 11046 52250 11102 52252
rect 11126 52250 11182 52252
rect 10886 52198 10932 52250
rect 10932 52198 10942 52250
rect 10966 52198 10996 52250
rect 10996 52198 11008 52250
rect 11008 52198 11022 52250
rect 11046 52198 11060 52250
rect 11060 52198 11072 52250
rect 11072 52198 11102 52250
rect 11126 52198 11136 52250
rect 11136 52198 11182 52250
rect 10886 52196 10942 52198
rect 10966 52196 11022 52198
rect 11046 52196 11102 52198
rect 11126 52196 11182 52198
rect 10886 51162 10942 51164
rect 10966 51162 11022 51164
rect 11046 51162 11102 51164
rect 11126 51162 11182 51164
rect 10886 51110 10932 51162
rect 10932 51110 10942 51162
rect 10966 51110 10996 51162
rect 10996 51110 11008 51162
rect 11008 51110 11022 51162
rect 11046 51110 11060 51162
rect 11060 51110 11072 51162
rect 11072 51110 11102 51162
rect 11126 51110 11136 51162
rect 11136 51110 11182 51162
rect 10886 51108 10942 51110
rect 10966 51108 11022 51110
rect 11046 51108 11102 51110
rect 11126 51108 11182 51110
rect 9494 36760 9550 36816
rect 10414 36624 10470 36680
rect 10886 50074 10942 50076
rect 10966 50074 11022 50076
rect 11046 50074 11102 50076
rect 11126 50074 11182 50076
rect 10886 50022 10932 50074
rect 10932 50022 10942 50074
rect 10966 50022 10996 50074
rect 10996 50022 11008 50074
rect 11008 50022 11022 50074
rect 11046 50022 11060 50074
rect 11060 50022 11072 50074
rect 11072 50022 11102 50074
rect 11126 50022 11136 50074
rect 11136 50022 11182 50074
rect 10886 50020 10942 50022
rect 10966 50020 11022 50022
rect 11046 50020 11102 50022
rect 11126 50020 11182 50022
rect 10886 48986 10942 48988
rect 10966 48986 11022 48988
rect 11046 48986 11102 48988
rect 11126 48986 11182 48988
rect 10886 48934 10932 48986
rect 10932 48934 10942 48986
rect 10966 48934 10996 48986
rect 10996 48934 11008 48986
rect 11008 48934 11022 48986
rect 11046 48934 11060 48986
rect 11060 48934 11072 48986
rect 11072 48934 11102 48986
rect 11126 48934 11136 48986
rect 11136 48934 11182 48986
rect 10886 48932 10942 48934
rect 10966 48932 11022 48934
rect 11046 48932 11102 48934
rect 11126 48932 11182 48934
rect 10886 47898 10942 47900
rect 10966 47898 11022 47900
rect 11046 47898 11102 47900
rect 11126 47898 11182 47900
rect 10886 47846 10932 47898
rect 10932 47846 10942 47898
rect 10966 47846 10996 47898
rect 10996 47846 11008 47898
rect 11008 47846 11022 47898
rect 11046 47846 11060 47898
rect 11060 47846 11072 47898
rect 11072 47846 11102 47898
rect 11126 47846 11136 47898
rect 11136 47846 11182 47898
rect 10886 47844 10942 47846
rect 10966 47844 11022 47846
rect 11046 47844 11102 47846
rect 11126 47844 11182 47846
rect 10886 46810 10942 46812
rect 10966 46810 11022 46812
rect 11046 46810 11102 46812
rect 11126 46810 11182 46812
rect 10886 46758 10932 46810
rect 10932 46758 10942 46810
rect 10966 46758 10996 46810
rect 10996 46758 11008 46810
rect 11008 46758 11022 46810
rect 11046 46758 11060 46810
rect 11060 46758 11072 46810
rect 11072 46758 11102 46810
rect 11126 46758 11136 46810
rect 11136 46758 11182 46810
rect 10886 46756 10942 46758
rect 10966 46756 11022 46758
rect 11046 46756 11102 46758
rect 11126 46756 11182 46758
rect 10886 45722 10942 45724
rect 10966 45722 11022 45724
rect 11046 45722 11102 45724
rect 11126 45722 11182 45724
rect 10886 45670 10932 45722
rect 10932 45670 10942 45722
rect 10966 45670 10996 45722
rect 10996 45670 11008 45722
rect 11008 45670 11022 45722
rect 11046 45670 11060 45722
rect 11060 45670 11072 45722
rect 11072 45670 11102 45722
rect 11126 45670 11136 45722
rect 11136 45670 11182 45722
rect 10886 45668 10942 45670
rect 10966 45668 11022 45670
rect 11046 45668 11102 45670
rect 11126 45668 11182 45670
rect 10886 44634 10942 44636
rect 10966 44634 11022 44636
rect 11046 44634 11102 44636
rect 11126 44634 11182 44636
rect 10886 44582 10932 44634
rect 10932 44582 10942 44634
rect 10966 44582 10996 44634
rect 10996 44582 11008 44634
rect 11008 44582 11022 44634
rect 11046 44582 11060 44634
rect 11060 44582 11072 44634
rect 11072 44582 11102 44634
rect 11126 44582 11136 44634
rect 11136 44582 11182 44634
rect 10886 44580 10942 44582
rect 10966 44580 11022 44582
rect 11046 44580 11102 44582
rect 11126 44580 11182 44582
rect 11610 44240 11666 44296
rect 10886 43546 10942 43548
rect 10966 43546 11022 43548
rect 11046 43546 11102 43548
rect 11126 43546 11182 43548
rect 10886 43494 10932 43546
rect 10932 43494 10942 43546
rect 10966 43494 10996 43546
rect 10996 43494 11008 43546
rect 11008 43494 11022 43546
rect 11046 43494 11060 43546
rect 11060 43494 11072 43546
rect 11072 43494 11102 43546
rect 11126 43494 11136 43546
rect 11136 43494 11182 43546
rect 10886 43492 10942 43494
rect 10966 43492 11022 43494
rect 11046 43492 11102 43494
rect 11126 43492 11182 43494
rect 10886 42458 10942 42460
rect 10966 42458 11022 42460
rect 11046 42458 11102 42460
rect 11126 42458 11182 42460
rect 10886 42406 10932 42458
rect 10932 42406 10942 42458
rect 10966 42406 10996 42458
rect 10996 42406 11008 42458
rect 11008 42406 11022 42458
rect 11046 42406 11060 42458
rect 11060 42406 11072 42458
rect 11072 42406 11102 42458
rect 11126 42406 11136 42458
rect 11136 42406 11182 42458
rect 10886 42404 10942 42406
rect 10966 42404 11022 42406
rect 11046 42404 11102 42406
rect 11126 42404 11182 42406
rect 12346 44376 12402 44432
rect 12898 44376 12954 44432
rect 10886 41370 10942 41372
rect 10966 41370 11022 41372
rect 11046 41370 11102 41372
rect 11126 41370 11182 41372
rect 10886 41318 10932 41370
rect 10932 41318 10942 41370
rect 10966 41318 10996 41370
rect 10996 41318 11008 41370
rect 11008 41318 11022 41370
rect 11046 41318 11060 41370
rect 11060 41318 11072 41370
rect 11072 41318 11102 41370
rect 11126 41318 11136 41370
rect 11136 41318 11182 41370
rect 10886 41316 10942 41318
rect 10966 41316 11022 41318
rect 11046 41316 11102 41318
rect 11126 41316 11182 41318
rect 10886 40282 10942 40284
rect 10966 40282 11022 40284
rect 11046 40282 11102 40284
rect 11126 40282 11182 40284
rect 10886 40230 10932 40282
rect 10932 40230 10942 40282
rect 10966 40230 10996 40282
rect 10996 40230 11008 40282
rect 11008 40230 11022 40282
rect 11046 40230 11060 40282
rect 11060 40230 11072 40282
rect 11072 40230 11102 40282
rect 11126 40230 11136 40282
rect 11136 40230 11182 40282
rect 10886 40228 10942 40230
rect 10966 40228 11022 40230
rect 11046 40228 11102 40230
rect 11126 40228 11182 40230
rect 10886 39194 10942 39196
rect 10966 39194 11022 39196
rect 11046 39194 11102 39196
rect 11126 39194 11182 39196
rect 10886 39142 10932 39194
rect 10932 39142 10942 39194
rect 10966 39142 10996 39194
rect 10996 39142 11008 39194
rect 11008 39142 11022 39194
rect 11046 39142 11060 39194
rect 11060 39142 11072 39194
rect 11072 39142 11102 39194
rect 11126 39142 11136 39194
rect 11136 39142 11182 39194
rect 10886 39140 10942 39142
rect 10966 39140 11022 39142
rect 11046 39140 11102 39142
rect 11126 39140 11182 39142
rect 10886 38106 10942 38108
rect 10966 38106 11022 38108
rect 11046 38106 11102 38108
rect 11126 38106 11182 38108
rect 10886 38054 10932 38106
rect 10932 38054 10942 38106
rect 10966 38054 10996 38106
rect 10996 38054 11008 38106
rect 11008 38054 11022 38106
rect 11046 38054 11060 38106
rect 11060 38054 11072 38106
rect 11072 38054 11102 38106
rect 11126 38054 11136 38106
rect 11136 38054 11182 38106
rect 10886 38052 10942 38054
rect 10966 38052 11022 38054
rect 11046 38052 11102 38054
rect 11126 38052 11182 38054
rect 10886 37018 10942 37020
rect 10966 37018 11022 37020
rect 11046 37018 11102 37020
rect 11126 37018 11182 37020
rect 10886 36966 10932 37018
rect 10932 36966 10942 37018
rect 10966 36966 10996 37018
rect 10996 36966 11008 37018
rect 11008 36966 11022 37018
rect 11046 36966 11060 37018
rect 11060 36966 11072 37018
rect 11072 36966 11102 37018
rect 11126 36966 11136 37018
rect 11136 36966 11182 37018
rect 10886 36964 10942 36966
rect 10966 36964 11022 36966
rect 11046 36964 11102 36966
rect 11126 36964 11182 36966
rect 10886 35930 10942 35932
rect 10966 35930 11022 35932
rect 11046 35930 11102 35932
rect 11126 35930 11182 35932
rect 10886 35878 10932 35930
rect 10932 35878 10942 35930
rect 10966 35878 10996 35930
rect 10996 35878 11008 35930
rect 11008 35878 11022 35930
rect 11046 35878 11060 35930
rect 11060 35878 11072 35930
rect 11072 35878 11102 35930
rect 11126 35878 11136 35930
rect 11136 35878 11182 35930
rect 10886 35876 10942 35878
rect 10966 35876 11022 35878
rect 11046 35876 11102 35878
rect 11126 35876 11182 35878
rect 10886 34842 10942 34844
rect 10966 34842 11022 34844
rect 11046 34842 11102 34844
rect 11126 34842 11182 34844
rect 10886 34790 10932 34842
rect 10932 34790 10942 34842
rect 10966 34790 10996 34842
rect 10996 34790 11008 34842
rect 11008 34790 11022 34842
rect 11046 34790 11060 34842
rect 11060 34790 11072 34842
rect 11072 34790 11102 34842
rect 11126 34790 11136 34842
rect 11136 34790 11182 34842
rect 10886 34788 10942 34790
rect 10966 34788 11022 34790
rect 11046 34788 11102 34790
rect 11126 34788 11182 34790
rect 10886 33754 10942 33756
rect 10966 33754 11022 33756
rect 11046 33754 11102 33756
rect 11126 33754 11182 33756
rect 10886 33702 10932 33754
rect 10932 33702 10942 33754
rect 10966 33702 10996 33754
rect 10996 33702 11008 33754
rect 11008 33702 11022 33754
rect 11046 33702 11060 33754
rect 11060 33702 11072 33754
rect 11072 33702 11102 33754
rect 11126 33702 11136 33754
rect 11136 33702 11182 33754
rect 10886 33700 10942 33702
rect 10966 33700 11022 33702
rect 11046 33700 11102 33702
rect 11126 33700 11182 33702
rect 10886 32666 10942 32668
rect 10966 32666 11022 32668
rect 11046 32666 11102 32668
rect 11126 32666 11182 32668
rect 10886 32614 10932 32666
rect 10932 32614 10942 32666
rect 10966 32614 10996 32666
rect 10996 32614 11008 32666
rect 11008 32614 11022 32666
rect 11046 32614 11060 32666
rect 11060 32614 11072 32666
rect 11072 32614 11102 32666
rect 11126 32614 11136 32666
rect 11136 32614 11182 32666
rect 10886 32612 10942 32614
rect 10966 32612 11022 32614
rect 11046 32612 11102 32614
rect 11126 32612 11182 32614
rect 10886 31578 10942 31580
rect 10966 31578 11022 31580
rect 11046 31578 11102 31580
rect 11126 31578 11182 31580
rect 10886 31526 10932 31578
rect 10932 31526 10942 31578
rect 10966 31526 10996 31578
rect 10996 31526 11008 31578
rect 11008 31526 11022 31578
rect 11046 31526 11060 31578
rect 11060 31526 11072 31578
rect 11072 31526 11102 31578
rect 11126 31526 11136 31578
rect 11136 31526 11182 31578
rect 10886 31524 10942 31526
rect 10966 31524 11022 31526
rect 11046 31524 11102 31526
rect 11126 31524 11182 31526
rect 13082 43732 13084 43752
rect 13084 43732 13136 43752
rect 13136 43732 13138 43752
rect 13082 43696 13138 43732
rect 12070 38664 12126 38720
rect 15852 70202 15908 70204
rect 15932 70202 15988 70204
rect 16012 70202 16068 70204
rect 16092 70202 16148 70204
rect 15852 70150 15898 70202
rect 15898 70150 15908 70202
rect 15932 70150 15962 70202
rect 15962 70150 15974 70202
rect 15974 70150 15988 70202
rect 16012 70150 16026 70202
rect 16026 70150 16038 70202
rect 16038 70150 16068 70202
rect 16092 70150 16102 70202
rect 16102 70150 16148 70202
rect 15852 70148 15908 70150
rect 15932 70148 15988 70150
rect 16012 70148 16068 70150
rect 16092 70148 16148 70150
rect 15852 69114 15908 69116
rect 15932 69114 15988 69116
rect 16012 69114 16068 69116
rect 16092 69114 16148 69116
rect 15852 69062 15898 69114
rect 15898 69062 15908 69114
rect 15932 69062 15962 69114
rect 15962 69062 15974 69114
rect 15974 69062 15988 69114
rect 16012 69062 16026 69114
rect 16026 69062 16038 69114
rect 16038 69062 16068 69114
rect 16092 69062 16102 69114
rect 16102 69062 16148 69114
rect 15852 69060 15908 69062
rect 15932 69060 15988 69062
rect 16012 69060 16068 69062
rect 16092 69060 16148 69062
rect 15852 68026 15908 68028
rect 15932 68026 15988 68028
rect 16012 68026 16068 68028
rect 16092 68026 16148 68028
rect 15852 67974 15898 68026
rect 15898 67974 15908 68026
rect 15932 67974 15962 68026
rect 15962 67974 15974 68026
rect 15974 67974 15988 68026
rect 16012 67974 16026 68026
rect 16026 67974 16038 68026
rect 16038 67974 16068 68026
rect 16092 67974 16102 68026
rect 16102 67974 16148 68026
rect 15852 67972 15908 67974
rect 15932 67972 15988 67974
rect 16012 67972 16068 67974
rect 16092 67972 16148 67974
rect 15852 66938 15908 66940
rect 15932 66938 15988 66940
rect 16012 66938 16068 66940
rect 16092 66938 16148 66940
rect 15852 66886 15898 66938
rect 15898 66886 15908 66938
rect 15932 66886 15962 66938
rect 15962 66886 15974 66938
rect 15974 66886 15988 66938
rect 16012 66886 16026 66938
rect 16026 66886 16038 66938
rect 16038 66886 16068 66938
rect 16092 66886 16102 66938
rect 16102 66886 16148 66938
rect 15852 66884 15908 66886
rect 15932 66884 15988 66886
rect 16012 66884 16068 66886
rect 16092 66884 16148 66886
rect 20817 75098 20873 75100
rect 20897 75098 20953 75100
rect 20977 75098 21033 75100
rect 21057 75098 21113 75100
rect 20817 75046 20863 75098
rect 20863 75046 20873 75098
rect 20897 75046 20927 75098
rect 20927 75046 20939 75098
rect 20939 75046 20953 75098
rect 20977 75046 20991 75098
rect 20991 75046 21003 75098
rect 21003 75046 21033 75098
rect 21057 75046 21067 75098
rect 21067 75046 21113 75098
rect 20817 75044 20873 75046
rect 20897 75044 20953 75046
rect 20977 75044 21033 75046
rect 21057 75044 21113 75046
rect 17406 73108 17408 73128
rect 17408 73108 17460 73128
rect 17460 73108 17462 73128
rect 17406 73072 17462 73108
rect 17498 71440 17554 71496
rect 15852 65850 15908 65852
rect 15932 65850 15988 65852
rect 16012 65850 16068 65852
rect 16092 65850 16148 65852
rect 15852 65798 15898 65850
rect 15898 65798 15908 65850
rect 15932 65798 15962 65850
rect 15962 65798 15974 65850
rect 15974 65798 15988 65850
rect 16012 65798 16026 65850
rect 16026 65798 16038 65850
rect 16038 65798 16068 65850
rect 16092 65798 16102 65850
rect 16102 65798 16148 65850
rect 15852 65796 15908 65798
rect 15932 65796 15988 65798
rect 16012 65796 16068 65798
rect 16092 65796 16148 65798
rect 14554 51312 14610 51368
rect 15852 64762 15908 64764
rect 15932 64762 15988 64764
rect 16012 64762 16068 64764
rect 16092 64762 16148 64764
rect 15852 64710 15898 64762
rect 15898 64710 15908 64762
rect 15932 64710 15962 64762
rect 15962 64710 15974 64762
rect 15974 64710 15988 64762
rect 16012 64710 16026 64762
rect 16026 64710 16038 64762
rect 16038 64710 16068 64762
rect 16092 64710 16102 64762
rect 16102 64710 16148 64762
rect 15852 64708 15908 64710
rect 15932 64708 15988 64710
rect 16012 64708 16068 64710
rect 16092 64708 16148 64710
rect 15852 63674 15908 63676
rect 15932 63674 15988 63676
rect 16012 63674 16068 63676
rect 16092 63674 16148 63676
rect 15852 63622 15898 63674
rect 15898 63622 15908 63674
rect 15932 63622 15962 63674
rect 15962 63622 15974 63674
rect 15974 63622 15988 63674
rect 16012 63622 16026 63674
rect 16026 63622 16038 63674
rect 16038 63622 16068 63674
rect 16092 63622 16102 63674
rect 16102 63622 16148 63674
rect 15852 63620 15908 63622
rect 15932 63620 15988 63622
rect 16012 63620 16068 63622
rect 16092 63620 16148 63622
rect 15852 62586 15908 62588
rect 15932 62586 15988 62588
rect 16012 62586 16068 62588
rect 16092 62586 16148 62588
rect 15852 62534 15898 62586
rect 15898 62534 15908 62586
rect 15932 62534 15962 62586
rect 15962 62534 15974 62586
rect 15974 62534 15988 62586
rect 16012 62534 16026 62586
rect 16026 62534 16038 62586
rect 16038 62534 16068 62586
rect 16092 62534 16102 62586
rect 16102 62534 16148 62586
rect 15852 62532 15908 62534
rect 15932 62532 15988 62534
rect 16012 62532 16068 62534
rect 16092 62532 16148 62534
rect 18418 71476 18420 71496
rect 18420 71476 18472 71496
rect 18472 71476 18474 71496
rect 18418 71440 18474 71476
rect 18510 66136 18566 66192
rect 20817 74010 20873 74012
rect 20897 74010 20953 74012
rect 20977 74010 21033 74012
rect 21057 74010 21113 74012
rect 20817 73958 20863 74010
rect 20863 73958 20873 74010
rect 20897 73958 20927 74010
rect 20927 73958 20939 74010
rect 20939 73958 20953 74010
rect 20977 73958 20991 74010
rect 20991 73958 21003 74010
rect 21003 73958 21033 74010
rect 21057 73958 21067 74010
rect 21067 73958 21113 74010
rect 20817 73956 20873 73958
rect 20897 73956 20953 73958
rect 20977 73956 21033 73958
rect 21057 73956 21113 73958
rect 15852 61498 15908 61500
rect 15932 61498 15988 61500
rect 16012 61498 16068 61500
rect 16092 61498 16148 61500
rect 15852 61446 15898 61498
rect 15898 61446 15908 61498
rect 15932 61446 15962 61498
rect 15962 61446 15974 61498
rect 15974 61446 15988 61498
rect 16012 61446 16026 61498
rect 16026 61446 16038 61498
rect 16038 61446 16068 61498
rect 16092 61446 16102 61498
rect 16102 61446 16148 61498
rect 15852 61444 15908 61446
rect 15932 61444 15988 61446
rect 16012 61444 16068 61446
rect 16092 61444 16148 61446
rect 15106 51312 15162 51368
rect 15852 60410 15908 60412
rect 15932 60410 15988 60412
rect 16012 60410 16068 60412
rect 16092 60410 16148 60412
rect 15852 60358 15898 60410
rect 15898 60358 15908 60410
rect 15932 60358 15962 60410
rect 15962 60358 15974 60410
rect 15974 60358 15988 60410
rect 16012 60358 16026 60410
rect 16026 60358 16038 60410
rect 16038 60358 16068 60410
rect 16092 60358 16102 60410
rect 16102 60358 16148 60410
rect 15852 60356 15908 60358
rect 15932 60356 15988 60358
rect 16012 60356 16068 60358
rect 16092 60356 16148 60358
rect 15852 59322 15908 59324
rect 15932 59322 15988 59324
rect 16012 59322 16068 59324
rect 16092 59322 16148 59324
rect 15852 59270 15898 59322
rect 15898 59270 15908 59322
rect 15932 59270 15962 59322
rect 15962 59270 15974 59322
rect 15974 59270 15988 59322
rect 16012 59270 16026 59322
rect 16026 59270 16038 59322
rect 16038 59270 16068 59322
rect 16092 59270 16102 59322
rect 16102 59270 16148 59322
rect 15852 59268 15908 59270
rect 15932 59268 15988 59270
rect 16012 59268 16068 59270
rect 16092 59268 16148 59270
rect 15852 58234 15908 58236
rect 15932 58234 15988 58236
rect 16012 58234 16068 58236
rect 16092 58234 16148 58236
rect 15852 58182 15898 58234
rect 15898 58182 15908 58234
rect 15932 58182 15962 58234
rect 15962 58182 15974 58234
rect 15974 58182 15988 58234
rect 16012 58182 16026 58234
rect 16026 58182 16038 58234
rect 16038 58182 16068 58234
rect 16092 58182 16102 58234
rect 16102 58182 16148 58234
rect 15852 58180 15908 58182
rect 15932 58180 15988 58182
rect 16012 58180 16068 58182
rect 16092 58180 16148 58182
rect 10886 30490 10942 30492
rect 10966 30490 11022 30492
rect 11046 30490 11102 30492
rect 11126 30490 11182 30492
rect 10886 30438 10932 30490
rect 10932 30438 10942 30490
rect 10966 30438 10996 30490
rect 10996 30438 11008 30490
rect 11008 30438 11022 30490
rect 11046 30438 11060 30490
rect 11060 30438 11072 30490
rect 11072 30438 11102 30490
rect 11126 30438 11136 30490
rect 11136 30438 11182 30490
rect 10886 30436 10942 30438
rect 10966 30436 11022 30438
rect 11046 30436 11102 30438
rect 11126 30436 11182 30438
rect 14094 38664 14150 38720
rect 10886 29402 10942 29404
rect 10966 29402 11022 29404
rect 11046 29402 11102 29404
rect 11126 29402 11182 29404
rect 10886 29350 10932 29402
rect 10932 29350 10942 29402
rect 10966 29350 10996 29402
rect 10996 29350 11008 29402
rect 11008 29350 11022 29402
rect 11046 29350 11060 29402
rect 11060 29350 11072 29402
rect 11072 29350 11102 29402
rect 11126 29350 11136 29402
rect 11136 29350 11182 29402
rect 10886 29348 10942 29350
rect 10966 29348 11022 29350
rect 11046 29348 11102 29350
rect 11126 29348 11182 29350
rect 12622 29008 12678 29064
rect 10886 28314 10942 28316
rect 10966 28314 11022 28316
rect 11046 28314 11102 28316
rect 11126 28314 11182 28316
rect 10886 28262 10932 28314
rect 10932 28262 10942 28314
rect 10966 28262 10996 28314
rect 10996 28262 11008 28314
rect 11008 28262 11022 28314
rect 11046 28262 11060 28314
rect 11060 28262 11072 28314
rect 11072 28262 11102 28314
rect 11126 28262 11136 28314
rect 11136 28262 11182 28314
rect 10886 28260 10942 28262
rect 10966 28260 11022 28262
rect 11046 28260 11102 28262
rect 11126 28260 11182 28262
rect 10886 27226 10942 27228
rect 10966 27226 11022 27228
rect 11046 27226 11102 27228
rect 11126 27226 11182 27228
rect 10886 27174 10932 27226
rect 10932 27174 10942 27226
rect 10966 27174 10996 27226
rect 10996 27174 11008 27226
rect 11008 27174 11022 27226
rect 11046 27174 11060 27226
rect 11060 27174 11072 27226
rect 11072 27174 11102 27226
rect 11126 27174 11136 27226
rect 11136 27174 11182 27226
rect 10886 27172 10942 27174
rect 10966 27172 11022 27174
rect 11046 27172 11102 27174
rect 11126 27172 11182 27174
rect 10886 26138 10942 26140
rect 10966 26138 11022 26140
rect 11046 26138 11102 26140
rect 11126 26138 11182 26140
rect 10886 26086 10932 26138
rect 10932 26086 10942 26138
rect 10966 26086 10996 26138
rect 10996 26086 11008 26138
rect 11008 26086 11022 26138
rect 11046 26086 11060 26138
rect 11060 26086 11072 26138
rect 11072 26086 11102 26138
rect 11126 26086 11136 26138
rect 11136 26086 11182 26138
rect 10886 26084 10942 26086
rect 10966 26084 11022 26086
rect 11046 26084 11102 26086
rect 11126 26084 11182 26086
rect 10886 25050 10942 25052
rect 10966 25050 11022 25052
rect 11046 25050 11102 25052
rect 11126 25050 11182 25052
rect 10886 24998 10932 25050
rect 10932 24998 10942 25050
rect 10966 24998 10996 25050
rect 10996 24998 11008 25050
rect 11008 24998 11022 25050
rect 11046 24998 11060 25050
rect 11060 24998 11072 25050
rect 11072 24998 11102 25050
rect 11126 24998 11136 25050
rect 11136 24998 11182 25050
rect 10886 24996 10942 24998
rect 10966 24996 11022 24998
rect 11046 24996 11102 24998
rect 11126 24996 11182 24998
rect 10886 23962 10942 23964
rect 10966 23962 11022 23964
rect 11046 23962 11102 23964
rect 11126 23962 11182 23964
rect 10886 23910 10932 23962
rect 10932 23910 10942 23962
rect 10966 23910 10996 23962
rect 10996 23910 11008 23962
rect 11008 23910 11022 23962
rect 11046 23910 11060 23962
rect 11060 23910 11072 23962
rect 11072 23910 11102 23962
rect 11126 23910 11136 23962
rect 11136 23910 11182 23962
rect 10886 23908 10942 23910
rect 10966 23908 11022 23910
rect 11046 23908 11102 23910
rect 11126 23908 11182 23910
rect 10886 22874 10942 22876
rect 10966 22874 11022 22876
rect 11046 22874 11102 22876
rect 11126 22874 11182 22876
rect 10886 22822 10932 22874
rect 10932 22822 10942 22874
rect 10966 22822 10996 22874
rect 10996 22822 11008 22874
rect 11008 22822 11022 22874
rect 11046 22822 11060 22874
rect 11060 22822 11072 22874
rect 11072 22822 11102 22874
rect 11126 22822 11136 22874
rect 11136 22822 11182 22874
rect 10886 22820 10942 22822
rect 10966 22820 11022 22822
rect 11046 22820 11102 22822
rect 11126 22820 11182 22822
rect 10886 21786 10942 21788
rect 10966 21786 11022 21788
rect 11046 21786 11102 21788
rect 11126 21786 11182 21788
rect 10886 21734 10932 21786
rect 10932 21734 10942 21786
rect 10966 21734 10996 21786
rect 10996 21734 11008 21786
rect 11008 21734 11022 21786
rect 11046 21734 11060 21786
rect 11060 21734 11072 21786
rect 11072 21734 11102 21786
rect 11126 21734 11136 21786
rect 11136 21734 11182 21786
rect 10886 21732 10942 21734
rect 10966 21732 11022 21734
rect 11046 21732 11102 21734
rect 11126 21732 11182 21734
rect 12806 29008 12862 29064
rect 15852 57146 15908 57148
rect 15932 57146 15988 57148
rect 16012 57146 16068 57148
rect 16092 57146 16148 57148
rect 15852 57094 15898 57146
rect 15898 57094 15908 57146
rect 15932 57094 15962 57146
rect 15962 57094 15974 57146
rect 15974 57094 15988 57146
rect 16012 57094 16026 57146
rect 16026 57094 16038 57146
rect 16038 57094 16068 57146
rect 16092 57094 16102 57146
rect 16102 57094 16148 57146
rect 15852 57092 15908 57094
rect 15932 57092 15988 57094
rect 16012 57092 16068 57094
rect 16092 57092 16148 57094
rect 15852 56058 15908 56060
rect 15932 56058 15988 56060
rect 16012 56058 16068 56060
rect 16092 56058 16148 56060
rect 15852 56006 15898 56058
rect 15898 56006 15908 56058
rect 15932 56006 15962 56058
rect 15962 56006 15974 56058
rect 15974 56006 15988 56058
rect 16012 56006 16026 56058
rect 16026 56006 16038 56058
rect 16038 56006 16068 56058
rect 16092 56006 16102 56058
rect 16102 56006 16148 56058
rect 15852 56004 15908 56006
rect 15932 56004 15988 56006
rect 16012 56004 16068 56006
rect 16092 56004 16148 56006
rect 15852 54970 15908 54972
rect 15932 54970 15988 54972
rect 16012 54970 16068 54972
rect 16092 54970 16148 54972
rect 15852 54918 15898 54970
rect 15898 54918 15908 54970
rect 15932 54918 15962 54970
rect 15962 54918 15974 54970
rect 15974 54918 15988 54970
rect 16012 54918 16026 54970
rect 16026 54918 16038 54970
rect 16038 54918 16068 54970
rect 16092 54918 16102 54970
rect 16102 54918 16148 54970
rect 15852 54916 15908 54918
rect 15932 54916 15988 54918
rect 16012 54916 16068 54918
rect 16092 54916 16148 54918
rect 15852 53882 15908 53884
rect 15932 53882 15988 53884
rect 16012 53882 16068 53884
rect 16092 53882 16148 53884
rect 15852 53830 15898 53882
rect 15898 53830 15908 53882
rect 15932 53830 15962 53882
rect 15962 53830 15974 53882
rect 15974 53830 15988 53882
rect 16012 53830 16026 53882
rect 16026 53830 16038 53882
rect 16038 53830 16068 53882
rect 16092 53830 16102 53882
rect 16102 53830 16148 53882
rect 15852 53828 15908 53830
rect 15932 53828 15988 53830
rect 16012 53828 16068 53830
rect 16092 53828 16148 53830
rect 15852 52794 15908 52796
rect 15932 52794 15988 52796
rect 16012 52794 16068 52796
rect 16092 52794 16148 52796
rect 15852 52742 15898 52794
rect 15898 52742 15908 52794
rect 15932 52742 15962 52794
rect 15962 52742 15974 52794
rect 15974 52742 15988 52794
rect 16012 52742 16026 52794
rect 16026 52742 16038 52794
rect 16038 52742 16068 52794
rect 16092 52742 16102 52794
rect 16102 52742 16148 52794
rect 15852 52740 15908 52742
rect 15932 52740 15988 52742
rect 16012 52740 16068 52742
rect 16092 52740 16148 52742
rect 17314 62328 17370 62384
rect 15852 51706 15908 51708
rect 15932 51706 15988 51708
rect 16012 51706 16068 51708
rect 16092 51706 16148 51708
rect 15852 51654 15898 51706
rect 15898 51654 15908 51706
rect 15932 51654 15962 51706
rect 15962 51654 15974 51706
rect 15974 51654 15988 51706
rect 16012 51654 16026 51706
rect 16026 51654 16038 51706
rect 16038 51654 16068 51706
rect 16092 51654 16102 51706
rect 16102 51654 16148 51706
rect 15852 51652 15908 51654
rect 15932 51652 15988 51654
rect 16012 51652 16068 51654
rect 16092 51652 16148 51654
rect 15852 50618 15908 50620
rect 15932 50618 15988 50620
rect 16012 50618 16068 50620
rect 16092 50618 16148 50620
rect 15852 50566 15898 50618
rect 15898 50566 15908 50618
rect 15932 50566 15962 50618
rect 15962 50566 15974 50618
rect 15974 50566 15988 50618
rect 16012 50566 16026 50618
rect 16026 50566 16038 50618
rect 16038 50566 16068 50618
rect 16092 50566 16102 50618
rect 16102 50566 16148 50618
rect 15852 50564 15908 50566
rect 15932 50564 15988 50566
rect 16012 50564 16068 50566
rect 16092 50564 16148 50566
rect 15852 49530 15908 49532
rect 15932 49530 15988 49532
rect 16012 49530 16068 49532
rect 16092 49530 16148 49532
rect 15852 49478 15898 49530
rect 15898 49478 15908 49530
rect 15932 49478 15962 49530
rect 15962 49478 15974 49530
rect 15974 49478 15988 49530
rect 16012 49478 16026 49530
rect 16026 49478 16038 49530
rect 16038 49478 16068 49530
rect 16092 49478 16102 49530
rect 16102 49478 16148 49530
rect 15852 49476 15908 49478
rect 15932 49476 15988 49478
rect 16012 49476 16068 49478
rect 16092 49476 16148 49478
rect 15852 48442 15908 48444
rect 15932 48442 15988 48444
rect 16012 48442 16068 48444
rect 16092 48442 16148 48444
rect 15852 48390 15898 48442
rect 15898 48390 15908 48442
rect 15932 48390 15962 48442
rect 15962 48390 15974 48442
rect 15974 48390 15988 48442
rect 16012 48390 16026 48442
rect 16026 48390 16038 48442
rect 16038 48390 16068 48442
rect 16092 48390 16102 48442
rect 16102 48390 16148 48442
rect 15852 48388 15908 48390
rect 15932 48388 15988 48390
rect 16012 48388 16068 48390
rect 16092 48388 16148 48390
rect 15852 47354 15908 47356
rect 15932 47354 15988 47356
rect 16012 47354 16068 47356
rect 16092 47354 16148 47356
rect 15852 47302 15898 47354
rect 15898 47302 15908 47354
rect 15932 47302 15962 47354
rect 15962 47302 15974 47354
rect 15974 47302 15988 47354
rect 16012 47302 16026 47354
rect 16026 47302 16038 47354
rect 16038 47302 16068 47354
rect 16092 47302 16102 47354
rect 16102 47302 16148 47354
rect 15852 47300 15908 47302
rect 15932 47300 15988 47302
rect 16012 47300 16068 47302
rect 16092 47300 16148 47302
rect 15852 46266 15908 46268
rect 15932 46266 15988 46268
rect 16012 46266 16068 46268
rect 16092 46266 16148 46268
rect 15852 46214 15898 46266
rect 15898 46214 15908 46266
rect 15932 46214 15962 46266
rect 15962 46214 15974 46266
rect 15974 46214 15988 46266
rect 16012 46214 16026 46266
rect 16026 46214 16038 46266
rect 16038 46214 16068 46266
rect 16092 46214 16102 46266
rect 16102 46214 16148 46266
rect 15852 46212 15908 46214
rect 15932 46212 15988 46214
rect 16012 46212 16068 46214
rect 16092 46212 16148 46214
rect 15852 45178 15908 45180
rect 15932 45178 15988 45180
rect 16012 45178 16068 45180
rect 16092 45178 16148 45180
rect 15852 45126 15898 45178
rect 15898 45126 15908 45178
rect 15932 45126 15962 45178
rect 15962 45126 15974 45178
rect 15974 45126 15988 45178
rect 16012 45126 16026 45178
rect 16026 45126 16038 45178
rect 16038 45126 16068 45178
rect 16092 45126 16102 45178
rect 16102 45126 16148 45178
rect 15852 45124 15908 45126
rect 15932 45124 15988 45126
rect 16012 45124 16068 45126
rect 16092 45124 16148 45126
rect 15852 44090 15908 44092
rect 15932 44090 15988 44092
rect 16012 44090 16068 44092
rect 16092 44090 16148 44092
rect 15852 44038 15898 44090
rect 15898 44038 15908 44090
rect 15932 44038 15962 44090
rect 15962 44038 15974 44090
rect 15974 44038 15988 44090
rect 16012 44038 16026 44090
rect 16026 44038 16038 44090
rect 16038 44038 16068 44090
rect 16092 44038 16102 44090
rect 16102 44038 16148 44090
rect 15852 44036 15908 44038
rect 15932 44036 15988 44038
rect 16012 44036 16068 44038
rect 16092 44036 16148 44038
rect 16854 47776 16910 47832
rect 15852 43002 15908 43004
rect 15932 43002 15988 43004
rect 16012 43002 16068 43004
rect 16092 43002 16148 43004
rect 15852 42950 15898 43002
rect 15898 42950 15908 43002
rect 15932 42950 15962 43002
rect 15962 42950 15974 43002
rect 15974 42950 15988 43002
rect 16012 42950 16026 43002
rect 16026 42950 16038 43002
rect 16038 42950 16068 43002
rect 16092 42950 16102 43002
rect 16102 42950 16148 43002
rect 15852 42948 15908 42950
rect 15932 42948 15988 42950
rect 16012 42948 16068 42950
rect 16092 42948 16148 42950
rect 15852 41914 15908 41916
rect 15932 41914 15988 41916
rect 16012 41914 16068 41916
rect 16092 41914 16148 41916
rect 15852 41862 15898 41914
rect 15898 41862 15908 41914
rect 15932 41862 15962 41914
rect 15962 41862 15974 41914
rect 15974 41862 15988 41914
rect 16012 41862 16026 41914
rect 16026 41862 16038 41914
rect 16038 41862 16068 41914
rect 16092 41862 16102 41914
rect 16102 41862 16148 41914
rect 15852 41860 15908 41862
rect 15932 41860 15988 41862
rect 16012 41860 16068 41862
rect 16092 41860 16148 41862
rect 15852 40826 15908 40828
rect 15932 40826 15988 40828
rect 16012 40826 16068 40828
rect 16092 40826 16148 40828
rect 15852 40774 15898 40826
rect 15898 40774 15908 40826
rect 15932 40774 15962 40826
rect 15962 40774 15974 40826
rect 15974 40774 15988 40826
rect 16012 40774 16026 40826
rect 16026 40774 16038 40826
rect 16038 40774 16068 40826
rect 16092 40774 16102 40826
rect 16102 40774 16148 40826
rect 15852 40772 15908 40774
rect 15932 40772 15988 40774
rect 16012 40772 16068 40774
rect 16092 40772 16148 40774
rect 15382 36896 15438 36952
rect 13634 28736 13690 28792
rect 14738 28736 14794 28792
rect 14370 28192 14426 28248
rect 15852 39738 15908 39740
rect 15932 39738 15988 39740
rect 16012 39738 16068 39740
rect 16092 39738 16148 39740
rect 15852 39686 15898 39738
rect 15898 39686 15908 39738
rect 15932 39686 15962 39738
rect 15962 39686 15974 39738
rect 15974 39686 15988 39738
rect 16012 39686 16026 39738
rect 16026 39686 16038 39738
rect 16038 39686 16068 39738
rect 16092 39686 16102 39738
rect 16102 39686 16148 39738
rect 15852 39684 15908 39686
rect 15932 39684 15988 39686
rect 16012 39684 16068 39686
rect 16092 39684 16148 39686
rect 15852 38650 15908 38652
rect 15932 38650 15988 38652
rect 16012 38650 16068 38652
rect 16092 38650 16148 38652
rect 15852 38598 15898 38650
rect 15898 38598 15908 38650
rect 15932 38598 15962 38650
rect 15962 38598 15974 38650
rect 15974 38598 15988 38650
rect 16012 38598 16026 38650
rect 16026 38598 16038 38650
rect 16038 38598 16068 38650
rect 16092 38598 16102 38650
rect 16102 38598 16148 38650
rect 15852 38596 15908 38598
rect 15932 38596 15988 38598
rect 16012 38596 16068 38598
rect 16092 38596 16148 38598
rect 15852 37562 15908 37564
rect 15932 37562 15988 37564
rect 16012 37562 16068 37564
rect 16092 37562 16148 37564
rect 15852 37510 15898 37562
rect 15898 37510 15908 37562
rect 15932 37510 15962 37562
rect 15962 37510 15974 37562
rect 15974 37510 15988 37562
rect 16012 37510 16026 37562
rect 16026 37510 16038 37562
rect 16038 37510 16068 37562
rect 16092 37510 16102 37562
rect 16102 37510 16148 37562
rect 15852 37508 15908 37510
rect 15932 37508 15988 37510
rect 16012 37508 16068 37510
rect 16092 37508 16148 37510
rect 15934 36896 15990 36952
rect 25782 75642 25838 75644
rect 25862 75642 25918 75644
rect 25942 75642 25998 75644
rect 26022 75642 26078 75644
rect 25782 75590 25828 75642
rect 25828 75590 25838 75642
rect 25862 75590 25892 75642
rect 25892 75590 25904 75642
rect 25904 75590 25918 75642
rect 25942 75590 25956 75642
rect 25956 75590 25968 75642
rect 25968 75590 25998 75642
rect 26022 75590 26032 75642
rect 26032 75590 26078 75642
rect 25782 75588 25838 75590
rect 25862 75588 25918 75590
rect 25942 75588 25998 75590
rect 26022 75588 26078 75590
rect 20817 72922 20873 72924
rect 20897 72922 20953 72924
rect 20977 72922 21033 72924
rect 21057 72922 21113 72924
rect 20817 72870 20863 72922
rect 20863 72870 20873 72922
rect 20897 72870 20927 72922
rect 20927 72870 20939 72922
rect 20939 72870 20953 72922
rect 20977 72870 20991 72922
rect 20991 72870 21003 72922
rect 21003 72870 21033 72922
rect 21057 72870 21067 72922
rect 21067 72870 21113 72922
rect 20817 72868 20873 72870
rect 20897 72868 20953 72870
rect 20977 72868 21033 72870
rect 21057 72868 21113 72870
rect 20817 71834 20873 71836
rect 20897 71834 20953 71836
rect 20977 71834 21033 71836
rect 21057 71834 21113 71836
rect 20817 71782 20863 71834
rect 20863 71782 20873 71834
rect 20897 71782 20927 71834
rect 20927 71782 20939 71834
rect 20939 71782 20953 71834
rect 20977 71782 20991 71834
rect 20991 71782 21003 71834
rect 21003 71782 21033 71834
rect 21057 71782 21067 71834
rect 21067 71782 21113 71834
rect 20817 71780 20873 71782
rect 20897 71780 20953 71782
rect 20977 71780 21033 71782
rect 21057 71780 21113 71782
rect 20442 68856 20498 68912
rect 20442 68312 20498 68368
rect 18970 61104 19026 61160
rect 20817 70746 20873 70748
rect 20897 70746 20953 70748
rect 20977 70746 21033 70748
rect 21057 70746 21113 70748
rect 20817 70694 20863 70746
rect 20863 70694 20873 70746
rect 20897 70694 20927 70746
rect 20927 70694 20939 70746
rect 20939 70694 20953 70746
rect 20977 70694 20991 70746
rect 20991 70694 21003 70746
rect 21003 70694 21033 70746
rect 21057 70694 21067 70746
rect 21067 70694 21113 70746
rect 20817 70692 20873 70694
rect 20897 70692 20953 70694
rect 20977 70692 21033 70694
rect 21057 70692 21113 70694
rect 20817 69658 20873 69660
rect 20897 69658 20953 69660
rect 20977 69658 21033 69660
rect 21057 69658 21113 69660
rect 20817 69606 20863 69658
rect 20863 69606 20873 69658
rect 20897 69606 20927 69658
rect 20927 69606 20939 69658
rect 20939 69606 20953 69658
rect 20977 69606 20991 69658
rect 20991 69606 21003 69658
rect 21003 69606 21033 69658
rect 21057 69606 21067 69658
rect 21067 69606 21113 69658
rect 20817 69604 20873 69606
rect 20897 69604 20953 69606
rect 20977 69604 21033 69606
rect 21057 69604 21113 69606
rect 20817 68570 20873 68572
rect 20897 68570 20953 68572
rect 20977 68570 21033 68572
rect 21057 68570 21113 68572
rect 20817 68518 20863 68570
rect 20863 68518 20873 68570
rect 20897 68518 20927 68570
rect 20927 68518 20939 68570
rect 20939 68518 20953 68570
rect 20977 68518 20991 68570
rect 20991 68518 21003 68570
rect 21003 68518 21033 68570
rect 21057 68518 21067 68570
rect 21067 68518 21113 68570
rect 20817 68516 20873 68518
rect 20897 68516 20953 68518
rect 20977 68516 21033 68518
rect 21057 68516 21113 68518
rect 20817 67482 20873 67484
rect 20897 67482 20953 67484
rect 20977 67482 21033 67484
rect 21057 67482 21113 67484
rect 20817 67430 20863 67482
rect 20863 67430 20873 67482
rect 20897 67430 20927 67482
rect 20927 67430 20939 67482
rect 20939 67430 20953 67482
rect 20977 67430 20991 67482
rect 20991 67430 21003 67482
rect 21003 67430 21033 67482
rect 21057 67430 21067 67482
rect 21067 67430 21113 67482
rect 20817 67428 20873 67430
rect 20897 67428 20953 67430
rect 20977 67428 21033 67430
rect 21057 67428 21113 67430
rect 20817 66394 20873 66396
rect 20897 66394 20953 66396
rect 20977 66394 21033 66396
rect 21057 66394 21113 66396
rect 20817 66342 20863 66394
rect 20863 66342 20873 66394
rect 20897 66342 20927 66394
rect 20927 66342 20939 66394
rect 20939 66342 20953 66394
rect 20977 66342 20991 66394
rect 20991 66342 21003 66394
rect 21003 66342 21033 66394
rect 21057 66342 21067 66394
rect 21067 66342 21113 66394
rect 20817 66340 20873 66342
rect 20897 66340 20953 66342
rect 20977 66340 21033 66342
rect 21057 66340 21113 66342
rect 20817 65306 20873 65308
rect 20897 65306 20953 65308
rect 20977 65306 21033 65308
rect 21057 65306 21113 65308
rect 20817 65254 20863 65306
rect 20863 65254 20873 65306
rect 20897 65254 20927 65306
rect 20927 65254 20939 65306
rect 20939 65254 20953 65306
rect 20977 65254 20991 65306
rect 20991 65254 21003 65306
rect 21003 65254 21033 65306
rect 21057 65254 21067 65306
rect 21067 65254 21113 65306
rect 20817 65252 20873 65254
rect 20897 65252 20953 65254
rect 20977 65252 21033 65254
rect 21057 65252 21113 65254
rect 20817 64218 20873 64220
rect 20897 64218 20953 64220
rect 20977 64218 21033 64220
rect 21057 64218 21113 64220
rect 20817 64166 20863 64218
rect 20863 64166 20873 64218
rect 20897 64166 20927 64218
rect 20927 64166 20939 64218
rect 20939 64166 20953 64218
rect 20977 64166 20991 64218
rect 20991 64166 21003 64218
rect 21003 64166 21033 64218
rect 21057 64166 21067 64218
rect 21067 64166 21113 64218
rect 20817 64164 20873 64166
rect 20897 64164 20953 64166
rect 20977 64164 21033 64166
rect 21057 64164 21113 64166
rect 18970 60036 19026 60072
rect 18970 60016 18972 60036
rect 18972 60016 19024 60036
rect 19024 60016 19026 60036
rect 19338 60172 19394 60208
rect 19338 60152 19340 60172
rect 19340 60152 19392 60172
rect 19392 60152 19394 60172
rect 15842 36624 15898 36680
rect 15852 36474 15908 36476
rect 15932 36474 15988 36476
rect 16012 36474 16068 36476
rect 16092 36474 16148 36476
rect 15852 36422 15898 36474
rect 15898 36422 15908 36474
rect 15932 36422 15962 36474
rect 15962 36422 15974 36474
rect 15974 36422 15988 36474
rect 16012 36422 16026 36474
rect 16026 36422 16038 36474
rect 16038 36422 16068 36474
rect 16092 36422 16102 36474
rect 16102 36422 16148 36474
rect 15852 36420 15908 36422
rect 15932 36420 15988 36422
rect 16012 36420 16068 36422
rect 16092 36420 16148 36422
rect 15852 35386 15908 35388
rect 15932 35386 15988 35388
rect 16012 35386 16068 35388
rect 16092 35386 16148 35388
rect 15852 35334 15898 35386
rect 15898 35334 15908 35386
rect 15932 35334 15962 35386
rect 15962 35334 15974 35386
rect 15974 35334 15988 35386
rect 16012 35334 16026 35386
rect 16026 35334 16038 35386
rect 16038 35334 16068 35386
rect 16092 35334 16102 35386
rect 16102 35334 16148 35386
rect 15852 35332 15908 35334
rect 15932 35332 15988 35334
rect 16012 35332 16068 35334
rect 16092 35332 16148 35334
rect 15852 34298 15908 34300
rect 15932 34298 15988 34300
rect 16012 34298 16068 34300
rect 16092 34298 16148 34300
rect 15852 34246 15898 34298
rect 15898 34246 15908 34298
rect 15932 34246 15962 34298
rect 15962 34246 15974 34298
rect 15974 34246 15988 34298
rect 16012 34246 16026 34298
rect 16026 34246 16038 34298
rect 16038 34246 16068 34298
rect 16092 34246 16102 34298
rect 16102 34246 16148 34298
rect 15852 34244 15908 34246
rect 15932 34244 15988 34246
rect 16012 34244 16068 34246
rect 16092 34244 16148 34246
rect 15852 33210 15908 33212
rect 15932 33210 15988 33212
rect 16012 33210 16068 33212
rect 16092 33210 16148 33212
rect 15852 33158 15898 33210
rect 15898 33158 15908 33210
rect 15932 33158 15962 33210
rect 15962 33158 15974 33210
rect 15974 33158 15988 33210
rect 16012 33158 16026 33210
rect 16026 33158 16038 33210
rect 16038 33158 16068 33210
rect 16092 33158 16102 33210
rect 16102 33158 16148 33210
rect 15852 33156 15908 33158
rect 15932 33156 15988 33158
rect 16012 33156 16068 33158
rect 16092 33156 16148 33158
rect 15474 27784 15530 27840
rect 15382 27512 15438 27568
rect 10886 20698 10942 20700
rect 10966 20698 11022 20700
rect 11046 20698 11102 20700
rect 11126 20698 11182 20700
rect 10886 20646 10932 20698
rect 10932 20646 10942 20698
rect 10966 20646 10996 20698
rect 10996 20646 11008 20698
rect 11008 20646 11022 20698
rect 11046 20646 11060 20698
rect 11060 20646 11072 20698
rect 11072 20646 11102 20698
rect 11126 20646 11136 20698
rect 11136 20646 11182 20698
rect 10886 20644 10942 20646
rect 10966 20644 11022 20646
rect 11046 20644 11102 20646
rect 11126 20644 11182 20646
rect 10886 19610 10942 19612
rect 10966 19610 11022 19612
rect 11046 19610 11102 19612
rect 11126 19610 11182 19612
rect 10886 19558 10932 19610
rect 10932 19558 10942 19610
rect 10966 19558 10996 19610
rect 10996 19558 11008 19610
rect 11008 19558 11022 19610
rect 11046 19558 11060 19610
rect 11060 19558 11072 19610
rect 11072 19558 11102 19610
rect 11126 19558 11136 19610
rect 11136 19558 11182 19610
rect 10886 19556 10942 19558
rect 10966 19556 11022 19558
rect 11046 19556 11102 19558
rect 11126 19556 11182 19558
rect 10886 18522 10942 18524
rect 10966 18522 11022 18524
rect 11046 18522 11102 18524
rect 11126 18522 11182 18524
rect 10886 18470 10932 18522
rect 10932 18470 10942 18522
rect 10966 18470 10996 18522
rect 10996 18470 11008 18522
rect 11008 18470 11022 18522
rect 11046 18470 11060 18522
rect 11060 18470 11072 18522
rect 11072 18470 11102 18522
rect 11126 18470 11136 18522
rect 11136 18470 11182 18522
rect 10886 18468 10942 18470
rect 10966 18468 11022 18470
rect 11046 18468 11102 18470
rect 11126 18468 11182 18470
rect 10886 17434 10942 17436
rect 10966 17434 11022 17436
rect 11046 17434 11102 17436
rect 11126 17434 11182 17436
rect 10886 17382 10932 17434
rect 10932 17382 10942 17434
rect 10966 17382 10996 17434
rect 10996 17382 11008 17434
rect 11008 17382 11022 17434
rect 11046 17382 11060 17434
rect 11060 17382 11072 17434
rect 11072 17382 11102 17434
rect 11126 17382 11136 17434
rect 11136 17382 11182 17434
rect 10886 17380 10942 17382
rect 10966 17380 11022 17382
rect 11046 17380 11102 17382
rect 11126 17380 11182 17382
rect 10886 16346 10942 16348
rect 10966 16346 11022 16348
rect 11046 16346 11102 16348
rect 11126 16346 11182 16348
rect 10886 16294 10932 16346
rect 10932 16294 10942 16346
rect 10966 16294 10996 16346
rect 10996 16294 11008 16346
rect 11008 16294 11022 16346
rect 11046 16294 11060 16346
rect 11060 16294 11072 16346
rect 11072 16294 11102 16346
rect 11126 16294 11136 16346
rect 11136 16294 11182 16346
rect 10886 16292 10942 16294
rect 10966 16292 11022 16294
rect 11046 16292 11102 16294
rect 11126 16292 11182 16294
rect 10886 15258 10942 15260
rect 10966 15258 11022 15260
rect 11046 15258 11102 15260
rect 11126 15258 11182 15260
rect 10886 15206 10932 15258
rect 10932 15206 10942 15258
rect 10966 15206 10996 15258
rect 10996 15206 11008 15258
rect 11008 15206 11022 15258
rect 11046 15206 11060 15258
rect 11060 15206 11072 15258
rect 11072 15206 11102 15258
rect 11126 15206 11136 15258
rect 11136 15206 11182 15258
rect 10886 15204 10942 15206
rect 10966 15204 11022 15206
rect 11046 15204 11102 15206
rect 11126 15204 11182 15206
rect 10886 14170 10942 14172
rect 10966 14170 11022 14172
rect 11046 14170 11102 14172
rect 11126 14170 11182 14172
rect 10886 14118 10932 14170
rect 10932 14118 10942 14170
rect 10966 14118 10996 14170
rect 10996 14118 11008 14170
rect 11008 14118 11022 14170
rect 11046 14118 11060 14170
rect 11060 14118 11072 14170
rect 11072 14118 11102 14170
rect 11126 14118 11136 14170
rect 11136 14118 11182 14170
rect 10886 14116 10942 14118
rect 10966 14116 11022 14118
rect 11046 14116 11102 14118
rect 11126 14116 11182 14118
rect 10886 13082 10942 13084
rect 10966 13082 11022 13084
rect 11046 13082 11102 13084
rect 11126 13082 11182 13084
rect 10886 13030 10932 13082
rect 10932 13030 10942 13082
rect 10966 13030 10996 13082
rect 10996 13030 11008 13082
rect 11008 13030 11022 13082
rect 11046 13030 11060 13082
rect 11060 13030 11072 13082
rect 11072 13030 11102 13082
rect 11126 13030 11136 13082
rect 11136 13030 11182 13082
rect 10886 13028 10942 13030
rect 10966 13028 11022 13030
rect 11046 13028 11102 13030
rect 11126 13028 11182 13030
rect 10886 11994 10942 11996
rect 10966 11994 11022 11996
rect 11046 11994 11102 11996
rect 11126 11994 11182 11996
rect 10886 11942 10932 11994
rect 10932 11942 10942 11994
rect 10966 11942 10996 11994
rect 10996 11942 11008 11994
rect 11008 11942 11022 11994
rect 11046 11942 11060 11994
rect 11060 11942 11072 11994
rect 11072 11942 11102 11994
rect 11126 11942 11136 11994
rect 11136 11942 11182 11994
rect 10886 11940 10942 11942
rect 10966 11940 11022 11942
rect 11046 11940 11102 11942
rect 11126 11940 11182 11942
rect 10886 10906 10942 10908
rect 10966 10906 11022 10908
rect 11046 10906 11102 10908
rect 11126 10906 11182 10908
rect 10886 10854 10932 10906
rect 10932 10854 10942 10906
rect 10966 10854 10996 10906
rect 10996 10854 11008 10906
rect 11008 10854 11022 10906
rect 11046 10854 11060 10906
rect 11060 10854 11072 10906
rect 11072 10854 11102 10906
rect 11126 10854 11136 10906
rect 11136 10854 11182 10906
rect 10886 10852 10942 10854
rect 10966 10852 11022 10854
rect 11046 10852 11102 10854
rect 11126 10852 11182 10854
rect 10886 9818 10942 9820
rect 10966 9818 11022 9820
rect 11046 9818 11102 9820
rect 11126 9818 11182 9820
rect 10886 9766 10932 9818
rect 10932 9766 10942 9818
rect 10966 9766 10996 9818
rect 10996 9766 11008 9818
rect 11008 9766 11022 9818
rect 11046 9766 11060 9818
rect 11060 9766 11072 9818
rect 11072 9766 11102 9818
rect 11126 9766 11136 9818
rect 11136 9766 11182 9818
rect 10886 9764 10942 9766
rect 10966 9764 11022 9766
rect 11046 9764 11102 9766
rect 11126 9764 11182 9766
rect 10886 8730 10942 8732
rect 10966 8730 11022 8732
rect 11046 8730 11102 8732
rect 11126 8730 11182 8732
rect 10886 8678 10932 8730
rect 10932 8678 10942 8730
rect 10966 8678 10996 8730
rect 10996 8678 11008 8730
rect 11008 8678 11022 8730
rect 11046 8678 11060 8730
rect 11060 8678 11072 8730
rect 11072 8678 11102 8730
rect 11126 8678 11136 8730
rect 11136 8678 11182 8730
rect 10886 8676 10942 8678
rect 10966 8676 11022 8678
rect 11046 8676 11102 8678
rect 11126 8676 11182 8678
rect 15852 32122 15908 32124
rect 15932 32122 15988 32124
rect 16012 32122 16068 32124
rect 16092 32122 16148 32124
rect 15852 32070 15898 32122
rect 15898 32070 15908 32122
rect 15932 32070 15962 32122
rect 15962 32070 15974 32122
rect 15974 32070 15988 32122
rect 16012 32070 16026 32122
rect 16026 32070 16038 32122
rect 16038 32070 16068 32122
rect 16092 32070 16102 32122
rect 16102 32070 16148 32122
rect 15852 32068 15908 32070
rect 15932 32068 15988 32070
rect 16012 32068 16068 32070
rect 16092 32068 16148 32070
rect 15852 31034 15908 31036
rect 15932 31034 15988 31036
rect 16012 31034 16068 31036
rect 16092 31034 16148 31036
rect 15852 30982 15898 31034
rect 15898 30982 15908 31034
rect 15932 30982 15962 31034
rect 15962 30982 15974 31034
rect 15974 30982 15988 31034
rect 16012 30982 16026 31034
rect 16026 30982 16038 31034
rect 16038 30982 16068 31034
rect 16092 30982 16102 31034
rect 16102 30982 16148 31034
rect 15852 30980 15908 30982
rect 15932 30980 15988 30982
rect 16012 30980 16068 30982
rect 16092 30980 16148 30982
rect 15852 29946 15908 29948
rect 15932 29946 15988 29948
rect 16012 29946 16068 29948
rect 16092 29946 16148 29948
rect 15852 29894 15898 29946
rect 15898 29894 15908 29946
rect 15932 29894 15962 29946
rect 15962 29894 15974 29946
rect 15974 29894 15988 29946
rect 16012 29894 16026 29946
rect 16026 29894 16038 29946
rect 16038 29894 16068 29946
rect 16092 29894 16102 29946
rect 16102 29894 16148 29946
rect 15852 29892 15908 29894
rect 15932 29892 15988 29894
rect 16012 29892 16068 29894
rect 16092 29892 16148 29894
rect 15852 28858 15908 28860
rect 15932 28858 15988 28860
rect 16012 28858 16068 28860
rect 16092 28858 16148 28860
rect 15852 28806 15898 28858
rect 15898 28806 15908 28858
rect 15932 28806 15962 28858
rect 15962 28806 15974 28858
rect 15974 28806 15988 28858
rect 16012 28806 16026 28858
rect 16026 28806 16038 28858
rect 16038 28806 16068 28858
rect 16092 28806 16102 28858
rect 16102 28806 16148 28858
rect 15852 28804 15908 28806
rect 15932 28804 15988 28806
rect 16012 28804 16068 28806
rect 16092 28804 16148 28806
rect 15842 28212 15898 28248
rect 15842 28192 15844 28212
rect 15844 28192 15896 28212
rect 15896 28192 15898 28212
rect 15750 28056 15806 28112
rect 15852 27770 15908 27772
rect 15932 27770 15988 27772
rect 16012 27770 16068 27772
rect 16092 27770 16148 27772
rect 15852 27718 15898 27770
rect 15898 27718 15908 27770
rect 15932 27718 15962 27770
rect 15962 27718 15974 27770
rect 15974 27718 15988 27770
rect 16012 27718 16026 27770
rect 16026 27718 16038 27770
rect 16038 27718 16068 27770
rect 16092 27718 16102 27770
rect 16102 27718 16148 27770
rect 15852 27716 15908 27718
rect 15932 27716 15988 27718
rect 16012 27716 16068 27718
rect 16092 27716 16148 27718
rect 16210 26968 16266 27024
rect 15852 26682 15908 26684
rect 15932 26682 15988 26684
rect 16012 26682 16068 26684
rect 16092 26682 16148 26684
rect 15852 26630 15898 26682
rect 15898 26630 15908 26682
rect 15932 26630 15962 26682
rect 15962 26630 15974 26682
rect 15974 26630 15988 26682
rect 16012 26630 16026 26682
rect 16026 26630 16038 26682
rect 16038 26630 16068 26682
rect 16092 26630 16102 26682
rect 16102 26630 16148 26682
rect 15852 26628 15908 26630
rect 15932 26628 15988 26630
rect 16012 26628 16068 26630
rect 16092 26628 16148 26630
rect 15852 25594 15908 25596
rect 15932 25594 15988 25596
rect 16012 25594 16068 25596
rect 16092 25594 16148 25596
rect 15852 25542 15898 25594
rect 15898 25542 15908 25594
rect 15932 25542 15962 25594
rect 15962 25542 15974 25594
rect 15974 25542 15988 25594
rect 16012 25542 16026 25594
rect 16026 25542 16038 25594
rect 16038 25542 16068 25594
rect 16092 25542 16102 25594
rect 16102 25542 16148 25594
rect 15852 25540 15908 25542
rect 15932 25540 15988 25542
rect 16012 25540 16068 25542
rect 16092 25540 16148 25542
rect 15852 24506 15908 24508
rect 15932 24506 15988 24508
rect 16012 24506 16068 24508
rect 16092 24506 16148 24508
rect 15852 24454 15898 24506
rect 15898 24454 15908 24506
rect 15932 24454 15962 24506
rect 15962 24454 15974 24506
rect 15974 24454 15988 24506
rect 16012 24454 16026 24506
rect 16026 24454 16038 24506
rect 16038 24454 16068 24506
rect 16092 24454 16102 24506
rect 16102 24454 16148 24506
rect 15852 24452 15908 24454
rect 15932 24452 15988 24454
rect 16012 24452 16068 24454
rect 16092 24452 16148 24454
rect 15852 23418 15908 23420
rect 15932 23418 15988 23420
rect 16012 23418 16068 23420
rect 16092 23418 16148 23420
rect 15852 23366 15898 23418
rect 15898 23366 15908 23418
rect 15932 23366 15962 23418
rect 15962 23366 15974 23418
rect 15974 23366 15988 23418
rect 16012 23366 16026 23418
rect 16026 23366 16038 23418
rect 16038 23366 16068 23418
rect 16092 23366 16102 23418
rect 16102 23366 16148 23418
rect 15852 23364 15908 23366
rect 15932 23364 15988 23366
rect 16012 23364 16068 23366
rect 16092 23364 16148 23366
rect 15852 22330 15908 22332
rect 15932 22330 15988 22332
rect 16012 22330 16068 22332
rect 16092 22330 16148 22332
rect 15852 22278 15898 22330
rect 15898 22278 15908 22330
rect 15932 22278 15962 22330
rect 15962 22278 15974 22330
rect 15974 22278 15988 22330
rect 16012 22278 16026 22330
rect 16026 22278 16038 22330
rect 16038 22278 16068 22330
rect 16092 22278 16102 22330
rect 16102 22278 16148 22330
rect 15852 22276 15908 22278
rect 15932 22276 15988 22278
rect 16012 22276 16068 22278
rect 16092 22276 16148 22278
rect 15852 21242 15908 21244
rect 15932 21242 15988 21244
rect 16012 21242 16068 21244
rect 16092 21242 16148 21244
rect 15852 21190 15898 21242
rect 15898 21190 15908 21242
rect 15932 21190 15962 21242
rect 15962 21190 15974 21242
rect 15974 21190 15988 21242
rect 16012 21190 16026 21242
rect 16026 21190 16038 21242
rect 16038 21190 16068 21242
rect 16092 21190 16102 21242
rect 16102 21190 16148 21242
rect 15852 21188 15908 21190
rect 15932 21188 15988 21190
rect 16012 21188 16068 21190
rect 16092 21188 16148 21190
rect 15852 20154 15908 20156
rect 15932 20154 15988 20156
rect 16012 20154 16068 20156
rect 16092 20154 16148 20156
rect 15852 20102 15898 20154
rect 15898 20102 15908 20154
rect 15932 20102 15962 20154
rect 15962 20102 15974 20154
rect 15974 20102 15988 20154
rect 16012 20102 16026 20154
rect 16026 20102 16038 20154
rect 16038 20102 16068 20154
rect 16092 20102 16102 20154
rect 16102 20102 16148 20154
rect 15852 20100 15908 20102
rect 15932 20100 15988 20102
rect 16012 20100 16068 20102
rect 16092 20100 16148 20102
rect 15852 19066 15908 19068
rect 15932 19066 15988 19068
rect 16012 19066 16068 19068
rect 16092 19066 16148 19068
rect 15852 19014 15898 19066
rect 15898 19014 15908 19066
rect 15932 19014 15962 19066
rect 15962 19014 15974 19066
rect 15974 19014 15988 19066
rect 16012 19014 16026 19066
rect 16026 19014 16038 19066
rect 16038 19014 16068 19066
rect 16092 19014 16102 19066
rect 16102 19014 16148 19066
rect 15852 19012 15908 19014
rect 15932 19012 15988 19014
rect 16012 19012 16068 19014
rect 16092 19012 16148 19014
rect 15852 17978 15908 17980
rect 15932 17978 15988 17980
rect 16012 17978 16068 17980
rect 16092 17978 16148 17980
rect 15852 17926 15898 17978
rect 15898 17926 15908 17978
rect 15932 17926 15962 17978
rect 15962 17926 15974 17978
rect 15974 17926 15988 17978
rect 16012 17926 16026 17978
rect 16026 17926 16038 17978
rect 16038 17926 16068 17978
rect 16092 17926 16102 17978
rect 16102 17926 16148 17978
rect 15852 17924 15908 17926
rect 15932 17924 15988 17926
rect 16012 17924 16068 17926
rect 16092 17924 16148 17926
rect 15852 16890 15908 16892
rect 15932 16890 15988 16892
rect 16012 16890 16068 16892
rect 16092 16890 16148 16892
rect 15852 16838 15898 16890
rect 15898 16838 15908 16890
rect 15932 16838 15962 16890
rect 15962 16838 15974 16890
rect 15974 16838 15988 16890
rect 16012 16838 16026 16890
rect 16026 16838 16038 16890
rect 16038 16838 16068 16890
rect 16092 16838 16102 16890
rect 16102 16838 16148 16890
rect 15852 16836 15908 16838
rect 15932 16836 15988 16838
rect 16012 16836 16068 16838
rect 16092 16836 16148 16838
rect 16302 26696 16358 26752
rect 17314 47116 17370 47152
rect 17314 47096 17316 47116
rect 17316 47096 17368 47116
rect 17368 47096 17370 47116
rect 17866 47796 17922 47832
rect 17866 47776 17868 47796
rect 17868 47776 17920 47796
rect 17920 47776 17922 47796
rect 18602 44240 18658 44296
rect 19890 60152 19946 60208
rect 19798 57452 19854 57488
rect 19798 57432 19800 57452
rect 19800 57432 19852 57452
rect 19852 57432 19854 57452
rect 19154 47096 19210 47152
rect 20817 63130 20873 63132
rect 20897 63130 20953 63132
rect 20977 63130 21033 63132
rect 21057 63130 21113 63132
rect 20817 63078 20863 63130
rect 20863 63078 20873 63130
rect 20897 63078 20927 63130
rect 20927 63078 20939 63130
rect 20939 63078 20953 63130
rect 20977 63078 20991 63130
rect 20991 63078 21003 63130
rect 21003 63078 21033 63130
rect 21057 63078 21067 63130
rect 21067 63078 21113 63130
rect 20817 63076 20873 63078
rect 20897 63076 20953 63078
rect 20977 63076 21033 63078
rect 21057 63076 21113 63078
rect 20817 62042 20873 62044
rect 20897 62042 20953 62044
rect 20977 62042 21033 62044
rect 21057 62042 21113 62044
rect 20817 61990 20863 62042
rect 20863 61990 20873 62042
rect 20897 61990 20927 62042
rect 20927 61990 20939 62042
rect 20939 61990 20953 62042
rect 20977 61990 20991 62042
rect 20991 61990 21003 62042
rect 21003 61990 21033 62042
rect 21057 61990 21067 62042
rect 21067 61990 21113 62042
rect 20817 61988 20873 61990
rect 20897 61988 20953 61990
rect 20977 61988 21033 61990
rect 21057 61988 21113 61990
rect 20817 60954 20873 60956
rect 20897 60954 20953 60956
rect 20977 60954 21033 60956
rect 21057 60954 21113 60956
rect 20817 60902 20863 60954
rect 20863 60902 20873 60954
rect 20897 60902 20927 60954
rect 20927 60902 20939 60954
rect 20939 60902 20953 60954
rect 20977 60902 20991 60954
rect 20991 60902 21003 60954
rect 21003 60902 21033 60954
rect 21057 60902 21067 60954
rect 21067 60902 21113 60954
rect 20817 60900 20873 60902
rect 20897 60900 20953 60902
rect 20977 60900 21033 60902
rect 21057 60900 21113 60902
rect 20810 60716 20866 60752
rect 20810 60696 20812 60716
rect 20812 60696 20864 60716
rect 20864 60696 20866 60716
rect 20817 59866 20873 59868
rect 20897 59866 20953 59868
rect 20977 59866 21033 59868
rect 21057 59866 21113 59868
rect 20817 59814 20863 59866
rect 20863 59814 20873 59866
rect 20897 59814 20927 59866
rect 20927 59814 20939 59866
rect 20939 59814 20953 59866
rect 20977 59814 20991 59866
rect 20991 59814 21003 59866
rect 21003 59814 21033 59866
rect 21057 59814 21067 59866
rect 21067 59814 21113 59866
rect 20817 59812 20873 59814
rect 20897 59812 20953 59814
rect 20977 59812 21033 59814
rect 21057 59812 21113 59814
rect 20817 58778 20873 58780
rect 20897 58778 20953 58780
rect 20977 58778 21033 58780
rect 21057 58778 21113 58780
rect 20817 58726 20863 58778
rect 20863 58726 20873 58778
rect 20897 58726 20927 58778
rect 20927 58726 20939 58778
rect 20939 58726 20953 58778
rect 20977 58726 20991 58778
rect 20991 58726 21003 58778
rect 21003 58726 21033 58778
rect 21057 58726 21067 58778
rect 21067 58726 21113 58778
rect 20817 58724 20873 58726
rect 20897 58724 20953 58726
rect 20977 58724 21033 58726
rect 21057 58724 21113 58726
rect 20817 57690 20873 57692
rect 20897 57690 20953 57692
rect 20977 57690 21033 57692
rect 21057 57690 21113 57692
rect 20817 57638 20863 57690
rect 20863 57638 20873 57690
rect 20897 57638 20927 57690
rect 20927 57638 20939 57690
rect 20939 57638 20953 57690
rect 20977 57638 20991 57690
rect 20991 57638 21003 57690
rect 21003 57638 21033 57690
rect 21057 57638 21067 57690
rect 21067 57638 21113 57690
rect 20817 57636 20873 57638
rect 20897 57636 20953 57638
rect 20977 57636 21033 57638
rect 21057 57636 21113 57638
rect 18234 37324 18290 37360
rect 18234 37304 18236 37324
rect 18236 37304 18288 37324
rect 18288 37304 18290 37324
rect 15852 15802 15908 15804
rect 15932 15802 15988 15804
rect 16012 15802 16068 15804
rect 16092 15802 16148 15804
rect 15852 15750 15898 15802
rect 15898 15750 15908 15802
rect 15932 15750 15962 15802
rect 15962 15750 15974 15802
rect 15974 15750 15988 15802
rect 16012 15750 16026 15802
rect 16026 15750 16038 15802
rect 16038 15750 16068 15802
rect 16092 15750 16102 15802
rect 16102 15750 16148 15802
rect 15852 15748 15908 15750
rect 15932 15748 15988 15750
rect 16012 15748 16068 15750
rect 16092 15748 16148 15750
rect 18694 37440 18750 37496
rect 15852 14714 15908 14716
rect 15932 14714 15988 14716
rect 16012 14714 16068 14716
rect 16092 14714 16148 14716
rect 15852 14662 15898 14714
rect 15898 14662 15908 14714
rect 15932 14662 15962 14714
rect 15962 14662 15974 14714
rect 15974 14662 15988 14714
rect 16012 14662 16026 14714
rect 16026 14662 16038 14714
rect 16038 14662 16068 14714
rect 16092 14662 16102 14714
rect 16102 14662 16148 14714
rect 15852 14660 15908 14662
rect 15932 14660 15988 14662
rect 16012 14660 16068 14662
rect 16092 14660 16148 14662
rect 15852 13626 15908 13628
rect 15932 13626 15988 13628
rect 16012 13626 16068 13628
rect 16092 13626 16148 13628
rect 15852 13574 15898 13626
rect 15898 13574 15908 13626
rect 15932 13574 15962 13626
rect 15962 13574 15974 13626
rect 15974 13574 15988 13626
rect 16012 13574 16026 13626
rect 16026 13574 16038 13626
rect 16038 13574 16068 13626
rect 16092 13574 16102 13626
rect 16102 13574 16148 13626
rect 15852 13572 15908 13574
rect 15932 13572 15988 13574
rect 16012 13572 16068 13574
rect 16092 13572 16148 13574
rect 15852 12538 15908 12540
rect 15932 12538 15988 12540
rect 16012 12538 16068 12540
rect 16092 12538 16148 12540
rect 15852 12486 15898 12538
rect 15898 12486 15908 12538
rect 15932 12486 15962 12538
rect 15962 12486 15974 12538
rect 15974 12486 15988 12538
rect 16012 12486 16026 12538
rect 16026 12486 16038 12538
rect 16038 12486 16068 12538
rect 16092 12486 16102 12538
rect 16102 12486 16148 12538
rect 15852 12484 15908 12486
rect 15932 12484 15988 12486
rect 16012 12484 16068 12486
rect 16092 12484 16148 12486
rect 15852 11450 15908 11452
rect 15932 11450 15988 11452
rect 16012 11450 16068 11452
rect 16092 11450 16148 11452
rect 15852 11398 15898 11450
rect 15898 11398 15908 11450
rect 15932 11398 15962 11450
rect 15962 11398 15974 11450
rect 15974 11398 15988 11450
rect 16012 11398 16026 11450
rect 16026 11398 16038 11450
rect 16038 11398 16068 11450
rect 16092 11398 16102 11450
rect 16102 11398 16148 11450
rect 15852 11396 15908 11398
rect 15932 11396 15988 11398
rect 16012 11396 16068 11398
rect 16092 11396 16148 11398
rect 15852 10362 15908 10364
rect 15932 10362 15988 10364
rect 16012 10362 16068 10364
rect 16092 10362 16148 10364
rect 15852 10310 15898 10362
rect 15898 10310 15908 10362
rect 15932 10310 15962 10362
rect 15962 10310 15974 10362
rect 15974 10310 15988 10362
rect 16012 10310 16026 10362
rect 16026 10310 16038 10362
rect 16038 10310 16068 10362
rect 16092 10310 16102 10362
rect 16102 10310 16148 10362
rect 15852 10308 15908 10310
rect 15932 10308 15988 10310
rect 16012 10308 16068 10310
rect 16092 10308 16148 10310
rect 15852 9274 15908 9276
rect 15932 9274 15988 9276
rect 16012 9274 16068 9276
rect 16092 9274 16148 9276
rect 15852 9222 15898 9274
rect 15898 9222 15908 9274
rect 15932 9222 15962 9274
rect 15962 9222 15974 9274
rect 15974 9222 15988 9274
rect 16012 9222 16026 9274
rect 16026 9222 16038 9274
rect 16038 9222 16068 9274
rect 16092 9222 16102 9274
rect 16102 9222 16148 9274
rect 15852 9220 15908 9222
rect 15932 9220 15988 9222
rect 16012 9220 16068 9222
rect 16092 9220 16148 9222
rect 15852 8186 15908 8188
rect 15932 8186 15988 8188
rect 16012 8186 16068 8188
rect 16092 8186 16148 8188
rect 15852 8134 15898 8186
rect 15898 8134 15908 8186
rect 15932 8134 15962 8186
rect 15962 8134 15974 8186
rect 15974 8134 15988 8186
rect 16012 8134 16026 8186
rect 16026 8134 16038 8186
rect 16038 8134 16068 8186
rect 16092 8134 16102 8186
rect 16102 8134 16148 8186
rect 15852 8132 15908 8134
rect 15932 8132 15988 8134
rect 16012 8132 16068 8134
rect 16092 8132 16148 8134
rect 10886 7642 10942 7644
rect 10966 7642 11022 7644
rect 11046 7642 11102 7644
rect 11126 7642 11182 7644
rect 10886 7590 10932 7642
rect 10932 7590 10942 7642
rect 10966 7590 10996 7642
rect 10996 7590 11008 7642
rect 11008 7590 11022 7642
rect 11046 7590 11060 7642
rect 11060 7590 11072 7642
rect 11072 7590 11102 7642
rect 11126 7590 11136 7642
rect 11136 7590 11182 7642
rect 10886 7588 10942 7590
rect 10966 7588 11022 7590
rect 11046 7588 11102 7590
rect 11126 7588 11182 7590
rect 5921 7098 5977 7100
rect 6001 7098 6057 7100
rect 6081 7098 6137 7100
rect 6161 7098 6217 7100
rect 5921 7046 5967 7098
rect 5967 7046 5977 7098
rect 6001 7046 6031 7098
rect 6031 7046 6043 7098
rect 6043 7046 6057 7098
rect 6081 7046 6095 7098
rect 6095 7046 6107 7098
rect 6107 7046 6137 7098
rect 6161 7046 6171 7098
rect 6171 7046 6217 7098
rect 5921 7044 5977 7046
rect 6001 7044 6057 7046
rect 6081 7044 6137 7046
rect 6161 7044 6217 7046
rect 15852 7098 15908 7100
rect 15932 7098 15988 7100
rect 16012 7098 16068 7100
rect 16092 7098 16148 7100
rect 15852 7046 15898 7098
rect 15898 7046 15908 7098
rect 15932 7046 15962 7098
rect 15962 7046 15974 7098
rect 15974 7046 15988 7098
rect 16012 7046 16026 7098
rect 16026 7046 16038 7098
rect 16038 7046 16068 7098
rect 16092 7046 16102 7098
rect 16102 7046 16148 7098
rect 15852 7044 15908 7046
rect 15932 7044 15988 7046
rect 16012 7044 16068 7046
rect 16092 7044 16148 7046
rect 16854 16768 16910 16824
rect 18970 37324 19026 37360
rect 18970 37304 18972 37324
rect 18972 37304 19024 37324
rect 19024 37304 19026 37324
rect 19062 29008 19118 29064
rect 20810 57452 20866 57488
rect 20810 57432 20812 57452
rect 20812 57432 20864 57452
rect 20864 57432 20866 57452
rect 20817 56602 20873 56604
rect 20897 56602 20953 56604
rect 20977 56602 21033 56604
rect 21057 56602 21113 56604
rect 20817 56550 20863 56602
rect 20863 56550 20873 56602
rect 20897 56550 20927 56602
rect 20927 56550 20939 56602
rect 20939 56550 20953 56602
rect 20977 56550 20991 56602
rect 20991 56550 21003 56602
rect 21003 56550 21033 56602
rect 21057 56550 21067 56602
rect 21067 56550 21113 56602
rect 20817 56548 20873 56550
rect 20897 56548 20953 56550
rect 20977 56548 21033 56550
rect 21057 56548 21113 56550
rect 22558 66156 22614 66192
rect 22558 66136 22560 66156
rect 22560 66136 22612 66156
rect 22612 66136 22614 66156
rect 22650 66000 22706 66056
rect 22374 60696 22430 60752
rect 20817 55514 20873 55516
rect 20897 55514 20953 55516
rect 20977 55514 21033 55516
rect 21057 55514 21113 55516
rect 20817 55462 20863 55514
rect 20863 55462 20873 55514
rect 20897 55462 20927 55514
rect 20927 55462 20939 55514
rect 20939 55462 20953 55514
rect 20977 55462 20991 55514
rect 20991 55462 21003 55514
rect 21003 55462 21033 55514
rect 21057 55462 21067 55514
rect 21067 55462 21113 55514
rect 20817 55460 20873 55462
rect 20897 55460 20953 55462
rect 20977 55460 21033 55462
rect 21057 55460 21113 55462
rect 20817 54426 20873 54428
rect 20897 54426 20953 54428
rect 20977 54426 21033 54428
rect 21057 54426 21113 54428
rect 20817 54374 20863 54426
rect 20863 54374 20873 54426
rect 20897 54374 20927 54426
rect 20927 54374 20939 54426
rect 20939 54374 20953 54426
rect 20977 54374 20991 54426
rect 20991 54374 21003 54426
rect 21003 54374 21033 54426
rect 21057 54374 21067 54426
rect 21067 54374 21113 54426
rect 20817 54372 20873 54374
rect 20897 54372 20953 54374
rect 20977 54372 21033 54374
rect 21057 54372 21113 54374
rect 20817 53338 20873 53340
rect 20897 53338 20953 53340
rect 20977 53338 21033 53340
rect 21057 53338 21113 53340
rect 20817 53286 20863 53338
rect 20863 53286 20873 53338
rect 20897 53286 20927 53338
rect 20927 53286 20939 53338
rect 20939 53286 20953 53338
rect 20977 53286 20991 53338
rect 20991 53286 21003 53338
rect 21003 53286 21033 53338
rect 21057 53286 21067 53338
rect 21067 53286 21113 53338
rect 20817 53284 20873 53286
rect 20897 53284 20953 53286
rect 20977 53284 21033 53286
rect 21057 53284 21113 53286
rect 20350 48084 20352 48104
rect 20352 48084 20404 48104
rect 20404 48084 20406 48104
rect 20350 48048 20406 48084
rect 19890 40588 19946 40624
rect 19890 40568 19892 40588
rect 19892 40568 19944 40588
rect 19944 40568 19946 40588
rect 19890 37304 19946 37360
rect 19706 34992 19762 35048
rect 19706 34584 19762 34640
rect 20817 52250 20873 52252
rect 20897 52250 20953 52252
rect 20977 52250 21033 52252
rect 21057 52250 21113 52252
rect 20817 52198 20863 52250
rect 20863 52198 20873 52250
rect 20897 52198 20927 52250
rect 20927 52198 20939 52250
rect 20939 52198 20953 52250
rect 20977 52198 20991 52250
rect 20991 52198 21003 52250
rect 21003 52198 21033 52250
rect 21057 52198 21067 52250
rect 21067 52198 21113 52250
rect 20817 52196 20873 52198
rect 20897 52196 20953 52198
rect 20977 52196 21033 52198
rect 21057 52196 21113 52198
rect 20534 50360 20590 50416
rect 20817 51162 20873 51164
rect 20897 51162 20953 51164
rect 20977 51162 21033 51164
rect 21057 51162 21113 51164
rect 20817 51110 20863 51162
rect 20863 51110 20873 51162
rect 20897 51110 20927 51162
rect 20927 51110 20939 51162
rect 20939 51110 20953 51162
rect 20977 51110 20991 51162
rect 20991 51110 21003 51162
rect 21003 51110 21033 51162
rect 21057 51110 21067 51162
rect 21067 51110 21113 51162
rect 20817 51108 20873 51110
rect 20897 51108 20953 51110
rect 20977 51108 21033 51110
rect 21057 51108 21113 51110
rect 21086 50904 21142 50960
rect 20817 50074 20873 50076
rect 20897 50074 20953 50076
rect 20977 50074 21033 50076
rect 21057 50074 21113 50076
rect 20817 50022 20863 50074
rect 20863 50022 20873 50074
rect 20897 50022 20927 50074
rect 20927 50022 20939 50074
rect 20939 50022 20953 50074
rect 20977 50022 20991 50074
rect 20991 50022 21003 50074
rect 21003 50022 21033 50074
rect 21057 50022 21067 50074
rect 21067 50022 21113 50074
rect 20817 50020 20873 50022
rect 20897 50020 20953 50022
rect 20977 50020 21033 50022
rect 21057 50020 21113 50022
rect 20817 48986 20873 48988
rect 20897 48986 20953 48988
rect 20977 48986 21033 48988
rect 21057 48986 21113 48988
rect 20817 48934 20863 48986
rect 20863 48934 20873 48986
rect 20897 48934 20927 48986
rect 20927 48934 20939 48986
rect 20939 48934 20953 48986
rect 20977 48934 20991 48986
rect 20991 48934 21003 48986
rect 21003 48934 21033 48986
rect 21057 48934 21067 48986
rect 21067 48934 21113 48986
rect 20817 48932 20873 48934
rect 20897 48932 20953 48934
rect 20977 48932 21033 48934
rect 21057 48932 21113 48934
rect 20817 47898 20873 47900
rect 20897 47898 20953 47900
rect 20977 47898 21033 47900
rect 21057 47898 21113 47900
rect 20817 47846 20863 47898
rect 20863 47846 20873 47898
rect 20897 47846 20927 47898
rect 20927 47846 20939 47898
rect 20939 47846 20953 47898
rect 20977 47846 20991 47898
rect 20991 47846 21003 47898
rect 21003 47846 21033 47898
rect 21057 47846 21067 47898
rect 21067 47846 21113 47898
rect 20817 47844 20873 47846
rect 20897 47844 20953 47846
rect 20977 47844 21033 47846
rect 21057 47844 21113 47846
rect 20817 46810 20873 46812
rect 20897 46810 20953 46812
rect 20977 46810 21033 46812
rect 21057 46810 21113 46812
rect 20817 46758 20863 46810
rect 20863 46758 20873 46810
rect 20897 46758 20927 46810
rect 20927 46758 20939 46810
rect 20939 46758 20953 46810
rect 20977 46758 20991 46810
rect 20991 46758 21003 46810
rect 21003 46758 21033 46810
rect 21057 46758 21067 46810
rect 21067 46758 21113 46810
rect 20817 46756 20873 46758
rect 20897 46756 20953 46758
rect 20977 46756 21033 46758
rect 21057 46756 21113 46758
rect 20817 45722 20873 45724
rect 20897 45722 20953 45724
rect 20977 45722 21033 45724
rect 21057 45722 21113 45724
rect 20817 45670 20863 45722
rect 20863 45670 20873 45722
rect 20897 45670 20927 45722
rect 20927 45670 20939 45722
rect 20939 45670 20953 45722
rect 20977 45670 20991 45722
rect 20991 45670 21003 45722
rect 21003 45670 21033 45722
rect 21057 45670 21067 45722
rect 21067 45670 21113 45722
rect 20817 45668 20873 45670
rect 20897 45668 20953 45670
rect 20977 45668 21033 45670
rect 21057 45668 21113 45670
rect 20817 44634 20873 44636
rect 20897 44634 20953 44636
rect 20977 44634 21033 44636
rect 21057 44634 21113 44636
rect 20817 44582 20863 44634
rect 20863 44582 20873 44634
rect 20897 44582 20927 44634
rect 20927 44582 20939 44634
rect 20939 44582 20953 44634
rect 20977 44582 20991 44634
rect 20991 44582 21003 44634
rect 21003 44582 21033 44634
rect 21057 44582 21067 44634
rect 21067 44582 21113 44634
rect 20817 44580 20873 44582
rect 20897 44580 20953 44582
rect 20977 44580 21033 44582
rect 21057 44580 21113 44582
rect 20817 43546 20873 43548
rect 20897 43546 20953 43548
rect 20977 43546 21033 43548
rect 21057 43546 21113 43548
rect 20817 43494 20863 43546
rect 20863 43494 20873 43546
rect 20897 43494 20927 43546
rect 20927 43494 20939 43546
rect 20939 43494 20953 43546
rect 20977 43494 20991 43546
rect 20991 43494 21003 43546
rect 21003 43494 21033 43546
rect 21057 43494 21067 43546
rect 21067 43494 21113 43546
rect 20817 43492 20873 43494
rect 20897 43492 20953 43494
rect 20977 43492 21033 43494
rect 21057 43492 21113 43494
rect 21546 51032 21602 51088
rect 21546 50904 21602 50960
rect 21730 48592 21786 48648
rect 20817 42458 20873 42460
rect 20897 42458 20953 42460
rect 20977 42458 21033 42460
rect 21057 42458 21113 42460
rect 20817 42406 20863 42458
rect 20863 42406 20873 42458
rect 20897 42406 20927 42458
rect 20927 42406 20939 42458
rect 20939 42406 20953 42458
rect 20977 42406 20991 42458
rect 20991 42406 21003 42458
rect 21003 42406 21033 42458
rect 21057 42406 21067 42458
rect 21067 42406 21113 42458
rect 20817 42404 20873 42406
rect 20897 42404 20953 42406
rect 20977 42404 21033 42406
rect 21057 42404 21113 42406
rect 20817 41370 20873 41372
rect 20897 41370 20953 41372
rect 20977 41370 21033 41372
rect 21057 41370 21113 41372
rect 20817 41318 20863 41370
rect 20863 41318 20873 41370
rect 20897 41318 20927 41370
rect 20927 41318 20939 41370
rect 20939 41318 20953 41370
rect 20977 41318 20991 41370
rect 20991 41318 21003 41370
rect 21003 41318 21033 41370
rect 21057 41318 21067 41370
rect 21067 41318 21113 41370
rect 20817 41316 20873 41318
rect 20897 41316 20953 41318
rect 20977 41316 21033 41318
rect 21057 41316 21113 41318
rect 20817 40282 20873 40284
rect 20897 40282 20953 40284
rect 20977 40282 21033 40284
rect 21057 40282 21113 40284
rect 20817 40230 20863 40282
rect 20863 40230 20873 40282
rect 20897 40230 20927 40282
rect 20927 40230 20939 40282
rect 20939 40230 20953 40282
rect 20977 40230 20991 40282
rect 20991 40230 21003 40282
rect 21003 40230 21033 40282
rect 21057 40230 21067 40282
rect 21067 40230 21113 40282
rect 20817 40228 20873 40230
rect 20897 40228 20953 40230
rect 20977 40228 21033 40230
rect 21057 40228 21113 40230
rect 21270 40876 21272 40896
rect 21272 40876 21324 40896
rect 21324 40876 21326 40896
rect 21270 40840 21326 40876
rect 20817 39194 20873 39196
rect 20897 39194 20953 39196
rect 20977 39194 21033 39196
rect 21057 39194 21113 39196
rect 20817 39142 20863 39194
rect 20863 39142 20873 39194
rect 20897 39142 20927 39194
rect 20927 39142 20939 39194
rect 20939 39142 20953 39194
rect 20977 39142 20991 39194
rect 20991 39142 21003 39194
rect 21003 39142 21033 39194
rect 21057 39142 21067 39194
rect 21067 39142 21113 39194
rect 20817 39140 20873 39142
rect 20897 39140 20953 39142
rect 20977 39140 21033 39142
rect 21057 39140 21113 39142
rect 20817 38106 20873 38108
rect 20897 38106 20953 38108
rect 20977 38106 21033 38108
rect 21057 38106 21113 38108
rect 20817 38054 20863 38106
rect 20863 38054 20873 38106
rect 20897 38054 20927 38106
rect 20927 38054 20939 38106
rect 20939 38054 20953 38106
rect 20977 38054 20991 38106
rect 20991 38054 21003 38106
rect 21003 38054 21033 38106
rect 21057 38054 21067 38106
rect 21067 38054 21113 38106
rect 20817 38052 20873 38054
rect 20897 38052 20953 38054
rect 20977 38052 21033 38054
rect 21057 38052 21113 38054
rect 20817 37018 20873 37020
rect 20897 37018 20953 37020
rect 20977 37018 21033 37020
rect 21057 37018 21113 37020
rect 20817 36966 20863 37018
rect 20863 36966 20873 37018
rect 20897 36966 20927 37018
rect 20927 36966 20939 37018
rect 20939 36966 20953 37018
rect 20977 36966 20991 37018
rect 20991 36966 21003 37018
rect 21003 36966 21033 37018
rect 21057 36966 21067 37018
rect 21067 36966 21113 37018
rect 20817 36964 20873 36966
rect 20897 36964 20953 36966
rect 20977 36964 21033 36966
rect 21057 36964 21113 36966
rect 19614 29180 19616 29200
rect 19616 29180 19668 29200
rect 19668 29180 19670 29200
rect 19614 29144 19670 29180
rect 20817 35930 20873 35932
rect 20897 35930 20953 35932
rect 20977 35930 21033 35932
rect 21057 35930 21113 35932
rect 20817 35878 20863 35930
rect 20863 35878 20873 35930
rect 20897 35878 20927 35930
rect 20927 35878 20939 35930
rect 20939 35878 20953 35930
rect 20977 35878 20991 35930
rect 20991 35878 21003 35930
rect 21003 35878 21033 35930
rect 21057 35878 21067 35930
rect 21067 35878 21113 35930
rect 20817 35876 20873 35878
rect 20897 35876 20953 35878
rect 20977 35876 21033 35878
rect 21057 35876 21113 35878
rect 20817 34842 20873 34844
rect 20897 34842 20953 34844
rect 20977 34842 21033 34844
rect 21057 34842 21113 34844
rect 20817 34790 20863 34842
rect 20863 34790 20873 34842
rect 20897 34790 20927 34842
rect 20927 34790 20939 34842
rect 20939 34790 20953 34842
rect 20977 34790 20991 34842
rect 20991 34790 21003 34842
rect 21003 34790 21033 34842
rect 21057 34790 21067 34842
rect 21067 34790 21113 34842
rect 20817 34788 20873 34790
rect 20897 34788 20953 34790
rect 20977 34788 21033 34790
rect 21057 34788 21113 34790
rect 20817 33754 20873 33756
rect 20897 33754 20953 33756
rect 20977 33754 21033 33756
rect 21057 33754 21113 33756
rect 20817 33702 20863 33754
rect 20863 33702 20873 33754
rect 20897 33702 20927 33754
rect 20927 33702 20939 33754
rect 20939 33702 20953 33754
rect 20977 33702 20991 33754
rect 20991 33702 21003 33754
rect 21003 33702 21033 33754
rect 21057 33702 21067 33754
rect 21067 33702 21113 33754
rect 20817 33700 20873 33702
rect 20897 33700 20953 33702
rect 20977 33700 21033 33702
rect 21057 33700 21113 33702
rect 22006 50904 22062 50960
rect 21914 49544 21970 49600
rect 22190 46416 22246 46472
rect 22834 55256 22890 55312
rect 23478 57024 23534 57080
rect 23294 56480 23350 56536
rect 23202 55256 23258 55312
rect 23202 55156 23204 55176
rect 23204 55156 23256 55176
rect 23256 55156 23258 55176
rect 23202 55120 23258 55156
rect 22650 50224 22706 50280
rect 22834 49952 22890 50008
rect 22006 43288 22062 43344
rect 22282 42508 22284 42528
rect 22284 42508 22336 42528
rect 22336 42508 22338 42528
rect 22282 42472 22338 42508
rect 22098 41692 22100 41712
rect 22100 41692 22152 41712
rect 22152 41692 22154 41712
rect 22098 41656 22154 41692
rect 21730 38256 21786 38312
rect 22098 40160 22154 40216
rect 22190 38120 22246 38176
rect 21270 32852 21272 32872
rect 21272 32852 21324 32872
rect 21324 32852 21326 32872
rect 21270 32816 21326 32852
rect 20817 32666 20873 32668
rect 20897 32666 20953 32668
rect 20977 32666 21033 32668
rect 21057 32666 21113 32668
rect 20817 32614 20863 32666
rect 20863 32614 20873 32666
rect 20897 32614 20927 32666
rect 20927 32614 20939 32666
rect 20939 32614 20953 32666
rect 20977 32614 20991 32666
rect 20991 32614 21003 32666
rect 21003 32614 21033 32666
rect 21057 32614 21067 32666
rect 21067 32614 21113 32666
rect 20817 32612 20873 32614
rect 20897 32612 20953 32614
rect 20977 32612 21033 32614
rect 21057 32612 21113 32614
rect 20817 31578 20873 31580
rect 20897 31578 20953 31580
rect 20977 31578 21033 31580
rect 21057 31578 21113 31580
rect 20817 31526 20863 31578
rect 20863 31526 20873 31578
rect 20897 31526 20927 31578
rect 20927 31526 20939 31578
rect 20939 31526 20953 31578
rect 20977 31526 20991 31578
rect 20991 31526 21003 31578
rect 21003 31526 21033 31578
rect 21057 31526 21067 31578
rect 21067 31526 21113 31578
rect 20817 31524 20873 31526
rect 20897 31524 20953 31526
rect 20977 31524 21033 31526
rect 21057 31524 21113 31526
rect 20817 30490 20873 30492
rect 20897 30490 20953 30492
rect 20977 30490 21033 30492
rect 21057 30490 21113 30492
rect 20817 30438 20863 30490
rect 20863 30438 20873 30490
rect 20897 30438 20927 30490
rect 20927 30438 20939 30490
rect 20939 30438 20953 30490
rect 20977 30438 20991 30490
rect 20991 30438 21003 30490
rect 21003 30438 21033 30490
rect 21057 30438 21067 30490
rect 21067 30438 21113 30490
rect 20817 30436 20873 30438
rect 20897 30436 20953 30438
rect 20977 30436 21033 30438
rect 21057 30436 21113 30438
rect 20817 29402 20873 29404
rect 20897 29402 20953 29404
rect 20977 29402 21033 29404
rect 21057 29402 21113 29404
rect 20817 29350 20863 29402
rect 20863 29350 20873 29402
rect 20897 29350 20927 29402
rect 20927 29350 20939 29402
rect 20939 29350 20953 29402
rect 20977 29350 20991 29402
rect 20991 29350 21003 29402
rect 21003 29350 21033 29402
rect 21057 29350 21067 29402
rect 21067 29350 21113 29402
rect 20817 29348 20873 29350
rect 20897 29348 20953 29350
rect 20977 29348 21033 29350
rect 21057 29348 21113 29350
rect 18142 15816 18198 15872
rect 18694 16360 18750 16416
rect 19246 16788 19302 16824
rect 19246 16768 19248 16788
rect 19248 16768 19300 16788
rect 19300 16768 19302 16788
rect 18878 16668 18880 16688
rect 18880 16668 18932 16688
rect 18932 16668 18934 16688
rect 18878 16632 18934 16668
rect 18878 16516 18934 16552
rect 18878 16496 18880 16516
rect 18880 16496 18932 16516
rect 18932 16496 18934 16516
rect 19522 16496 19578 16552
rect 19522 14492 19524 14512
rect 19524 14492 19576 14512
rect 19576 14492 19578 14512
rect 19522 14456 19578 14492
rect 19890 16652 19946 16688
rect 19890 16632 19892 16652
rect 19892 16632 19944 16652
rect 19944 16632 19946 16652
rect 19890 16396 19892 16416
rect 19892 16396 19944 16416
rect 19944 16396 19946 16416
rect 19890 16360 19946 16396
rect 19614 11228 19616 11248
rect 19616 11228 19668 11248
rect 19668 11228 19670 11248
rect 19614 11192 19670 11228
rect 20817 28314 20873 28316
rect 20897 28314 20953 28316
rect 20977 28314 21033 28316
rect 21057 28314 21113 28316
rect 20817 28262 20863 28314
rect 20863 28262 20873 28314
rect 20897 28262 20927 28314
rect 20927 28262 20939 28314
rect 20939 28262 20953 28314
rect 20977 28262 20991 28314
rect 20991 28262 21003 28314
rect 21003 28262 21033 28314
rect 21057 28262 21067 28314
rect 21067 28262 21113 28314
rect 20817 28260 20873 28262
rect 20897 28260 20953 28262
rect 20977 28260 21033 28262
rect 21057 28260 21113 28262
rect 20817 27226 20873 27228
rect 20897 27226 20953 27228
rect 20977 27226 21033 27228
rect 21057 27226 21113 27228
rect 20817 27174 20863 27226
rect 20863 27174 20873 27226
rect 20897 27174 20927 27226
rect 20927 27174 20939 27226
rect 20939 27174 20953 27226
rect 20977 27174 20991 27226
rect 20991 27174 21003 27226
rect 21003 27174 21033 27226
rect 21057 27174 21067 27226
rect 21067 27174 21113 27226
rect 20817 27172 20873 27174
rect 20897 27172 20953 27174
rect 20977 27172 21033 27174
rect 21057 27172 21113 27174
rect 20817 26138 20873 26140
rect 20897 26138 20953 26140
rect 20977 26138 21033 26140
rect 21057 26138 21113 26140
rect 20817 26086 20863 26138
rect 20863 26086 20873 26138
rect 20897 26086 20927 26138
rect 20927 26086 20939 26138
rect 20939 26086 20953 26138
rect 20977 26086 20991 26138
rect 20991 26086 21003 26138
rect 21003 26086 21033 26138
rect 21057 26086 21067 26138
rect 21067 26086 21113 26138
rect 20817 26084 20873 26086
rect 20897 26084 20953 26086
rect 20977 26084 21033 26086
rect 21057 26084 21113 26086
rect 20817 25050 20873 25052
rect 20897 25050 20953 25052
rect 20977 25050 21033 25052
rect 21057 25050 21113 25052
rect 20817 24998 20863 25050
rect 20863 24998 20873 25050
rect 20897 24998 20927 25050
rect 20927 24998 20939 25050
rect 20939 24998 20953 25050
rect 20977 24998 20991 25050
rect 20991 24998 21003 25050
rect 21003 24998 21033 25050
rect 21057 24998 21067 25050
rect 21067 24998 21113 25050
rect 20817 24996 20873 24998
rect 20897 24996 20953 24998
rect 20977 24996 21033 24998
rect 21057 24996 21113 24998
rect 20817 23962 20873 23964
rect 20897 23962 20953 23964
rect 20977 23962 21033 23964
rect 21057 23962 21113 23964
rect 20817 23910 20863 23962
rect 20863 23910 20873 23962
rect 20897 23910 20927 23962
rect 20927 23910 20939 23962
rect 20939 23910 20953 23962
rect 20977 23910 20991 23962
rect 20991 23910 21003 23962
rect 21003 23910 21033 23962
rect 21057 23910 21067 23962
rect 21067 23910 21113 23962
rect 20817 23908 20873 23910
rect 20897 23908 20953 23910
rect 20977 23908 21033 23910
rect 21057 23908 21113 23910
rect 20817 22874 20873 22876
rect 20897 22874 20953 22876
rect 20977 22874 21033 22876
rect 21057 22874 21113 22876
rect 20817 22822 20863 22874
rect 20863 22822 20873 22874
rect 20897 22822 20927 22874
rect 20927 22822 20939 22874
rect 20939 22822 20953 22874
rect 20977 22822 20991 22874
rect 20991 22822 21003 22874
rect 21003 22822 21033 22874
rect 21057 22822 21067 22874
rect 21067 22822 21113 22874
rect 20817 22820 20873 22822
rect 20897 22820 20953 22822
rect 20977 22820 21033 22822
rect 21057 22820 21113 22822
rect 20817 21786 20873 21788
rect 20897 21786 20953 21788
rect 20977 21786 21033 21788
rect 21057 21786 21113 21788
rect 20817 21734 20863 21786
rect 20863 21734 20873 21786
rect 20897 21734 20927 21786
rect 20927 21734 20939 21786
rect 20939 21734 20953 21786
rect 20977 21734 20991 21786
rect 20991 21734 21003 21786
rect 21003 21734 21033 21786
rect 21057 21734 21067 21786
rect 21067 21734 21113 21786
rect 20817 21732 20873 21734
rect 20897 21732 20953 21734
rect 20977 21732 21033 21734
rect 21057 21732 21113 21734
rect 20817 20698 20873 20700
rect 20897 20698 20953 20700
rect 20977 20698 21033 20700
rect 21057 20698 21113 20700
rect 20817 20646 20863 20698
rect 20863 20646 20873 20698
rect 20897 20646 20927 20698
rect 20927 20646 20939 20698
rect 20939 20646 20953 20698
rect 20977 20646 20991 20698
rect 20991 20646 21003 20698
rect 21003 20646 21033 20698
rect 21057 20646 21067 20698
rect 21067 20646 21113 20698
rect 20817 20644 20873 20646
rect 20897 20644 20953 20646
rect 20977 20644 21033 20646
rect 21057 20644 21113 20646
rect 20817 19610 20873 19612
rect 20897 19610 20953 19612
rect 20977 19610 21033 19612
rect 21057 19610 21113 19612
rect 20817 19558 20863 19610
rect 20863 19558 20873 19610
rect 20897 19558 20927 19610
rect 20927 19558 20939 19610
rect 20939 19558 20953 19610
rect 20977 19558 20991 19610
rect 20991 19558 21003 19610
rect 21003 19558 21033 19610
rect 21057 19558 21067 19610
rect 21067 19558 21113 19610
rect 20817 19556 20873 19558
rect 20897 19556 20953 19558
rect 20977 19556 21033 19558
rect 21057 19556 21113 19558
rect 20817 18522 20873 18524
rect 20897 18522 20953 18524
rect 20977 18522 21033 18524
rect 21057 18522 21113 18524
rect 20817 18470 20863 18522
rect 20863 18470 20873 18522
rect 20897 18470 20927 18522
rect 20927 18470 20939 18522
rect 20939 18470 20953 18522
rect 20977 18470 20991 18522
rect 20991 18470 21003 18522
rect 21003 18470 21033 18522
rect 21057 18470 21067 18522
rect 21067 18470 21113 18522
rect 20817 18468 20873 18470
rect 20897 18468 20953 18470
rect 20977 18468 21033 18470
rect 21057 18468 21113 18470
rect 20817 17434 20873 17436
rect 20897 17434 20953 17436
rect 20977 17434 21033 17436
rect 21057 17434 21113 17436
rect 20817 17382 20863 17434
rect 20863 17382 20873 17434
rect 20897 17382 20927 17434
rect 20927 17382 20939 17434
rect 20939 17382 20953 17434
rect 20977 17382 20991 17434
rect 20991 17382 21003 17434
rect 21003 17382 21033 17434
rect 21057 17382 21067 17434
rect 21067 17382 21113 17434
rect 20817 17380 20873 17382
rect 20897 17380 20953 17382
rect 20977 17380 21033 17382
rect 21057 17380 21113 17382
rect 23018 49816 23074 49872
rect 22098 29824 22154 29880
rect 21914 24792 21970 24848
rect 20817 16346 20873 16348
rect 20897 16346 20953 16348
rect 20977 16346 21033 16348
rect 21057 16346 21113 16348
rect 20817 16294 20863 16346
rect 20863 16294 20873 16346
rect 20897 16294 20927 16346
rect 20927 16294 20939 16346
rect 20939 16294 20953 16346
rect 20977 16294 20991 16346
rect 20991 16294 21003 16346
rect 21003 16294 21033 16346
rect 21057 16294 21067 16346
rect 21067 16294 21113 16346
rect 20817 16292 20873 16294
rect 20897 16292 20953 16294
rect 20977 16292 21033 16294
rect 21057 16292 21113 16294
rect 21178 15816 21234 15872
rect 20817 15258 20873 15260
rect 20897 15258 20953 15260
rect 20977 15258 21033 15260
rect 21057 15258 21113 15260
rect 20817 15206 20863 15258
rect 20863 15206 20873 15258
rect 20897 15206 20927 15258
rect 20927 15206 20939 15258
rect 20939 15206 20953 15258
rect 20977 15206 20991 15258
rect 20991 15206 21003 15258
rect 21003 15206 21033 15258
rect 21057 15206 21067 15258
rect 21067 15206 21113 15258
rect 20817 15204 20873 15206
rect 20897 15204 20953 15206
rect 20977 15204 21033 15206
rect 21057 15204 21113 15206
rect 20817 14170 20873 14172
rect 20897 14170 20953 14172
rect 20977 14170 21033 14172
rect 21057 14170 21113 14172
rect 20817 14118 20863 14170
rect 20863 14118 20873 14170
rect 20897 14118 20927 14170
rect 20927 14118 20939 14170
rect 20939 14118 20953 14170
rect 20977 14118 20991 14170
rect 20991 14118 21003 14170
rect 21003 14118 21033 14170
rect 21057 14118 21067 14170
rect 21067 14118 21113 14170
rect 20817 14116 20873 14118
rect 20897 14116 20953 14118
rect 20977 14116 21033 14118
rect 21057 14116 21113 14118
rect 20817 13082 20873 13084
rect 20897 13082 20953 13084
rect 20977 13082 21033 13084
rect 21057 13082 21113 13084
rect 20817 13030 20863 13082
rect 20863 13030 20873 13082
rect 20897 13030 20927 13082
rect 20927 13030 20939 13082
rect 20939 13030 20953 13082
rect 20977 13030 20991 13082
rect 20991 13030 21003 13082
rect 21003 13030 21033 13082
rect 21057 13030 21067 13082
rect 21067 13030 21113 13082
rect 20817 13028 20873 13030
rect 20897 13028 20953 13030
rect 20977 13028 21033 13030
rect 21057 13028 21113 13030
rect 20817 11994 20873 11996
rect 20897 11994 20953 11996
rect 20977 11994 21033 11996
rect 21057 11994 21113 11996
rect 20817 11942 20863 11994
rect 20863 11942 20873 11994
rect 20897 11942 20927 11994
rect 20927 11942 20939 11994
rect 20939 11942 20953 11994
rect 20977 11942 20991 11994
rect 20991 11942 21003 11994
rect 21003 11942 21033 11994
rect 21057 11942 21067 11994
rect 21067 11942 21113 11994
rect 20817 11940 20873 11942
rect 20897 11940 20953 11942
rect 20977 11940 21033 11942
rect 21057 11940 21113 11942
rect 21362 11192 21418 11248
rect 20817 10906 20873 10908
rect 20897 10906 20953 10908
rect 20977 10906 21033 10908
rect 21057 10906 21113 10908
rect 20817 10854 20863 10906
rect 20863 10854 20873 10906
rect 20897 10854 20927 10906
rect 20927 10854 20939 10906
rect 20939 10854 20953 10906
rect 20977 10854 20991 10906
rect 20991 10854 21003 10906
rect 21003 10854 21033 10906
rect 21057 10854 21067 10906
rect 21067 10854 21113 10906
rect 20817 10852 20873 10854
rect 20897 10852 20953 10854
rect 20977 10852 21033 10854
rect 21057 10852 21113 10854
rect 23018 41656 23074 41712
rect 23570 56616 23626 56672
rect 23662 52944 23718 53000
rect 23662 52844 23664 52864
rect 23664 52844 23716 52864
rect 23716 52844 23718 52864
rect 23662 52808 23718 52844
rect 23846 55800 23902 55856
rect 23846 55120 23902 55176
rect 23846 53624 23902 53680
rect 23478 51312 23534 51368
rect 23386 49816 23442 49872
rect 23294 43152 23350 43208
rect 23294 42356 23350 42392
rect 23294 42336 23296 42356
rect 23296 42336 23348 42356
rect 23348 42336 23350 42356
rect 22926 37848 22982 37904
rect 22926 36896 22982 36952
rect 22926 32852 22928 32872
rect 22928 32852 22980 32872
rect 22980 32852 22982 32872
rect 22926 32816 22982 32852
rect 24122 59064 24178 59120
rect 24122 57296 24178 57352
rect 24030 53352 24086 53408
rect 23938 52264 23994 52320
rect 23846 51448 23902 51504
rect 23754 50904 23810 50960
rect 23754 50380 23810 50416
rect 23754 50360 23756 50380
rect 23756 50360 23808 50380
rect 23808 50360 23810 50380
rect 23662 49952 23718 50008
rect 23754 43732 23756 43752
rect 23756 43732 23808 43752
rect 23808 43732 23810 43752
rect 23754 43696 23810 43732
rect 23478 41520 23534 41576
rect 23294 40876 23296 40896
rect 23296 40876 23348 40896
rect 23348 40876 23350 40896
rect 23294 40840 23350 40876
rect 23386 38412 23442 38448
rect 23386 38392 23388 38412
rect 23388 38392 23440 38412
rect 23440 38392 23442 38412
rect 23202 32136 23258 32192
rect 22926 31456 22982 31512
rect 22374 23160 22430 23216
rect 22926 24812 22982 24848
rect 22926 24792 22928 24812
rect 22928 24792 22980 24812
rect 22980 24792 22982 24812
rect 22650 22616 22706 22672
rect 23386 31712 23442 31768
rect 23294 31456 23350 31512
rect 23938 49952 23994 50008
rect 24030 43188 24032 43208
rect 24032 43188 24084 43208
rect 24084 43188 24086 43208
rect 24030 43152 24086 43188
rect 24030 43016 24086 43072
rect 24030 42200 24086 42256
rect 24030 40704 24086 40760
rect 23846 38936 23902 38992
rect 24214 55392 24270 55448
rect 24214 54848 24270 54904
rect 25782 74554 25838 74556
rect 25862 74554 25918 74556
rect 25942 74554 25998 74556
rect 26022 74554 26078 74556
rect 25782 74502 25828 74554
rect 25828 74502 25838 74554
rect 25862 74502 25892 74554
rect 25892 74502 25904 74554
rect 25904 74502 25918 74554
rect 25942 74502 25956 74554
rect 25956 74502 25968 74554
rect 25968 74502 25998 74554
rect 26022 74502 26032 74554
rect 26032 74502 26078 74554
rect 25782 74500 25838 74502
rect 25862 74500 25918 74502
rect 25942 74500 25998 74502
rect 26022 74500 26078 74502
rect 25782 73466 25838 73468
rect 25862 73466 25918 73468
rect 25942 73466 25998 73468
rect 26022 73466 26078 73468
rect 25782 73414 25828 73466
rect 25828 73414 25838 73466
rect 25862 73414 25892 73466
rect 25892 73414 25904 73466
rect 25904 73414 25918 73466
rect 25942 73414 25956 73466
rect 25956 73414 25968 73466
rect 25968 73414 25998 73466
rect 26022 73414 26032 73466
rect 26032 73414 26078 73466
rect 25782 73412 25838 73414
rect 25862 73412 25918 73414
rect 25942 73412 25998 73414
rect 26022 73412 26078 73414
rect 25782 72378 25838 72380
rect 25862 72378 25918 72380
rect 25942 72378 25998 72380
rect 26022 72378 26078 72380
rect 25782 72326 25828 72378
rect 25828 72326 25838 72378
rect 25862 72326 25892 72378
rect 25892 72326 25904 72378
rect 25904 72326 25918 72378
rect 25942 72326 25956 72378
rect 25956 72326 25968 72378
rect 25968 72326 25998 72378
rect 26022 72326 26032 72378
rect 26032 72326 26078 72378
rect 25782 72324 25838 72326
rect 25862 72324 25918 72326
rect 25942 72324 25998 72326
rect 26022 72324 26078 72326
rect 25782 71290 25838 71292
rect 25862 71290 25918 71292
rect 25942 71290 25998 71292
rect 26022 71290 26078 71292
rect 25782 71238 25828 71290
rect 25828 71238 25838 71290
rect 25862 71238 25892 71290
rect 25892 71238 25904 71290
rect 25904 71238 25918 71290
rect 25942 71238 25956 71290
rect 25956 71238 25968 71290
rect 25968 71238 25998 71290
rect 26022 71238 26032 71290
rect 26032 71238 26078 71290
rect 25782 71236 25838 71238
rect 25862 71236 25918 71238
rect 25942 71236 25998 71238
rect 26022 71236 26078 71238
rect 25782 70202 25838 70204
rect 25862 70202 25918 70204
rect 25942 70202 25998 70204
rect 26022 70202 26078 70204
rect 25782 70150 25828 70202
rect 25828 70150 25838 70202
rect 25862 70150 25892 70202
rect 25892 70150 25904 70202
rect 25904 70150 25918 70202
rect 25942 70150 25956 70202
rect 25956 70150 25968 70202
rect 25968 70150 25998 70202
rect 26022 70150 26032 70202
rect 26032 70150 26078 70202
rect 25782 70148 25838 70150
rect 25862 70148 25918 70150
rect 25942 70148 25998 70150
rect 26022 70148 26078 70150
rect 25042 68176 25098 68232
rect 24858 62328 24914 62384
rect 24766 62056 24822 62112
rect 24858 61648 24914 61704
rect 25042 61648 25098 61704
rect 24582 60424 24638 60480
rect 24582 60288 24638 60344
rect 24674 60016 24730 60072
rect 24582 56888 24638 56944
rect 24398 56772 24454 56808
rect 24398 56752 24400 56772
rect 24400 56752 24452 56772
rect 24452 56752 24454 56772
rect 24582 54984 24638 55040
rect 24306 43696 24362 43752
rect 24306 41248 24362 41304
rect 24214 41112 24270 41168
rect 23570 37984 23626 38040
rect 20817 9818 20873 9820
rect 20897 9818 20953 9820
rect 20977 9818 21033 9820
rect 21057 9818 21113 9820
rect 20817 9766 20863 9818
rect 20863 9766 20873 9818
rect 20897 9766 20927 9818
rect 20927 9766 20939 9818
rect 20939 9766 20953 9818
rect 20977 9766 20991 9818
rect 20991 9766 21003 9818
rect 21003 9766 21033 9818
rect 21057 9766 21067 9818
rect 21067 9766 21113 9818
rect 20817 9764 20873 9766
rect 20897 9764 20953 9766
rect 20977 9764 21033 9766
rect 21057 9764 21113 9766
rect 20817 8730 20873 8732
rect 20897 8730 20953 8732
rect 20977 8730 21033 8732
rect 21057 8730 21113 8732
rect 20817 8678 20863 8730
rect 20863 8678 20873 8730
rect 20897 8678 20927 8730
rect 20927 8678 20939 8730
rect 20939 8678 20953 8730
rect 20977 8678 20991 8730
rect 20991 8678 21003 8730
rect 21003 8678 21033 8730
rect 21057 8678 21067 8730
rect 21067 8678 21113 8730
rect 20817 8676 20873 8678
rect 20897 8676 20953 8678
rect 20977 8676 21033 8678
rect 21057 8676 21113 8678
rect 20817 7642 20873 7644
rect 20897 7642 20953 7644
rect 20977 7642 21033 7644
rect 21057 7642 21113 7644
rect 20817 7590 20863 7642
rect 20863 7590 20873 7642
rect 20897 7590 20927 7642
rect 20927 7590 20939 7642
rect 20939 7590 20953 7642
rect 20977 7590 20991 7642
rect 20991 7590 21003 7642
rect 21003 7590 21033 7642
rect 21057 7590 21067 7642
rect 21067 7590 21113 7642
rect 20817 7588 20873 7590
rect 20897 7588 20953 7590
rect 20977 7588 21033 7590
rect 21057 7588 21113 7590
rect 10886 6554 10942 6556
rect 10966 6554 11022 6556
rect 11046 6554 11102 6556
rect 11126 6554 11182 6556
rect 10886 6502 10932 6554
rect 10932 6502 10942 6554
rect 10966 6502 10996 6554
rect 10996 6502 11008 6554
rect 11008 6502 11022 6554
rect 11046 6502 11060 6554
rect 11060 6502 11072 6554
rect 11072 6502 11102 6554
rect 11126 6502 11136 6554
rect 11136 6502 11182 6554
rect 10886 6500 10942 6502
rect 10966 6500 11022 6502
rect 11046 6500 11102 6502
rect 11126 6500 11182 6502
rect 1582 6180 1638 6216
rect 1582 6160 1584 6180
rect 1584 6160 1636 6180
rect 1636 6160 1638 6180
rect 5921 6010 5977 6012
rect 6001 6010 6057 6012
rect 6081 6010 6137 6012
rect 6161 6010 6217 6012
rect 5921 5958 5967 6010
rect 5967 5958 5977 6010
rect 6001 5958 6031 6010
rect 6031 5958 6043 6010
rect 6043 5958 6057 6010
rect 6081 5958 6095 6010
rect 6095 5958 6107 6010
rect 6107 5958 6137 6010
rect 6161 5958 6171 6010
rect 6171 5958 6217 6010
rect 5921 5956 5977 5958
rect 6001 5956 6057 5958
rect 6081 5956 6137 5958
rect 6161 5956 6217 5958
rect 15852 6010 15908 6012
rect 15932 6010 15988 6012
rect 16012 6010 16068 6012
rect 16092 6010 16148 6012
rect 15852 5958 15898 6010
rect 15898 5958 15908 6010
rect 15932 5958 15962 6010
rect 15962 5958 15974 6010
rect 15974 5958 15988 6010
rect 16012 5958 16026 6010
rect 16026 5958 16038 6010
rect 16038 5958 16068 6010
rect 16092 5958 16102 6010
rect 16102 5958 16148 6010
rect 15852 5956 15908 5958
rect 15932 5956 15988 5958
rect 16012 5956 16068 5958
rect 16092 5956 16148 5958
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 1582 5480 1638 5516
rect 10886 5466 10942 5468
rect 10966 5466 11022 5468
rect 11046 5466 11102 5468
rect 11126 5466 11182 5468
rect 10886 5414 10932 5466
rect 10932 5414 10942 5466
rect 10966 5414 10996 5466
rect 10996 5414 11008 5466
rect 11008 5414 11022 5466
rect 11046 5414 11060 5466
rect 11060 5414 11072 5466
rect 11072 5414 11102 5466
rect 11126 5414 11136 5466
rect 11136 5414 11182 5466
rect 10886 5412 10942 5414
rect 10966 5412 11022 5414
rect 11046 5412 11102 5414
rect 11126 5412 11182 5414
rect 1582 4972 1584 4992
rect 1584 4972 1636 4992
rect 1636 4972 1638 4992
rect 1582 4936 1638 4972
rect 5921 4922 5977 4924
rect 6001 4922 6057 4924
rect 6081 4922 6137 4924
rect 6161 4922 6217 4924
rect 5921 4870 5967 4922
rect 5967 4870 5977 4922
rect 6001 4870 6031 4922
rect 6031 4870 6043 4922
rect 6043 4870 6057 4922
rect 6081 4870 6095 4922
rect 6095 4870 6107 4922
rect 6107 4870 6137 4922
rect 6161 4870 6171 4922
rect 6171 4870 6217 4922
rect 5921 4868 5977 4870
rect 6001 4868 6057 4870
rect 6081 4868 6137 4870
rect 6161 4868 6217 4870
rect 15852 4922 15908 4924
rect 15932 4922 15988 4924
rect 16012 4922 16068 4924
rect 16092 4922 16148 4924
rect 15852 4870 15898 4922
rect 15898 4870 15908 4922
rect 15932 4870 15962 4922
rect 15962 4870 15974 4922
rect 15974 4870 15988 4922
rect 16012 4870 16026 4922
rect 16026 4870 16038 4922
rect 16038 4870 16068 4922
rect 16092 4870 16102 4922
rect 16102 4870 16148 4922
rect 15852 4868 15908 4870
rect 15932 4868 15988 4870
rect 16012 4868 16068 4870
rect 16092 4868 16148 4870
rect 10886 4378 10942 4380
rect 10966 4378 11022 4380
rect 11046 4378 11102 4380
rect 11126 4378 11182 4380
rect 10886 4326 10932 4378
rect 10932 4326 10942 4378
rect 10966 4326 10996 4378
rect 10996 4326 11008 4378
rect 11008 4326 11022 4378
rect 11046 4326 11060 4378
rect 11060 4326 11072 4378
rect 11072 4326 11102 4378
rect 11126 4326 11136 4378
rect 11136 4326 11182 4378
rect 10886 4324 10942 4326
rect 10966 4324 11022 4326
rect 11046 4324 11102 4326
rect 11126 4324 11182 4326
rect 1582 4256 1638 4312
rect 5921 3834 5977 3836
rect 6001 3834 6057 3836
rect 6081 3834 6137 3836
rect 6161 3834 6217 3836
rect 5921 3782 5967 3834
rect 5967 3782 5977 3834
rect 6001 3782 6031 3834
rect 6031 3782 6043 3834
rect 6043 3782 6057 3834
rect 6081 3782 6095 3834
rect 6095 3782 6107 3834
rect 6107 3782 6137 3834
rect 6161 3782 6171 3834
rect 6171 3782 6217 3834
rect 5921 3780 5977 3782
rect 6001 3780 6057 3782
rect 6081 3780 6137 3782
rect 6161 3780 6217 3782
rect 15852 3834 15908 3836
rect 15932 3834 15988 3836
rect 16012 3834 16068 3836
rect 16092 3834 16148 3836
rect 15852 3782 15898 3834
rect 15898 3782 15908 3834
rect 15932 3782 15962 3834
rect 15962 3782 15974 3834
rect 15974 3782 15988 3834
rect 16012 3782 16026 3834
rect 16026 3782 16038 3834
rect 16038 3782 16068 3834
rect 16092 3782 16102 3834
rect 16102 3782 16148 3834
rect 15852 3780 15908 3782
rect 15932 3780 15988 3782
rect 16012 3780 16068 3782
rect 16092 3780 16148 3782
rect 1582 3576 1638 3632
rect 1582 2896 1638 2952
rect 10886 3290 10942 3292
rect 10966 3290 11022 3292
rect 11046 3290 11102 3292
rect 11126 3290 11182 3292
rect 10886 3238 10932 3290
rect 10932 3238 10942 3290
rect 10966 3238 10996 3290
rect 10996 3238 11008 3290
rect 11008 3238 11022 3290
rect 11046 3238 11060 3290
rect 11060 3238 11072 3290
rect 11072 3238 11102 3290
rect 11126 3238 11136 3290
rect 11136 3238 11182 3290
rect 10886 3236 10942 3238
rect 10966 3236 11022 3238
rect 11046 3236 11102 3238
rect 11126 3236 11182 3238
rect 5921 2746 5977 2748
rect 6001 2746 6057 2748
rect 6081 2746 6137 2748
rect 6161 2746 6217 2748
rect 5921 2694 5967 2746
rect 5967 2694 5977 2746
rect 6001 2694 6031 2746
rect 6031 2694 6043 2746
rect 6043 2694 6057 2746
rect 6081 2694 6095 2746
rect 6095 2694 6107 2746
rect 6107 2694 6137 2746
rect 6161 2694 6171 2746
rect 6171 2694 6217 2746
rect 5921 2692 5977 2694
rect 6001 2692 6057 2694
rect 6081 2692 6137 2694
rect 6161 2692 6217 2694
rect 15852 2746 15908 2748
rect 15932 2746 15988 2748
rect 16012 2746 16068 2748
rect 16092 2746 16148 2748
rect 15852 2694 15898 2746
rect 15898 2694 15908 2746
rect 15932 2694 15962 2746
rect 15962 2694 15974 2746
rect 15974 2694 15988 2746
rect 16012 2694 16026 2746
rect 16026 2694 16038 2746
rect 16038 2694 16068 2746
rect 16092 2694 16102 2746
rect 16102 2694 16148 2746
rect 15852 2692 15908 2694
rect 15932 2692 15988 2694
rect 16012 2692 16068 2694
rect 16092 2692 16148 2694
rect 20817 6554 20873 6556
rect 20897 6554 20953 6556
rect 20977 6554 21033 6556
rect 21057 6554 21113 6556
rect 20817 6502 20863 6554
rect 20863 6502 20873 6554
rect 20897 6502 20927 6554
rect 20927 6502 20939 6554
rect 20939 6502 20953 6554
rect 20977 6502 20991 6554
rect 20991 6502 21003 6554
rect 21003 6502 21033 6554
rect 21057 6502 21067 6554
rect 21067 6502 21113 6554
rect 20817 6500 20873 6502
rect 20897 6500 20953 6502
rect 20977 6500 21033 6502
rect 21057 6500 21113 6502
rect 20817 5466 20873 5468
rect 20897 5466 20953 5468
rect 20977 5466 21033 5468
rect 21057 5466 21113 5468
rect 20817 5414 20863 5466
rect 20863 5414 20873 5466
rect 20897 5414 20927 5466
rect 20927 5414 20939 5466
rect 20939 5414 20953 5466
rect 20977 5414 20991 5466
rect 20991 5414 21003 5466
rect 21003 5414 21033 5466
rect 21057 5414 21067 5466
rect 21067 5414 21113 5466
rect 20817 5412 20873 5414
rect 20897 5412 20953 5414
rect 20977 5412 21033 5414
rect 21057 5412 21113 5414
rect 20817 4378 20873 4380
rect 20897 4378 20953 4380
rect 20977 4378 21033 4380
rect 21057 4378 21113 4380
rect 20817 4326 20863 4378
rect 20863 4326 20873 4378
rect 20897 4326 20927 4378
rect 20927 4326 20939 4378
rect 20939 4326 20953 4378
rect 20977 4326 20991 4378
rect 20991 4326 21003 4378
rect 21003 4326 21033 4378
rect 21057 4326 21067 4378
rect 21067 4326 21113 4378
rect 20817 4324 20873 4326
rect 20897 4324 20953 4326
rect 20977 4324 21033 4326
rect 21057 4324 21113 4326
rect 20817 3290 20873 3292
rect 20897 3290 20953 3292
rect 20977 3290 21033 3292
rect 21057 3290 21113 3292
rect 20817 3238 20863 3290
rect 20863 3238 20873 3290
rect 20897 3238 20927 3290
rect 20927 3238 20939 3290
rect 20939 3238 20953 3290
rect 20977 3238 20991 3290
rect 20991 3238 21003 3290
rect 21003 3238 21033 3290
rect 21057 3238 21067 3290
rect 21067 3238 21113 3290
rect 20817 3236 20873 3238
rect 20897 3236 20953 3238
rect 20977 3236 21033 3238
rect 21057 3236 21113 3238
rect 2318 2252 2320 2272
rect 2320 2252 2372 2272
rect 2372 2252 2374 2272
rect 1398 1536 1454 1592
rect 2318 2216 2374 2252
rect 1582 856 1638 912
rect 10886 2202 10942 2204
rect 10966 2202 11022 2204
rect 11046 2202 11102 2204
rect 11126 2202 11182 2204
rect 10886 2150 10932 2202
rect 10932 2150 10942 2202
rect 10966 2150 10996 2202
rect 10996 2150 11008 2202
rect 11008 2150 11022 2202
rect 11046 2150 11060 2202
rect 11060 2150 11072 2202
rect 11072 2150 11102 2202
rect 11126 2150 11136 2202
rect 11136 2150 11182 2202
rect 10886 2148 10942 2150
rect 10966 2148 11022 2150
rect 11046 2148 11102 2150
rect 11126 2148 11182 2150
rect 20817 2202 20873 2204
rect 20897 2202 20953 2204
rect 20977 2202 21033 2204
rect 21057 2202 21113 2204
rect 20817 2150 20863 2202
rect 20863 2150 20873 2202
rect 20897 2150 20927 2202
rect 20927 2150 20939 2202
rect 20939 2150 20953 2202
rect 20977 2150 20991 2202
rect 20991 2150 21003 2202
rect 21003 2150 21033 2202
rect 21057 2150 21067 2202
rect 21067 2150 21113 2202
rect 20817 2148 20873 2150
rect 20897 2148 20953 2150
rect 20977 2148 21033 2150
rect 21057 2148 21113 2150
rect 24030 37712 24086 37768
rect 24122 35284 24178 35320
rect 24122 35264 24124 35284
rect 24124 35264 24176 35284
rect 24176 35264 24178 35284
rect 24214 33768 24270 33824
rect 24582 51348 24584 51368
rect 24584 51348 24636 51368
rect 24636 51348 24638 51368
rect 24582 51312 24638 51348
rect 24490 51040 24546 51096
rect 25042 60424 25098 60480
rect 25226 62328 25282 62384
rect 25782 69114 25838 69116
rect 25862 69114 25918 69116
rect 25942 69114 25998 69116
rect 26022 69114 26078 69116
rect 25782 69062 25828 69114
rect 25828 69062 25838 69114
rect 25862 69062 25892 69114
rect 25892 69062 25904 69114
rect 25904 69062 25918 69114
rect 25942 69062 25956 69114
rect 25956 69062 25968 69114
rect 25968 69062 25998 69114
rect 26022 69062 26032 69114
rect 26032 69062 26078 69114
rect 25782 69060 25838 69062
rect 25862 69060 25918 69062
rect 25942 69060 25998 69062
rect 26022 69060 26078 69062
rect 25782 68026 25838 68028
rect 25862 68026 25918 68028
rect 25942 68026 25998 68028
rect 26022 68026 26078 68028
rect 25782 67974 25828 68026
rect 25828 67974 25838 68026
rect 25862 67974 25892 68026
rect 25892 67974 25904 68026
rect 25904 67974 25918 68026
rect 25942 67974 25956 68026
rect 25956 67974 25968 68026
rect 25968 67974 25998 68026
rect 26022 67974 26032 68026
rect 26032 67974 26078 68026
rect 25782 67972 25838 67974
rect 25862 67972 25918 67974
rect 25942 67972 25998 67974
rect 26022 67972 26078 67974
rect 26054 67804 26056 67824
rect 26056 67804 26108 67824
rect 26108 67804 26110 67824
rect 26054 67768 26110 67804
rect 25686 67632 25742 67688
rect 25410 66000 25466 66056
rect 25318 60832 25374 60888
rect 25226 56652 25228 56672
rect 25228 56652 25280 56672
rect 25280 56652 25282 56672
rect 25226 56616 25282 56652
rect 25134 55800 25190 55856
rect 25782 66938 25838 66940
rect 25862 66938 25918 66940
rect 25942 66938 25998 66940
rect 26022 66938 26078 66940
rect 25782 66886 25828 66938
rect 25828 66886 25838 66938
rect 25862 66886 25892 66938
rect 25892 66886 25904 66938
rect 25904 66886 25918 66938
rect 25942 66886 25956 66938
rect 25956 66886 25968 66938
rect 25968 66886 25998 66938
rect 26022 66886 26032 66938
rect 26032 66886 26078 66938
rect 25782 66884 25838 66886
rect 25862 66884 25918 66886
rect 25942 66884 25998 66886
rect 26022 66884 26078 66886
rect 26238 67088 26294 67144
rect 25782 65850 25838 65852
rect 25862 65850 25918 65852
rect 25942 65850 25998 65852
rect 26022 65850 26078 65852
rect 25782 65798 25828 65850
rect 25828 65798 25838 65850
rect 25862 65798 25892 65850
rect 25892 65798 25904 65850
rect 25904 65798 25918 65850
rect 25942 65798 25956 65850
rect 25956 65798 25968 65850
rect 25968 65798 25998 65850
rect 26022 65798 26032 65850
rect 26032 65798 26078 65850
rect 25782 65796 25838 65798
rect 25862 65796 25918 65798
rect 25942 65796 25998 65798
rect 26022 65796 26078 65798
rect 25782 64762 25838 64764
rect 25862 64762 25918 64764
rect 25942 64762 25998 64764
rect 26022 64762 26078 64764
rect 25782 64710 25828 64762
rect 25828 64710 25838 64762
rect 25862 64710 25892 64762
rect 25892 64710 25904 64762
rect 25904 64710 25918 64762
rect 25942 64710 25956 64762
rect 25956 64710 25968 64762
rect 25968 64710 25998 64762
rect 26022 64710 26032 64762
rect 26032 64710 26078 64762
rect 25782 64708 25838 64710
rect 25862 64708 25918 64710
rect 25942 64708 25998 64710
rect 26022 64708 26078 64710
rect 25782 63674 25838 63676
rect 25862 63674 25918 63676
rect 25942 63674 25998 63676
rect 26022 63674 26078 63676
rect 25782 63622 25828 63674
rect 25828 63622 25838 63674
rect 25862 63622 25892 63674
rect 25892 63622 25904 63674
rect 25904 63622 25918 63674
rect 25942 63622 25956 63674
rect 25956 63622 25968 63674
rect 25968 63622 25998 63674
rect 26022 63622 26032 63674
rect 26032 63622 26078 63674
rect 25782 63620 25838 63622
rect 25862 63620 25918 63622
rect 25942 63620 25998 63622
rect 26022 63620 26078 63622
rect 25782 62586 25838 62588
rect 25862 62586 25918 62588
rect 25942 62586 25998 62588
rect 26022 62586 26078 62588
rect 25782 62534 25828 62586
rect 25828 62534 25838 62586
rect 25862 62534 25892 62586
rect 25892 62534 25904 62586
rect 25904 62534 25918 62586
rect 25942 62534 25956 62586
rect 25956 62534 25968 62586
rect 25968 62534 25998 62586
rect 26022 62534 26032 62586
rect 26032 62534 26078 62586
rect 25782 62532 25838 62534
rect 25862 62532 25918 62534
rect 25942 62532 25998 62534
rect 26022 62532 26078 62534
rect 25782 61498 25838 61500
rect 25862 61498 25918 61500
rect 25942 61498 25998 61500
rect 26022 61498 26078 61500
rect 25782 61446 25828 61498
rect 25828 61446 25838 61498
rect 25862 61446 25892 61498
rect 25892 61446 25904 61498
rect 25904 61446 25918 61498
rect 25942 61446 25956 61498
rect 25956 61446 25968 61498
rect 25968 61446 25998 61498
rect 26022 61446 26032 61498
rect 26032 61446 26078 61498
rect 25782 61444 25838 61446
rect 25862 61444 25918 61446
rect 25942 61444 25998 61446
rect 26022 61444 26078 61446
rect 25778 61124 25834 61160
rect 25778 61104 25780 61124
rect 25780 61104 25832 61124
rect 25832 61104 25834 61124
rect 25594 60832 25650 60888
rect 25042 55392 25098 55448
rect 24950 55120 25006 55176
rect 25042 54848 25098 54904
rect 24950 51584 25006 51640
rect 24858 50904 24914 50960
rect 24858 50632 24914 50688
rect 24858 50496 24914 50552
rect 24490 48728 24546 48784
rect 24582 48456 24638 48512
rect 24490 43968 24546 44024
rect 24766 49972 24822 50008
rect 24766 49952 24768 49972
rect 24768 49952 24820 49972
rect 24820 49952 24822 49972
rect 24674 45056 24730 45112
rect 24490 43016 24546 43072
rect 24766 43152 24822 43208
rect 24766 42880 24822 42936
rect 24674 42608 24730 42664
rect 24950 49680 25006 49736
rect 25502 55800 25558 55856
rect 25226 54032 25282 54088
rect 25134 51040 25190 51096
rect 24858 42608 24914 42664
rect 24766 41248 24822 41304
rect 24582 38800 24638 38856
rect 24674 38612 24730 38668
rect 24582 38392 24638 38448
rect 24674 38256 24730 38312
rect 24306 24656 24362 24712
rect 25226 46144 25282 46200
rect 24858 38612 24914 38668
rect 24858 38120 24914 38176
rect 24858 37884 24878 37904
rect 24878 37884 24914 37904
rect 24858 37848 24914 37884
rect 24858 37576 24914 37632
rect 24766 36116 24768 36136
rect 24768 36116 24820 36136
rect 24820 36116 24822 36136
rect 24766 36080 24822 36116
rect 25134 43016 25190 43072
rect 25870 60696 25926 60752
rect 26330 64404 26332 64424
rect 26332 64404 26384 64424
rect 26384 64404 26386 64424
rect 26330 64368 26386 64404
rect 26514 63008 26570 63064
rect 26238 61104 26294 61160
rect 25962 60560 26018 60616
rect 25782 60410 25838 60412
rect 25862 60410 25918 60412
rect 25942 60410 25998 60412
rect 26022 60410 26078 60412
rect 25782 60358 25828 60410
rect 25828 60358 25838 60410
rect 25862 60358 25892 60410
rect 25892 60358 25904 60410
rect 25904 60358 25918 60410
rect 25942 60358 25956 60410
rect 25956 60358 25968 60410
rect 25968 60358 25998 60410
rect 26022 60358 26032 60410
rect 26032 60358 26078 60410
rect 25782 60356 25838 60358
rect 25862 60356 25918 60358
rect 25942 60356 25998 60358
rect 26022 60356 26078 60358
rect 25778 60152 25834 60208
rect 25870 59880 25926 59936
rect 26146 60152 26202 60208
rect 25870 59608 25926 59664
rect 26054 59608 26110 59664
rect 25782 59322 25838 59324
rect 25862 59322 25918 59324
rect 25942 59322 25998 59324
rect 26022 59322 26078 59324
rect 25782 59270 25828 59322
rect 25828 59270 25838 59322
rect 25862 59270 25892 59322
rect 25892 59270 25904 59322
rect 25904 59270 25918 59322
rect 25942 59270 25956 59322
rect 25956 59270 25968 59322
rect 25968 59270 25998 59322
rect 26022 59270 26032 59322
rect 26032 59270 26078 59322
rect 25782 59268 25838 59270
rect 25862 59268 25918 59270
rect 25942 59268 25998 59270
rect 26022 59268 26078 59270
rect 25782 58234 25838 58236
rect 25862 58234 25918 58236
rect 25942 58234 25998 58236
rect 26022 58234 26078 58236
rect 25782 58182 25828 58234
rect 25828 58182 25838 58234
rect 25862 58182 25892 58234
rect 25892 58182 25904 58234
rect 25904 58182 25918 58234
rect 25942 58182 25956 58234
rect 25956 58182 25968 58234
rect 25968 58182 25998 58234
rect 26022 58182 26032 58234
rect 26032 58182 26078 58234
rect 25782 58180 25838 58182
rect 25862 58180 25918 58182
rect 25942 58180 25998 58182
rect 26022 58180 26078 58182
rect 25962 57976 26018 58032
rect 26054 57452 26110 57488
rect 26054 57432 26056 57452
rect 26056 57432 26108 57452
rect 26108 57432 26110 57452
rect 25962 57296 26018 57352
rect 25782 57146 25838 57148
rect 25862 57146 25918 57148
rect 25942 57146 25998 57148
rect 26022 57146 26078 57148
rect 25782 57094 25828 57146
rect 25828 57094 25838 57146
rect 25862 57094 25892 57146
rect 25892 57094 25904 57146
rect 25904 57094 25918 57146
rect 25942 57094 25956 57146
rect 25956 57094 25968 57146
rect 25968 57094 25998 57146
rect 26022 57094 26032 57146
rect 26032 57094 26078 57146
rect 25782 57092 25838 57094
rect 25862 57092 25918 57094
rect 25942 57092 25998 57094
rect 26022 57092 26078 57094
rect 26054 56888 26110 56944
rect 25782 56058 25838 56060
rect 25862 56058 25918 56060
rect 25942 56058 25998 56060
rect 26022 56058 26078 56060
rect 25782 56006 25828 56058
rect 25828 56006 25838 56058
rect 25862 56006 25892 56058
rect 25892 56006 25904 56058
rect 25904 56006 25918 56058
rect 25942 56006 25956 56058
rect 25956 56006 25968 56058
rect 25968 56006 25998 56058
rect 26022 56006 26032 56058
rect 26032 56006 26078 56058
rect 25782 56004 25838 56006
rect 25862 56004 25918 56006
rect 25942 56004 25998 56006
rect 26022 56004 26078 56006
rect 25962 55820 26018 55856
rect 25962 55800 25964 55820
rect 25964 55800 26016 55820
rect 26016 55800 26018 55820
rect 25870 55392 25926 55448
rect 25778 55256 25834 55312
rect 25962 55120 26018 55176
rect 25782 54970 25838 54972
rect 25862 54970 25918 54972
rect 25942 54970 25998 54972
rect 26022 54970 26078 54972
rect 25782 54918 25828 54970
rect 25828 54918 25838 54970
rect 25862 54918 25892 54970
rect 25892 54918 25904 54970
rect 25904 54918 25918 54970
rect 25942 54918 25956 54970
rect 25956 54918 25968 54970
rect 25968 54918 25998 54970
rect 26022 54918 26032 54970
rect 26032 54918 26078 54970
rect 25782 54916 25838 54918
rect 25862 54916 25918 54918
rect 25942 54916 25998 54918
rect 26022 54916 26078 54918
rect 26422 60968 26478 61024
rect 26330 58556 26332 58576
rect 26332 58556 26384 58576
rect 26384 58556 26386 58576
rect 26330 58520 26386 58556
rect 26330 57568 26386 57624
rect 26146 54712 26202 54768
rect 26146 54304 26202 54360
rect 26054 54168 26110 54224
rect 25782 53882 25838 53884
rect 25862 53882 25918 53884
rect 25942 53882 25998 53884
rect 26022 53882 26078 53884
rect 25782 53830 25828 53882
rect 25828 53830 25838 53882
rect 25862 53830 25892 53882
rect 25892 53830 25904 53882
rect 25904 53830 25918 53882
rect 25942 53830 25956 53882
rect 25956 53830 25968 53882
rect 25968 53830 25998 53882
rect 26022 53830 26032 53882
rect 26032 53830 26078 53882
rect 25782 53828 25838 53830
rect 25862 53828 25918 53830
rect 25942 53828 25998 53830
rect 26022 53828 26078 53830
rect 25962 53080 26018 53136
rect 25782 52794 25838 52796
rect 25862 52794 25918 52796
rect 25942 52794 25998 52796
rect 26022 52794 26078 52796
rect 25782 52742 25828 52794
rect 25828 52742 25838 52794
rect 25862 52742 25892 52794
rect 25892 52742 25904 52794
rect 25904 52742 25918 52794
rect 25942 52742 25956 52794
rect 25956 52742 25968 52794
rect 25968 52742 25998 52794
rect 26022 52742 26032 52794
rect 26032 52742 26078 52794
rect 25782 52740 25838 52742
rect 25862 52740 25918 52742
rect 25942 52740 25998 52742
rect 26022 52740 26078 52742
rect 25502 48864 25558 48920
rect 25502 46452 25504 46472
rect 25504 46452 25556 46472
rect 25556 46452 25558 46472
rect 25502 46416 25558 46452
rect 25318 42336 25374 42392
rect 25318 41520 25374 41576
rect 25226 40840 25282 40896
rect 25226 40704 25282 40760
rect 25134 40432 25190 40488
rect 25226 37440 25282 37496
rect 25134 32000 25190 32056
rect 24858 31320 24914 31376
rect 24582 24792 24638 24848
rect 25134 31184 25190 31240
rect 25042 30640 25098 30696
rect 25042 28600 25098 28656
rect 24858 25336 24914 25392
rect 24950 24112 25006 24168
rect 25134 26832 25190 26888
rect 25042 22344 25098 22400
rect 24950 22072 25006 22128
rect 25042 21936 25098 21992
rect 24950 21664 25006 21720
rect 24858 18128 24914 18184
rect 25134 21392 25190 21448
rect 25502 41384 25558 41440
rect 25410 41112 25466 41168
rect 25782 51706 25838 51708
rect 25862 51706 25918 51708
rect 25942 51706 25998 51708
rect 26022 51706 26078 51708
rect 25782 51654 25828 51706
rect 25828 51654 25838 51706
rect 25862 51654 25892 51706
rect 25892 51654 25904 51706
rect 25904 51654 25918 51706
rect 25942 51654 25956 51706
rect 25956 51654 25968 51706
rect 25968 51654 25998 51706
rect 26022 51654 26032 51706
rect 26032 51654 26078 51706
rect 25782 51652 25838 51654
rect 25862 51652 25918 51654
rect 25942 51652 25998 51654
rect 26022 51652 26078 51654
rect 25778 51060 25834 51096
rect 25778 51040 25780 51060
rect 25780 51040 25832 51060
rect 25832 51040 25834 51060
rect 25778 50788 25834 50824
rect 25778 50768 25780 50788
rect 25780 50768 25832 50788
rect 25832 50768 25834 50788
rect 25782 50618 25838 50620
rect 25862 50618 25918 50620
rect 25942 50618 25998 50620
rect 26022 50618 26078 50620
rect 25782 50566 25828 50618
rect 25828 50566 25838 50618
rect 25862 50566 25892 50618
rect 25892 50566 25904 50618
rect 25904 50566 25918 50618
rect 25942 50566 25956 50618
rect 25956 50566 25968 50618
rect 25968 50566 25998 50618
rect 26022 50566 26032 50618
rect 26032 50566 26078 50618
rect 25782 50564 25838 50566
rect 25862 50564 25918 50566
rect 25942 50564 25998 50566
rect 26022 50564 26078 50566
rect 25870 50224 25926 50280
rect 25778 49972 25834 50008
rect 25778 49952 25780 49972
rect 25780 49952 25832 49972
rect 25832 49952 25834 49972
rect 25782 49530 25838 49532
rect 25862 49530 25918 49532
rect 25942 49530 25998 49532
rect 26022 49530 26078 49532
rect 25782 49478 25828 49530
rect 25828 49478 25838 49530
rect 25862 49478 25892 49530
rect 25892 49478 25904 49530
rect 25904 49478 25918 49530
rect 25942 49478 25956 49530
rect 25956 49478 25968 49530
rect 25968 49478 25998 49530
rect 26022 49478 26032 49530
rect 26032 49478 26078 49530
rect 25782 49476 25838 49478
rect 25862 49476 25918 49478
rect 25942 49476 25998 49478
rect 26022 49476 26078 49478
rect 26146 48728 26202 48784
rect 26606 61240 26662 61296
rect 26882 66816 26938 66872
rect 27250 67224 27306 67280
rect 26790 61376 26846 61432
rect 27526 68176 27582 68232
rect 27526 67768 27582 67824
rect 29274 77696 29330 77752
rect 28906 77324 28908 77344
rect 28908 77324 28960 77344
rect 28960 77324 28962 77344
rect 28906 77288 28962 77324
rect 27802 67668 27804 67688
rect 27804 67668 27856 67688
rect 27856 67668 27858 67688
rect 27802 67632 27858 67668
rect 27802 67532 27804 67552
rect 27804 67532 27856 67552
rect 27856 67532 27858 67552
rect 27802 67496 27858 67532
rect 27894 65592 27950 65648
rect 27894 64404 27896 64424
rect 27896 64404 27948 64424
rect 27948 64404 27950 64424
rect 27434 63688 27490 63744
rect 27618 63144 27674 63200
rect 27526 62872 27582 62928
rect 27250 62328 27306 62384
rect 27710 62736 27766 62792
rect 27618 62192 27674 62248
rect 26974 60968 27030 61024
rect 27158 60968 27214 61024
rect 26606 60052 26608 60072
rect 26608 60052 26660 60072
rect 26660 60052 26662 60072
rect 26606 60016 26662 60052
rect 26790 60016 26846 60072
rect 26974 60560 27030 60616
rect 27066 60288 27122 60344
rect 26606 57568 26662 57624
rect 26330 52944 26386 53000
rect 26790 55936 26846 55992
rect 26422 51176 26478 51232
rect 26606 52028 26608 52048
rect 26608 52028 26660 52048
rect 26660 52028 26662 52048
rect 26606 51992 26662 52028
rect 26330 48728 26386 48784
rect 25962 48592 26018 48648
rect 25782 48442 25838 48444
rect 25862 48442 25918 48444
rect 25942 48442 25998 48444
rect 26022 48442 26078 48444
rect 25782 48390 25828 48442
rect 25828 48390 25838 48442
rect 25862 48390 25892 48442
rect 25892 48390 25904 48442
rect 25904 48390 25918 48442
rect 25942 48390 25956 48442
rect 25956 48390 25968 48442
rect 25968 48390 25998 48442
rect 26022 48390 26032 48442
rect 26032 48390 26078 48442
rect 25782 48388 25838 48390
rect 25862 48388 25918 48390
rect 25942 48388 25998 48390
rect 26022 48388 26078 48390
rect 25962 47796 26018 47832
rect 25962 47776 25964 47796
rect 25964 47776 26016 47796
rect 26016 47776 26018 47796
rect 26330 48184 26386 48240
rect 26238 48048 26294 48104
rect 25782 47354 25838 47356
rect 25862 47354 25918 47356
rect 25942 47354 25998 47356
rect 26022 47354 26078 47356
rect 25782 47302 25828 47354
rect 25828 47302 25838 47354
rect 25862 47302 25892 47354
rect 25892 47302 25904 47354
rect 25904 47302 25918 47354
rect 25942 47302 25956 47354
rect 25956 47302 25968 47354
rect 25968 47302 25998 47354
rect 26022 47302 26032 47354
rect 26032 47302 26078 47354
rect 25782 47300 25838 47302
rect 25862 47300 25918 47302
rect 25942 47300 25998 47302
rect 26022 47300 26078 47302
rect 25778 46452 25780 46472
rect 25780 46452 25832 46472
rect 25832 46452 25834 46472
rect 25778 46416 25834 46452
rect 25782 46266 25838 46268
rect 25862 46266 25918 46268
rect 25942 46266 25998 46268
rect 26022 46266 26078 46268
rect 25782 46214 25828 46266
rect 25828 46214 25838 46266
rect 25862 46214 25892 46266
rect 25892 46214 25904 46266
rect 25904 46214 25918 46266
rect 25942 46214 25956 46266
rect 25956 46214 25968 46266
rect 25968 46214 25998 46266
rect 26022 46214 26032 46266
rect 26032 46214 26078 46266
rect 25782 46212 25838 46214
rect 25862 46212 25918 46214
rect 25942 46212 25998 46214
rect 26022 46212 26078 46214
rect 25782 45178 25838 45180
rect 25862 45178 25918 45180
rect 25942 45178 25998 45180
rect 26022 45178 26078 45180
rect 25782 45126 25828 45178
rect 25828 45126 25838 45178
rect 25862 45126 25892 45178
rect 25892 45126 25904 45178
rect 25904 45126 25918 45178
rect 25942 45126 25956 45178
rect 25956 45126 25968 45178
rect 25968 45126 25998 45178
rect 26022 45126 26032 45178
rect 26032 45126 26078 45178
rect 25782 45124 25838 45126
rect 25862 45124 25918 45126
rect 25942 45124 25998 45126
rect 26022 45124 26078 45126
rect 25782 44090 25838 44092
rect 25862 44090 25918 44092
rect 25942 44090 25998 44092
rect 26022 44090 26078 44092
rect 25782 44038 25828 44090
rect 25828 44038 25838 44090
rect 25862 44038 25892 44090
rect 25892 44038 25904 44090
rect 25904 44038 25918 44090
rect 25942 44038 25956 44090
rect 25956 44038 25968 44090
rect 25968 44038 25998 44090
rect 26022 44038 26032 44090
rect 26032 44038 26078 44090
rect 25782 44036 25838 44038
rect 25862 44036 25918 44038
rect 25942 44036 25998 44038
rect 26022 44036 26078 44038
rect 25782 43002 25838 43004
rect 25862 43002 25918 43004
rect 25942 43002 25998 43004
rect 26022 43002 26078 43004
rect 25782 42950 25828 43002
rect 25828 42950 25838 43002
rect 25862 42950 25892 43002
rect 25892 42950 25904 43002
rect 25904 42950 25918 43002
rect 25942 42950 25956 43002
rect 25956 42950 25968 43002
rect 25968 42950 25998 43002
rect 26022 42950 26032 43002
rect 26032 42950 26078 43002
rect 25782 42948 25838 42950
rect 25862 42948 25918 42950
rect 25942 42948 25998 42950
rect 26022 42948 26078 42950
rect 25870 42744 25926 42800
rect 25778 42472 25834 42528
rect 25870 42200 25926 42256
rect 25782 41914 25838 41916
rect 25862 41914 25918 41916
rect 25942 41914 25998 41916
rect 26022 41914 26078 41916
rect 25782 41862 25828 41914
rect 25828 41862 25838 41914
rect 25862 41862 25892 41914
rect 25892 41862 25904 41914
rect 25904 41862 25918 41914
rect 25942 41862 25956 41914
rect 25956 41862 25968 41914
rect 25968 41862 25998 41914
rect 26022 41862 26032 41914
rect 26032 41862 26078 41914
rect 25782 41860 25838 41862
rect 25862 41860 25918 41862
rect 25942 41860 25998 41862
rect 26022 41860 26078 41862
rect 25686 41520 25742 41576
rect 25594 38528 25650 38584
rect 25962 40976 26018 41032
rect 26974 59492 27030 59528
rect 26974 59472 26976 59492
rect 26976 59472 27028 59492
rect 27028 59472 27030 59492
rect 26974 54732 27030 54768
rect 26974 54712 26976 54732
rect 26976 54712 27028 54732
rect 27028 54712 27030 54732
rect 26882 49544 26938 49600
rect 26974 49408 27030 49464
rect 27158 60188 27160 60208
rect 27160 60188 27212 60208
rect 27212 60188 27214 60208
rect 27158 60152 27214 60188
rect 27158 58792 27214 58848
rect 27434 62056 27490 62112
rect 27342 60968 27398 61024
rect 27710 61104 27766 61160
rect 27434 57740 27436 57760
rect 27436 57740 27488 57760
rect 27488 57740 27490 57760
rect 27434 57704 27490 57740
rect 27434 57432 27490 57488
rect 27342 57160 27398 57216
rect 27342 57024 27398 57080
rect 27434 55528 27490 55584
rect 27894 64368 27950 64404
rect 27894 62092 27896 62112
rect 27896 62092 27948 62112
rect 27948 62092 27950 62112
rect 27894 62056 27950 62092
rect 27894 60968 27950 61024
rect 27618 58520 27674 58576
rect 27434 54576 27490 54632
rect 27434 54440 27490 54496
rect 27710 53216 27766 53272
rect 26790 49136 26846 49192
rect 27066 49136 27122 49192
rect 27434 49700 27490 49736
rect 27434 49680 27436 49700
rect 27436 49680 27488 49700
rect 27488 49680 27490 49700
rect 27434 49408 27490 49464
rect 27342 49000 27398 49056
rect 26790 48456 26846 48512
rect 26514 46860 26516 46880
rect 26516 46860 26568 46880
rect 26568 46860 26570 46880
rect 26514 46824 26570 46860
rect 26330 45056 26386 45112
rect 26146 41384 26202 41440
rect 25782 40826 25838 40828
rect 25862 40826 25918 40828
rect 25942 40826 25998 40828
rect 26022 40826 26078 40828
rect 25782 40774 25828 40826
rect 25828 40774 25838 40826
rect 25862 40774 25892 40826
rect 25892 40774 25904 40826
rect 25904 40774 25918 40826
rect 25942 40774 25956 40826
rect 25956 40774 25968 40826
rect 25968 40774 25998 40826
rect 26022 40774 26032 40826
rect 26032 40774 26078 40826
rect 25782 40772 25838 40774
rect 25862 40772 25918 40774
rect 25942 40772 25998 40774
rect 26022 40772 26078 40774
rect 25870 40452 25926 40488
rect 25870 40432 25872 40452
rect 25872 40432 25924 40452
rect 25924 40432 25926 40452
rect 26054 40452 26110 40488
rect 26054 40432 26056 40452
rect 26056 40432 26108 40452
rect 26108 40432 26110 40452
rect 25778 40296 25834 40352
rect 26514 41420 26516 41440
rect 26516 41420 26568 41440
rect 26568 41420 26570 41440
rect 26514 41384 26570 41420
rect 26514 41248 26570 41304
rect 26330 40432 26386 40488
rect 25782 39738 25838 39740
rect 25862 39738 25918 39740
rect 25942 39738 25998 39740
rect 26022 39738 26078 39740
rect 25782 39686 25828 39738
rect 25828 39686 25838 39738
rect 25862 39686 25892 39738
rect 25892 39686 25904 39738
rect 25904 39686 25918 39738
rect 25942 39686 25956 39738
rect 25956 39686 25968 39738
rect 25968 39686 25998 39738
rect 26022 39686 26032 39738
rect 26032 39686 26078 39738
rect 25782 39684 25838 39686
rect 25862 39684 25918 39686
rect 25942 39684 25998 39686
rect 26022 39684 26078 39686
rect 25962 39344 26018 39400
rect 26146 39480 26202 39536
rect 25870 38936 25926 38992
rect 25870 38836 25872 38856
rect 25872 38836 25924 38856
rect 25924 38836 25926 38856
rect 25870 38800 25926 38836
rect 25782 38650 25838 38652
rect 25862 38650 25918 38652
rect 25942 38650 25998 38652
rect 26022 38650 26078 38652
rect 25782 38598 25828 38650
rect 25828 38598 25838 38650
rect 25862 38598 25892 38650
rect 25892 38598 25904 38650
rect 25904 38598 25918 38650
rect 25942 38598 25956 38650
rect 25956 38598 25968 38650
rect 25968 38598 25998 38650
rect 26022 38598 26032 38650
rect 26032 38598 26078 38650
rect 25782 38596 25838 38598
rect 25862 38596 25918 38598
rect 25942 38596 25998 38598
rect 26022 38596 26078 38598
rect 25778 38392 25834 38448
rect 26054 38392 26110 38448
rect 25594 38120 25650 38176
rect 25502 37168 25558 37224
rect 25410 32816 25466 32872
rect 25782 37562 25838 37564
rect 25862 37562 25918 37564
rect 25942 37562 25998 37564
rect 26022 37562 26078 37564
rect 25782 37510 25828 37562
rect 25828 37510 25838 37562
rect 25862 37510 25892 37562
rect 25892 37510 25904 37562
rect 25904 37510 25918 37562
rect 25942 37510 25956 37562
rect 25956 37510 25968 37562
rect 25968 37510 25998 37562
rect 26022 37510 26032 37562
rect 26032 37510 26078 37562
rect 25782 37508 25838 37510
rect 25862 37508 25918 37510
rect 25942 37508 25998 37510
rect 26022 37508 26078 37510
rect 26054 37068 26056 37088
rect 26056 37068 26108 37088
rect 26108 37068 26110 37088
rect 26054 37032 26110 37068
rect 26422 39208 26478 39264
rect 26330 39072 26386 39128
rect 26698 41928 26754 41984
rect 26514 38936 26570 38992
rect 26514 38800 26570 38856
rect 26330 38664 26386 38720
rect 25686 36624 25742 36680
rect 25782 36474 25838 36476
rect 25862 36474 25918 36476
rect 25942 36474 25998 36476
rect 26022 36474 26078 36476
rect 25782 36422 25828 36474
rect 25828 36422 25838 36474
rect 25862 36422 25892 36474
rect 25892 36422 25904 36474
rect 25904 36422 25918 36474
rect 25942 36422 25956 36474
rect 25956 36422 25968 36474
rect 25968 36422 25998 36474
rect 26022 36422 26032 36474
rect 26032 36422 26078 36474
rect 25782 36420 25838 36422
rect 25862 36420 25918 36422
rect 25942 36420 25998 36422
rect 26022 36420 26078 36422
rect 25594 36080 25650 36136
rect 25870 35808 25926 35864
rect 26054 35980 26056 36000
rect 26056 35980 26108 36000
rect 26108 35980 26110 36000
rect 26054 35944 26110 35980
rect 25778 35672 25834 35728
rect 26422 38528 26478 38584
rect 26422 36624 26478 36680
rect 26606 38156 26608 38176
rect 26608 38156 26660 38176
rect 26660 38156 26662 38176
rect 26606 38120 26662 38156
rect 26698 36624 26754 36680
rect 25782 35386 25838 35388
rect 25862 35386 25918 35388
rect 25942 35386 25998 35388
rect 26022 35386 26078 35388
rect 25782 35334 25828 35386
rect 25828 35334 25838 35386
rect 25862 35334 25892 35386
rect 25892 35334 25904 35386
rect 25904 35334 25918 35386
rect 25942 35334 25956 35386
rect 25956 35334 25968 35386
rect 25968 35334 25998 35386
rect 26022 35334 26032 35386
rect 26032 35334 26078 35386
rect 25782 35332 25838 35334
rect 25862 35332 25918 35334
rect 25942 35332 25998 35334
rect 26022 35332 26078 35334
rect 25782 34298 25838 34300
rect 25862 34298 25918 34300
rect 25942 34298 25998 34300
rect 26022 34298 26078 34300
rect 25782 34246 25828 34298
rect 25828 34246 25838 34298
rect 25862 34246 25892 34298
rect 25892 34246 25904 34298
rect 25904 34246 25918 34298
rect 25942 34246 25956 34298
rect 25956 34246 25968 34298
rect 25968 34246 25998 34298
rect 26022 34246 26032 34298
rect 26032 34246 26078 34298
rect 25782 34244 25838 34246
rect 25862 34244 25918 34246
rect 25942 34244 25998 34246
rect 26022 34244 26078 34246
rect 25778 34040 25834 34096
rect 25594 31728 25650 31784
rect 25410 27104 25466 27160
rect 25594 30132 25596 30152
rect 25596 30132 25648 30152
rect 25648 30132 25650 30152
rect 25594 30096 25650 30132
rect 25782 33210 25838 33212
rect 25862 33210 25918 33212
rect 25942 33210 25998 33212
rect 26022 33210 26078 33212
rect 25782 33158 25828 33210
rect 25828 33158 25838 33210
rect 25862 33158 25892 33210
rect 25892 33158 25904 33210
rect 25904 33158 25918 33210
rect 25942 33158 25956 33210
rect 25956 33158 25968 33210
rect 25968 33158 25998 33210
rect 26022 33158 26032 33210
rect 26032 33158 26078 33210
rect 25782 33156 25838 33158
rect 25862 33156 25918 33158
rect 25942 33156 25998 33158
rect 26022 33156 26078 33158
rect 25778 32988 25780 33008
rect 25780 32988 25832 33008
rect 25832 32988 25834 33008
rect 25778 32952 25834 32988
rect 25782 32122 25838 32124
rect 25862 32122 25918 32124
rect 25942 32122 25998 32124
rect 26022 32122 26078 32124
rect 25782 32070 25828 32122
rect 25828 32070 25838 32122
rect 25862 32070 25892 32122
rect 25892 32070 25904 32122
rect 25904 32070 25918 32122
rect 25942 32070 25956 32122
rect 25956 32070 25968 32122
rect 25968 32070 25998 32122
rect 26022 32070 26032 32122
rect 26032 32070 26078 32122
rect 25782 32068 25838 32070
rect 25862 32068 25918 32070
rect 25942 32068 25998 32070
rect 26022 32068 26078 32070
rect 26054 31900 26056 31920
rect 26056 31900 26108 31920
rect 26108 31900 26110 31920
rect 26054 31864 26110 31900
rect 26238 31592 26294 31648
rect 26146 31320 26202 31376
rect 25782 31034 25838 31036
rect 25862 31034 25918 31036
rect 25942 31034 25998 31036
rect 26022 31034 26078 31036
rect 25782 30982 25828 31034
rect 25828 30982 25838 31034
rect 25862 30982 25892 31034
rect 25892 30982 25904 31034
rect 25904 30982 25918 31034
rect 25942 30982 25956 31034
rect 25956 30982 25968 31034
rect 25968 30982 25998 31034
rect 26022 30982 26032 31034
rect 26032 30982 26078 31034
rect 25782 30980 25838 30982
rect 25862 30980 25918 30982
rect 25942 30980 25998 30982
rect 26022 30980 26078 30982
rect 26054 30776 26110 30832
rect 25782 29946 25838 29948
rect 25862 29946 25918 29948
rect 25942 29946 25998 29948
rect 26022 29946 26078 29948
rect 25782 29894 25828 29946
rect 25828 29894 25838 29946
rect 25862 29894 25892 29946
rect 25892 29894 25904 29946
rect 25904 29894 25918 29946
rect 25942 29894 25956 29946
rect 25956 29894 25968 29946
rect 25968 29894 25998 29946
rect 26022 29894 26032 29946
rect 26032 29894 26078 29946
rect 25782 29892 25838 29894
rect 25862 29892 25918 29894
rect 25942 29892 25998 29894
rect 26022 29892 26078 29894
rect 25778 29688 25834 29744
rect 25962 29416 26018 29472
rect 26054 29280 26110 29336
rect 26054 29164 26110 29200
rect 26054 29144 26056 29164
rect 26056 29144 26108 29164
rect 26108 29144 26110 29164
rect 25594 27920 25650 27976
rect 25782 28858 25838 28860
rect 25862 28858 25918 28860
rect 25942 28858 25998 28860
rect 26022 28858 26078 28860
rect 25782 28806 25828 28858
rect 25828 28806 25838 28858
rect 25862 28806 25892 28858
rect 25892 28806 25904 28858
rect 25904 28806 25918 28858
rect 25942 28806 25956 28858
rect 25956 28806 25968 28858
rect 25968 28806 25998 28858
rect 26022 28806 26032 28858
rect 26032 28806 26078 28858
rect 25782 28804 25838 28806
rect 25862 28804 25918 28806
rect 25942 28804 25998 28806
rect 26022 28804 26078 28806
rect 25782 27770 25838 27772
rect 25862 27770 25918 27772
rect 25942 27770 25998 27772
rect 26022 27770 26078 27772
rect 25782 27718 25828 27770
rect 25828 27718 25838 27770
rect 25862 27718 25892 27770
rect 25892 27718 25904 27770
rect 25904 27718 25918 27770
rect 25942 27718 25956 27770
rect 25956 27718 25968 27770
rect 25968 27718 25998 27770
rect 26022 27718 26032 27770
rect 26032 27718 26078 27770
rect 25782 27716 25838 27718
rect 25862 27716 25918 27718
rect 25942 27716 25998 27718
rect 26022 27716 26078 27718
rect 25686 26968 25742 27024
rect 25318 25200 25374 25256
rect 25410 23060 25412 23080
rect 25412 23060 25464 23080
rect 25464 23060 25466 23080
rect 25410 23024 25466 23060
rect 25318 21800 25374 21856
rect 25594 22480 25650 22536
rect 25782 26682 25838 26684
rect 25862 26682 25918 26684
rect 25942 26682 25998 26684
rect 26022 26682 26078 26684
rect 25782 26630 25828 26682
rect 25828 26630 25838 26682
rect 25862 26630 25892 26682
rect 25892 26630 25904 26682
rect 25904 26630 25918 26682
rect 25942 26630 25956 26682
rect 25956 26630 25968 26682
rect 25968 26630 25998 26682
rect 26022 26630 26032 26682
rect 26032 26630 26078 26682
rect 25782 26628 25838 26630
rect 25862 26628 25918 26630
rect 25942 26628 25998 26630
rect 26022 26628 26078 26630
rect 26054 26424 26110 26480
rect 26238 26424 26294 26480
rect 25782 25594 25838 25596
rect 25862 25594 25918 25596
rect 25942 25594 25998 25596
rect 26022 25594 26078 25596
rect 25782 25542 25828 25594
rect 25828 25542 25838 25594
rect 25862 25542 25892 25594
rect 25892 25542 25904 25594
rect 25904 25542 25918 25594
rect 25942 25542 25956 25594
rect 25956 25542 25968 25594
rect 25968 25542 25998 25594
rect 26022 25542 26032 25594
rect 26032 25542 26078 25594
rect 25782 25540 25838 25542
rect 25862 25540 25918 25542
rect 25942 25540 25998 25542
rect 26022 25540 26078 25542
rect 25782 24506 25838 24508
rect 25862 24506 25918 24508
rect 25942 24506 25998 24508
rect 26022 24506 26078 24508
rect 25782 24454 25828 24506
rect 25828 24454 25838 24506
rect 25862 24454 25892 24506
rect 25892 24454 25904 24506
rect 25904 24454 25918 24506
rect 25942 24454 25956 24506
rect 25956 24454 25968 24506
rect 25968 24454 25998 24506
rect 26022 24454 26032 24506
rect 26032 24454 26078 24506
rect 25782 24452 25838 24454
rect 25862 24452 25918 24454
rect 25942 24452 25998 24454
rect 26022 24452 26078 24454
rect 25782 23418 25838 23420
rect 25862 23418 25918 23420
rect 25942 23418 25998 23420
rect 26022 23418 26078 23420
rect 25782 23366 25828 23418
rect 25828 23366 25838 23418
rect 25862 23366 25892 23418
rect 25892 23366 25904 23418
rect 25904 23366 25918 23418
rect 25942 23366 25956 23418
rect 25956 23366 25968 23418
rect 25968 23366 25998 23418
rect 26022 23366 26032 23418
rect 26032 23366 26078 23418
rect 25782 23364 25838 23366
rect 25862 23364 25918 23366
rect 25942 23364 25998 23366
rect 26022 23364 26078 23366
rect 26238 24656 26294 24712
rect 25782 22330 25838 22332
rect 25862 22330 25918 22332
rect 25942 22330 25998 22332
rect 26022 22330 26078 22332
rect 25782 22278 25828 22330
rect 25828 22278 25838 22330
rect 25862 22278 25892 22330
rect 25892 22278 25904 22330
rect 25904 22278 25918 22330
rect 25942 22278 25956 22330
rect 25956 22278 25968 22330
rect 25968 22278 25998 22330
rect 26022 22278 26032 22330
rect 26032 22278 26078 22330
rect 25782 22276 25838 22278
rect 25862 22276 25918 22278
rect 25942 22276 25998 22278
rect 26022 22276 26078 22278
rect 26238 22092 26294 22128
rect 26238 22072 26240 22092
rect 26240 22072 26292 22092
rect 26292 22072 26294 22092
rect 25782 21242 25838 21244
rect 25862 21242 25918 21244
rect 25942 21242 25998 21244
rect 26022 21242 26078 21244
rect 25782 21190 25828 21242
rect 25828 21190 25838 21242
rect 25862 21190 25892 21242
rect 25892 21190 25904 21242
rect 25904 21190 25918 21242
rect 25942 21190 25956 21242
rect 25956 21190 25968 21242
rect 25968 21190 25998 21242
rect 26022 21190 26032 21242
rect 26032 21190 26078 21242
rect 25782 21188 25838 21190
rect 25862 21188 25918 21190
rect 25942 21188 25998 21190
rect 26022 21188 26078 21190
rect 25778 20984 25834 21040
rect 25782 20154 25838 20156
rect 25862 20154 25918 20156
rect 25942 20154 25998 20156
rect 26022 20154 26078 20156
rect 25782 20102 25828 20154
rect 25828 20102 25838 20154
rect 25862 20102 25892 20154
rect 25892 20102 25904 20154
rect 25904 20102 25918 20154
rect 25942 20102 25956 20154
rect 25956 20102 25968 20154
rect 25968 20102 25998 20154
rect 26022 20102 26032 20154
rect 26032 20102 26078 20154
rect 25782 20100 25838 20102
rect 25862 20100 25918 20102
rect 25942 20100 25998 20102
rect 26022 20100 26078 20102
rect 25318 18400 25374 18456
rect 25042 16108 25098 16144
rect 25042 16088 25044 16108
rect 25044 16088 25096 16108
rect 25096 16088 25098 16108
rect 25782 19066 25838 19068
rect 25862 19066 25918 19068
rect 25942 19066 25998 19068
rect 26022 19066 26078 19068
rect 25782 19014 25828 19066
rect 25828 19014 25838 19066
rect 25862 19014 25892 19066
rect 25892 19014 25904 19066
rect 25904 19014 25918 19066
rect 25942 19014 25956 19066
rect 25956 19014 25968 19066
rect 25968 19014 25998 19066
rect 26022 19014 26032 19066
rect 26032 19014 26078 19066
rect 25782 19012 25838 19014
rect 25862 19012 25918 19014
rect 25942 19012 25998 19014
rect 26022 19012 26078 19014
rect 25962 18692 26018 18728
rect 25962 18672 25964 18692
rect 25964 18672 26016 18692
rect 26016 18672 26018 18692
rect 25778 18128 25834 18184
rect 25782 17978 25838 17980
rect 25862 17978 25918 17980
rect 25942 17978 25998 17980
rect 26022 17978 26078 17980
rect 25782 17926 25828 17978
rect 25828 17926 25838 17978
rect 25862 17926 25892 17978
rect 25892 17926 25904 17978
rect 25904 17926 25918 17978
rect 25942 17926 25956 17978
rect 25956 17926 25968 17978
rect 25968 17926 25998 17978
rect 26022 17926 26032 17978
rect 26032 17926 26078 17978
rect 25782 17924 25838 17926
rect 25862 17924 25918 17926
rect 25942 17924 25998 17926
rect 26022 17924 26078 17926
rect 26054 17620 26056 17640
rect 26056 17620 26108 17640
rect 26108 17620 26110 17640
rect 26054 17584 26110 17620
rect 25594 15272 25650 15328
rect 25782 16890 25838 16892
rect 25862 16890 25918 16892
rect 25942 16890 25998 16892
rect 26022 16890 26078 16892
rect 25782 16838 25828 16890
rect 25828 16838 25838 16890
rect 25862 16838 25892 16890
rect 25892 16838 25904 16890
rect 25904 16838 25918 16890
rect 25942 16838 25956 16890
rect 25956 16838 25968 16890
rect 25968 16838 25998 16890
rect 26022 16838 26032 16890
rect 26032 16838 26078 16890
rect 25782 16836 25838 16838
rect 25862 16836 25918 16838
rect 25942 16836 25998 16838
rect 26022 16836 26078 16838
rect 25782 15802 25838 15804
rect 25862 15802 25918 15804
rect 25942 15802 25998 15804
rect 26022 15802 26078 15804
rect 25782 15750 25828 15802
rect 25828 15750 25838 15802
rect 25862 15750 25892 15802
rect 25892 15750 25904 15802
rect 25904 15750 25918 15802
rect 25942 15750 25956 15802
rect 25956 15750 25968 15802
rect 25968 15750 25998 15802
rect 26022 15750 26032 15802
rect 26032 15750 26078 15802
rect 25782 15748 25838 15750
rect 25862 15748 25918 15750
rect 25942 15748 25998 15750
rect 26022 15748 26078 15750
rect 25782 14714 25838 14716
rect 25862 14714 25918 14716
rect 25942 14714 25998 14716
rect 26022 14714 26078 14716
rect 25782 14662 25828 14714
rect 25828 14662 25838 14714
rect 25862 14662 25892 14714
rect 25892 14662 25904 14714
rect 25904 14662 25918 14714
rect 25942 14662 25956 14714
rect 25956 14662 25968 14714
rect 25968 14662 25998 14714
rect 26022 14662 26032 14714
rect 26032 14662 26078 14714
rect 25782 14660 25838 14662
rect 25862 14660 25918 14662
rect 25942 14660 25998 14662
rect 26022 14660 26078 14662
rect 25778 14048 25834 14104
rect 26606 36352 26662 36408
rect 26514 36252 26516 36272
rect 26516 36252 26568 36272
rect 26568 36252 26570 36272
rect 26514 36216 26570 36252
rect 26422 20712 26478 20768
rect 25782 13626 25838 13628
rect 25862 13626 25918 13628
rect 25942 13626 25998 13628
rect 26022 13626 26078 13628
rect 25782 13574 25828 13626
rect 25828 13574 25838 13626
rect 25862 13574 25892 13626
rect 25892 13574 25904 13626
rect 25904 13574 25918 13626
rect 25942 13574 25956 13626
rect 25956 13574 25968 13626
rect 25968 13574 25998 13626
rect 26022 13574 26032 13626
rect 26032 13574 26078 13626
rect 25782 13572 25838 13574
rect 25862 13572 25918 13574
rect 25942 13572 25998 13574
rect 26022 13572 26078 13574
rect 25782 12538 25838 12540
rect 25862 12538 25918 12540
rect 25942 12538 25998 12540
rect 26022 12538 26078 12540
rect 25782 12486 25828 12538
rect 25828 12486 25838 12538
rect 25862 12486 25892 12538
rect 25892 12486 25904 12538
rect 25904 12486 25918 12538
rect 25942 12486 25956 12538
rect 25956 12486 25968 12538
rect 25968 12486 25998 12538
rect 26022 12486 26032 12538
rect 26032 12486 26078 12538
rect 25782 12484 25838 12486
rect 25862 12484 25918 12486
rect 25942 12484 25998 12486
rect 26022 12484 26078 12486
rect 26146 12008 26202 12064
rect 25782 11450 25838 11452
rect 25862 11450 25918 11452
rect 25942 11450 25998 11452
rect 26022 11450 26078 11452
rect 25782 11398 25828 11450
rect 25828 11398 25838 11450
rect 25862 11398 25892 11450
rect 25892 11398 25904 11450
rect 25904 11398 25918 11450
rect 25942 11398 25956 11450
rect 25956 11398 25968 11450
rect 25968 11398 25998 11450
rect 26022 11398 26032 11450
rect 26032 11398 26078 11450
rect 25782 11396 25838 11398
rect 25862 11396 25918 11398
rect 25942 11396 25998 11398
rect 26022 11396 26078 11398
rect 25782 10362 25838 10364
rect 25862 10362 25918 10364
rect 25942 10362 25998 10364
rect 26022 10362 26078 10364
rect 25782 10310 25828 10362
rect 25828 10310 25838 10362
rect 25862 10310 25892 10362
rect 25892 10310 25904 10362
rect 25904 10310 25918 10362
rect 25942 10310 25956 10362
rect 25956 10310 25968 10362
rect 25968 10310 25998 10362
rect 26022 10310 26032 10362
rect 26032 10310 26078 10362
rect 25782 10308 25838 10310
rect 25862 10308 25918 10310
rect 25942 10308 25998 10310
rect 26022 10308 26078 10310
rect 25782 9274 25838 9276
rect 25862 9274 25918 9276
rect 25942 9274 25998 9276
rect 26022 9274 26078 9276
rect 25782 9222 25828 9274
rect 25828 9222 25838 9274
rect 25862 9222 25892 9274
rect 25892 9222 25904 9274
rect 25904 9222 25918 9274
rect 25942 9222 25956 9274
rect 25956 9222 25968 9274
rect 25968 9222 25998 9274
rect 26022 9222 26032 9274
rect 26032 9222 26078 9274
rect 25782 9220 25838 9222
rect 25862 9220 25918 9222
rect 25942 9220 25998 9222
rect 26022 9220 26078 9222
rect 26514 19760 26570 19816
rect 26514 19624 26570 19680
rect 26882 48272 26938 48328
rect 26882 41520 26938 41576
rect 27066 48592 27122 48648
rect 27066 48456 27122 48512
rect 26974 41112 27030 41168
rect 27618 52536 27674 52592
rect 27618 52400 27674 52456
rect 28078 65456 28134 65512
rect 28078 64948 28080 64968
rect 28080 64948 28132 64968
rect 28132 64948 28134 64968
rect 28078 64912 28134 64948
rect 28170 64096 28226 64152
rect 28446 65592 28502 65648
rect 28262 63960 28318 64016
rect 28078 63860 28080 63880
rect 28080 63860 28132 63880
rect 28132 63860 28134 63880
rect 28078 63824 28134 63860
rect 28078 60968 28134 61024
rect 27894 53760 27950 53816
rect 28078 60152 28134 60208
rect 28078 59628 28134 59664
rect 28078 59608 28080 59628
rect 28080 59608 28132 59628
rect 28132 59608 28134 59628
rect 28078 59472 28134 59528
rect 27802 51176 27858 51232
rect 27710 51040 27766 51096
rect 27618 48728 27674 48784
rect 27434 48456 27490 48512
rect 27250 48048 27306 48104
rect 27342 47912 27398 47968
rect 26974 32136 27030 32192
rect 27158 33496 27214 33552
rect 26790 30368 26846 30424
rect 26790 29688 26846 29744
rect 26974 31728 27030 31784
rect 27066 29824 27122 29880
rect 27618 48272 27674 48328
rect 27434 44376 27490 44432
rect 27434 42336 27490 42392
rect 27986 52808 28042 52864
rect 27986 52672 28042 52728
rect 27986 50904 28042 50960
rect 27986 49544 28042 49600
rect 27802 44648 27858 44704
rect 27710 42608 27766 42664
rect 27618 42200 27674 42256
rect 27526 41656 27582 41712
rect 27802 41928 27858 41984
rect 27710 41112 27766 41168
rect 27526 40976 27582 41032
rect 27710 40976 27766 41032
rect 27618 39616 27674 39672
rect 26790 25200 26846 25256
rect 26698 22752 26754 22808
rect 26882 24928 26938 24984
rect 26790 22072 26846 22128
rect 26882 21936 26938 21992
rect 26606 17584 26662 17640
rect 26790 14048 26846 14104
rect 26514 10784 26570 10840
rect 26790 10784 26846 10840
rect 25782 8186 25838 8188
rect 25862 8186 25918 8188
rect 25942 8186 25998 8188
rect 26022 8186 26078 8188
rect 25782 8134 25828 8186
rect 25828 8134 25838 8186
rect 25862 8134 25892 8186
rect 25892 8134 25904 8186
rect 25904 8134 25918 8186
rect 25942 8134 25956 8186
rect 25956 8134 25968 8186
rect 25968 8134 25998 8186
rect 26022 8134 26032 8186
rect 26032 8134 26078 8186
rect 25782 8132 25838 8134
rect 25862 8132 25918 8134
rect 25942 8132 25998 8134
rect 26022 8132 26078 8134
rect 25782 7098 25838 7100
rect 25862 7098 25918 7100
rect 25942 7098 25998 7100
rect 26022 7098 26078 7100
rect 25782 7046 25828 7098
rect 25828 7046 25838 7098
rect 25862 7046 25892 7098
rect 25892 7046 25904 7098
rect 25904 7046 25918 7098
rect 25942 7046 25956 7098
rect 25956 7046 25968 7098
rect 25968 7046 25998 7098
rect 26022 7046 26032 7098
rect 26032 7046 26078 7098
rect 25782 7044 25838 7046
rect 25862 7044 25918 7046
rect 25942 7044 25998 7046
rect 26022 7044 26078 7046
rect 25782 6010 25838 6012
rect 25862 6010 25918 6012
rect 25942 6010 25998 6012
rect 26022 6010 26078 6012
rect 25782 5958 25828 6010
rect 25828 5958 25838 6010
rect 25862 5958 25892 6010
rect 25892 5958 25904 6010
rect 25904 5958 25918 6010
rect 25942 5958 25956 6010
rect 25956 5958 25968 6010
rect 25968 5958 25998 6010
rect 26022 5958 26032 6010
rect 26032 5958 26078 6010
rect 25782 5956 25838 5958
rect 25862 5956 25918 5958
rect 25942 5956 25998 5958
rect 26022 5956 26078 5958
rect 27342 29960 27398 30016
rect 27250 29044 27252 29064
rect 27252 29044 27304 29064
rect 27304 29044 27306 29064
rect 27250 29008 27306 29044
rect 27250 27920 27306 27976
rect 27526 35672 27582 35728
rect 27618 35436 27620 35456
rect 27620 35436 27672 35456
rect 27672 35436 27674 35456
rect 27618 35400 27674 35436
rect 27618 32408 27674 32464
rect 27986 44512 28042 44568
rect 27986 43152 28042 43208
rect 28354 63008 28410 63064
rect 29274 75792 29330 75848
rect 29182 69944 29238 70000
rect 28906 68720 28962 68776
rect 28906 67360 28962 67416
rect 28630 64504 28686 64560
rect 28538 63436 28594 63472
rect 28538 63416 28540 63436
rect 28540 63416 28592 63436
rect 28592 63416 28594 63436
rect 28538 63008 28594 63064
rect 28538 62892 28594 62928
rect 28538 62872 28540 62892
rect 28540 62872 28592 62892
rect 28592 62872 28594 62892
rect 28446 61240 28502 61296
rect 28630 61784 28686 61840
rect 28906 66408 28962 66464
rect 28814 64096 28870 64152
rect 28630 61648 28686 61704
rect 28722 61512 28778 61568
rect 28538 60968 28594 61024
rect 28538 60288 28594 60344
rect 28814 61376 28870 61432
rect 28814 61276 28816 61296
rect 28816 61276 28868 61296
rect 28868 61276 28870 61296
rect 28814 61240 28870 61276
rect 28814 61140 28816 61160
rect 28816 61140 28868 61160
rect 28868 61140 28870 61160
rect 28814 61104 28870 61140
rect 28814 60560 28870 60616
rect 28814 60016 28870 60072
rect 28170 57024 28226 57080
rect 28170 56652 28172 56672
rect 28172 56652 28224 56672
rect 28224 56652 28226 56672
rect 28170 56616 28226 56652
rect 28170 56480 28226 56536
rect 28170 51040 28226 51096
rect 28354 56752 28410 56808
rect 28446 51856 28502 51912
rect 28262 48884 28318 48920
rect 28262 48864 28264 48884
rect 28264 48864 28316 48884
rect 28316 48864 28318 48884
rect 28262 48748 28318 48784
rect 28262 48728 28264 48748
rect 28264 48728 28316 48748
rect 28316 48728 28318 48748
rect 28170 41656 28226 41712
rect 28078 41384 28134 41440
rect 28262 41384 28318 41440
rect 27986 40976 28042 41032
rect 27986 40840 28042 40896
rect 27802 40160 27858 40216
rect 27802 40024 27858 40080
rect 27710 32272 27766 32328
rect 27710 32000 27766 32056
rect 27618 31728 27674 31784
rect 27526 30912 27582 30968
rect 27526 30776 27582 30832
rect 28170 39924 28172 39944
rect 28172 39924 28224 39944
rect 28224 39924 28226 39944
rect 28170 39888 28226 39924
rect 27986 38392 28042 38448
rect 27986 37304 28042 37360
rect 28170 39244 28172 39264
rect 28172 39244 28224 39264
rect 28224 39244 28226 39264
rect 28170 39208 28226 39244
rect 28170 38256 28226 38312
rect 28262 37168 28318 37224
rect 28262 36916 28318 36952
rect 28262 36896 28264 36916
rect 28264 36896 28316 36916
rect 28316 36896 28318 36916
rect 28262 35692 28318 35728
rect 28262 35672 28264 35692
rect 28264 35672 28316 35692
rect 28316 35672 28318 35692
rect 28170 34856 28226 34912
rect 28078 32680 28134 32736
rect 28078 32544 28134 32600
rect 28078 32272 28134 32328
rect 28630 59220 28686 59256
rect 28630 59200 28632 59220
rect 28632 59200 28684 59220
rect 28684 59200 28686 59220
rect 28630 58948 28686 58984
rect 28630 58928 28632 58948
rect 28632 58928 28684 58948
rect 28684 58928 28686 58948
rect 28630 58676 28686 58712
rect 28630 58656 28632 58676
rect 28632 58656 28684 58676
rect 28684 58656 28686 58676
rect 28722 57160 28778 57216
rect 28722 56888 28778 56944
rect 28630 56072 28686 56128
rect 28906 59336 28962 59392
rect 28906 58792 28962 58848
rect 28814 55528 28870 55584
rect 28722 55392 28778 55448
rect 28814 55276 28870 55312
rect 28814 55256 28816 55276
rect 28816 55256 28868 55276
rect 28868 55256 28870 55276
rect 28814 55120 28870 55176
rect 28630 54168 28686 54224
rect 28630 52672 28686 52728
rect 28722 52264 28778 52320
rect 28630 52128 28686 52184
rect 28722 51992 28778 52048
rect 28722 51856 28778 51912
rect 28630 51312 28686 51368
rect 30102 76744 30158 76800
rect 29274 69284 29330 69320
rect 29274 69264 29276 69284
rect 29276 69264 29328 69284
rect 29328 69264 29330 69284
rect 29090 61140 29092 61160
rect 29092 61140 29144 61160
rect 29144 61140 29146 61160
rect 29090 61104 29146 61140
rect 29274 60832 29330 60888
rect 29182 60696 29238 60752
rect 30010 76336 30066 76392
rect 30010 74840 30066 74896
rect 30010 74024 30066 74080
rect 30010 73072 30066 73128
rect 30010 72528 30066 72584
rect 30010 72120 30066 72176
rect 30010 71576 30066 71632
rect 30010 71168 30066 71224
rect 30010 70624 30066 70680
rect 30010 70252 30012 70272
rect 30012 70252 30064 70272
rect 30064 70252 30066 70272
rect 30010 70216 30066 70252
rect 30010 69708 30012 69728
rect 30012 69708 30064 69728
rect 30064 69708 30066 69728
rect 30010 69672 30066 69708
rect 29918 68312 29974 68368
rect 30010 67904 30066 67960
rect 29918 66952 29974 67008
rect 30194 75384 30250 75440
rect 30194 74432 30250 74488
rect 30194 73480 30250 73536
rect 30010 66000 30066 66056
rect 29826 65048 29882 65104
rect 29918 63552 29974 63608
rect 29734 61240 29790 61296
rect 29642 61104 29698 61160
rect 29090 60560 29146 60616
rect 29182 55528 29238 55584
rect 29182 53488 29238 53544
rect 29090 53388 29092 53408
rect 29092 53388 29144 53408
rect 29144 53388 29146 53408
rect 29090 53352 29146 53388
rect 29366 60424 29422 60480
rect 29366 60152 29422 60208
rect 29366 56616 29422 56672
rect 28906 52944 28962 53000
rect 29274 53080 29330 53136
rect 29274 52672 29330 52728
rect 29458 54032 29514 54088
rect 29366 52536 29422 52592
rect 28538 45464 28594 45520
rect 28906 51212 28908 51232
rect 28908 51212 28960 51232
rect 28960 51212 28962 51232
rect 28906 51176 28962 51212
rect 29182 52128 29238 52184
rect 29090 51992 29146 52048
rect 29458 52400 29514 52456
rect 29182 51176 29238 51232
rect 28722 49816 28778 49872
rect 28814 49000 28870 49056
rect 28814 48592 28870 48648
rect 28722 48184 28778 48240
rect 28722 48048 28778 48104
rect 29090 51040 29146 51096
rect 28998 50360 29054 50416
rect 28998 47948 29000 47968
rect 29000 47948 29052 47968
rect 29052 47948 29054 47968
rect 28998 47912 29054 47948
rect 28906 45872 28962 45928
rect 28814 44784 28870 44840
rect 28722 44376 28778 44432
rect 28538 41384 28594 41440
rect 28538 41112 28594 41168
rect 28906 44240 28962 44296
rect 28906 44104 28962 44160
rect 29090 45600 29146 45656
rect 29090 45464 29146 45520
rect 28998 43288 29054 43344
rect 29826 60832 29882 60888
rect 30010 60968 30066 61024
rect 29826 59744 29882 59800
rect 29826 58384 29882 58440
rect 29734 57976 29790 58032
rect 29734 57840 29790 57896
rect 29734 57452 29790 57488
rect 29734 57432 29736 57452
rect 29736 57432 29788 57452
rect 29788 57432 29790 57452
rect 29734 57160 29790 57216
rect 29734 55120 29790 55176
rect 29734 54712 29790 54768
rect 29734 53760 29790 53816
rect 29642 53624 29698 53680
rect 29918 56616 29974 56672
rect 29918 55256 29974 55312
rect 29642 52944 29698 53000
rect 29550 51720 29606 51776
rect 29366 51312 29422 51368
rect 29366 43288 29422 43344
rect 29274 43152 29330 43208
rect 29274 42880 29330 42936
rect 29734 51448 29790 51504
rect 29642 51312 29698 51368
rect 29550 48320 29606 48376
rect 29550 48184 29606 48240
rect 30010 53100 30066 53136
rect 30010 53080 30012 53100
rect 30012 53080 30064 53100
rect 30064 53080 30066 53100
rect 29918 51584 29974 51640
rect 29918 50768 29974 50824
rect 30286 55256 30342 55312
rect 30286 54440 30342 54496
rect 29826 50668 29828 50688
rect 29828 50668 29880 50688
rect 29880 50668 29882 50688
rect 29826 50632 29882 50668
rect 29734 50360 29790 50416
rect 29826 50124 29828 50144
rect 29828 50124 29880 50144
rect 29880 50124 29882 50144
rect 29826 50088 29882 50124
rect 29734 49952 29790 50008
rect 29734 49408 29790 49464
rect 29734 47096 29790 47152
rect 29734 46688 29790 46744
rect 29734 46144 29790 46200
rect 29734 46008 29790 46064
rect 29642 45600 29698 45656
rect 29182 42200 29238 42256
rect 29090 41928 29146 41984
rect 28722 41384 28778 41440
rect 28906 41112 28962 41168
rect 28814 40976 28870 41032
rect 28630 40840 28686 40896
rect 28538 39752 28594 39808
rect 28078 31728 28134 31784
rect 28078 31320 28134 31376
rect 28446 31456 28502 31512
rect 28262 29996 28264 30016
rect 28264 29996 28316 30016
rect 28316 29996 28318 30016
rect 28262 29960 28318 29996
rect 27526 29280 27582 29336
rect 27526 28736 27582 28792
rect 27158 26968 27214 27024
rect 27066 19760 27122 19816
rect 27250 26832 27306 26888
rect 27434 26696 27490 26752
rect 27434 26560 27490 26616
rect 27250 21800 27306 21856
rect 27710 27940 27766 27976
rect 27710 27920 27712 27940
rect 27712 27920 27764 27940
rect 27764 27920 27766 27940
rect 27710 27532 27766 27568
rect 27710 27512 27712 27532
rect 27712 27512 27764 27532
rect 27764 27512 27766 27532
rect 27710 27376 27766 27432
rect 27894 29552 27950 29608
rect 28078 29416 28134 29472
rect 27894 28872 27950 28928
rect 27618 25220 27674 25256
rect 27618 25200 27620 25220
rect 27620 25200 27672 25220
rect 27672 25200 27674 25220
rect 27802 24012 27804 24032
rect 27804 24012 27856 24032
rect 27856 24012 27858 24032
rect 27802 23976 27858 24012
rect 27802 23704 27858 23760
rect 27434 22208 27490 22264
rect 27526 22072 27582 22128
rect 27342 18264 27398 18320
rect 27802 21956 27858 21992
rect 27802 21936 27804 21956
rect 27804 21936 27856 21956
rect 27856 21936 27858 21956
rect 27618 21256 27674 21312
rect 27526 18672 27582 18728
rect 27618 16224 27674 16280
rect 27618 15428 27674 15464
rect 27618 15408 27620 15428
rect 27620 15408 27672 15428
rect 27672 15408 27674 15428
rect 25782 4922 25838 4924
rect 25862 4922 25918 4924
rect 25942 4922 25998 4924
rect 26022 4922 26078 4924
rect 25782 4870 25828 4922
rect 25828 4870 25838 4922
rect 25862 4870 25892 4922
rect 25892 4870 25904 4922
rect 25904 4870 25918 4922
rect 25942 4870 25956 4922
rect 25956 4870 25968 4922
rect 25968 4870 25998 4922
rect 26022 4870 26032 4922
rect 26032 4870 26078 4922
rect 25782 4868 25838 4870
rect 25862 4868 25918 4870
rect 25942 4868 25998 4870
rect 26022 4868 26078 4870
rect 25782 3834 25838 3836
rect 25862 3834 25918 3836
rect 25942 3834 25998 3836
rect 26022 3834 26078 3836
rect 25782 3782 25828 3834
rect 25828 3782 25838 3834
rect 25862 3782 25892 3834
rect 25892 3782 25904 3834
rect 25904 3782 25918 3834
rect 25942 3782 25956 3834
rect 25956 3782 25968 3834
rect 25968 3782 25998 3834
rect 26022 3782 26032 3834
rect 26032 3782 26078 3834
rect 25782 3780 25838 3782
rect 25862 3780 25918 3782
rect 25942 3780 25998 3782
rect 26022 3780 26078 3782
rect 27618 13776 27674 13832
rect 28354 29688 28410 29744
rect 28170 29144 28226 29200
rect 28446 27412 28448 27432
rect 28448 27412 28500 27432
rect 28500 27412 28502 27432
rect 28446 27376 28502 27412
rect 28354 25064 28410 25120
rect 28078 21800 28134 21856
rect 27894 16224 27950 16280
rect 28262 20884 28264 20904
rect 28264 20884 28316 20904
rect 28316 20884 28318 20904
rect 28262 20848 28318 20884
rect 28446 22072 28502 22128
rect 28446 21800 28502 21856
rect 27986 14492 27988 14512
rect 27988 14492 28040 14512
rect 28040 14492 28042 14512
rect 27986 14456 28042 14492
rect 28354 17448 28410 17504
rect 28262 15156 28318 15192
rect 28262 15136 28264 15156
rect 28264 15136 28316 15156
rect 28316 15136 28318 15156
rect 28630 38256 28686 38312
rect 28630 37984 28686 38040
rect 28998 40840 29054 40896
rect 28906 38664 28962 38720
rect 28722 37712 28778 37768
rect 28906 34448 28962 34504
rect 28722 32680 28778 32736
rect 28906 33496 28962 33552
rect 28814 32544 28870 32600
rect 28630 32000 28686 32056
rect 28998 32544 29054 32600
rect 29366 42608 29422 42664
rect 29826 43832 29882 43888
rect 30102 48320 30158 48376
rect 30010 44532 30066 44568
rect 30010 44512 30012 44532
rect 30012 44512 30064 44532
rect 30064 44512 30066 44532
rect 30010 44260 30066 44296
rect 30010 44240 30012 44260
rect 30012 44240 30064 44260
rect 30064 44240 30066 44260
rect 29918 43560 29974 43616
rect 29826 43424 29882 43480
rect 29642 42608 29698 42664
rect 29550 42336 29606 42392
rect 29458 42064 29514 42120
rect 29734 42200 29790 42256
rect 29550 41112 29606 41168
rect 29550 40976 29606 41032
rect 29458 38120 29514 38176
rect 29366 37304 29422 37360
rect 30010 42744 30066 42800
rect 29918 42472 29974 42528
rect 30010 42064 30066 42120
rect 29734 41384 29790 41440
rect 30010 41384 30066 41440
rect 29642 40432 29698 40488
rect 29274 33088 29330 33144
rect 28906 32136 28962 32192
rect 28998 32000 29054 32056
rect 28998 31864 29054 31920
rect 28814 30776 28870 30832
rect 28630 27376 28686 27432
rect 28630 25880 28686 25936
rect 28906 30368 28962 30424
rect 28906 28464 28962 28520
rect 29182 32272 29238 32328
rect 28722 23840 28778 23896
rect 28630 23568 28686 23624
rect 28998 27784 29054 27840
rect 28906 26560 28962 26616
rect 28906 26016 28962 26072
rect 28906 25880 28962 25936
rect 29090 25744 29146 25800
rect 28998 24520 29054 24576
rect 28906 24148 28908 24168
rect 28908 24148 28960 24168
rect 28960 24148 28962 24168
rect 28906 24112 28962 24148
rect 29182 23160 29238 23216
rect 28906 22344 28962 22400
rect 28906 21800 28962 21856
rect 28722 19760 28778 19816
rect 28538 14048 28594 14104
rect 28906 20304 28962 20360
rect 28814 19352 28870 19408
rect 28998 18128 29054 18184
rect 28814 17040 28870 17096
rect 28906 16632 28962 16688
rect 28170 11872 28226 11928
rect 27710 7656 27766 7712
rect 27618 7112 27674 7168
rect 25782 2746 25838 2748
rect 25862 2746 25918 2748
rect 25942 2746 25998 2748
rect 26022 2746 26078 2748
rect 25782 2694 25828 2746
rect 25828 2694 25838 2746
rect 25862 2694 25892 2746
rect 25892 2694 25904 2746
rect 25904 2694 25918 2746
rect 25942 2694 25956 2746
rect 25956 2694 25968 2746
rect 25968 2694 25998 2746
rect 26022 2694 26032 2746
rect 26032 2694 26078 2746
rect 25782 2692 25838 2694
rect 25862 2692 25918 2694
rect 25942 2692 25998 2694
rect 26022 2692 26078 2694
rect 27802 4392 27858 4448
rect 29366 32292 29422 32328
rect 29366 32272 29368 32292
rect 29368 32272 29420 32292
rect 29420 32272 29422 32292
rect 29550 31320 29606 31376
rect 29550 30504 29606 30560
rect 29550 29824 29606 29880
rect 29458 29008 29514 29064
rect 29366 28056 29422 28112
rect 29918 40976 29974 41032
rect 30286 41520 30342 41576
rect 29826 36780 29882 36816
rect 29826 36760 29828 36780
rect 29828 36760 29880 36780
rect 29880 36760 29882 36780
rect 30010 37712 30066 37768
rect 30010 36760 30066 36816
rect 30010 36624 30066 36680
rect 29918 36488 29974 36544
rect 29918 36252 29920 36272
rect 29920 36252 29972 36272
rect 29972 36252 29974 36272
rect 29918 36216 29974 36252
rect 30194 35808 30250 35864
rect 30654 57196 30656 57216
rect 30656 57196 30708 57216
rect 30708 57196 30710 57216
rect 30654 57160 30710 57196
rect 30470 52128 30526 52184
rect 30470 50904 30526 50960
rect 30470 50632 30526 50688
rect 30930 54984 30986 55040
rect 30930 51176 30986 51232
rect 30654 44104 30710 44160
rect 30654 43288 30710 43344
rect 30562 42200 30618 42256
rect 30102 34176 30158 34232
rect 30010 34040 30066 34096
rect 29918 32680 29974 32736
rect 30010 32544 30066 32600
rect 29734 31728 29790 31784
rect 29274 19896 29330 19952
rect 29642 22072 29698 22128
rect 28906 14184 28962 14240
rect 28814 12824 28870 12880
rect 28998 13232 29054 13288
rect 28906 12280 28962 12336
rect 28722 9560 28778 9616
rect 30102 31864 30158 31920
rect 30102 30640 30158 30696
rect 30010 30232 30066 30288
rect 30010 28736 30066 28792
rect 30010 26968 30066 27024
rect 30010 25492 30066 25528
rect 30010 25472 30012 25492
rect 30012 25472 30064 25492
rect 30064 25472 30066 25492
rect 29918 22752 29974 22808
rect 30102 24792 30158 24848
rect 30286 31048 30342 31104
rect 30378 30776 30434 30832
rect 30286 22480 30342 22536
rect 30102 22072 30158 22128
rect 29826 18400 29882 18456
rect 30010 18944 30066 19000
rect 29918 17992 29974 18048
rect 30102 16088 30158 16144
rect 29918 15680 29974 15736
rect 29918 15136 29974 15192
rect 29826 14728 29882 14784
rect 29366 11464 29422 11520
rect 29274 10920 29330 10976
rect 28906 9016 28962 9072
rect 28906 8608 28962 8664
rect 29918 10512 29974 10568
rect 29734 9988 29790 10024
rect 29734 9968 29736 9988
rect 29736 9968 29788 9988
rect 29788 9968 29790 9988
rect 28814 6704 28870 6760
rect 29826 8064 29882 8120
rect 30746 41656 30802 41712
rect 30654 40704 30710 40760
rect 30930 50904 30986 50960
rect 30930 50496 30986 50552
rect 30930 49272 30986 49328
rect 30930 47232 30986 47288
rect 31390 63824 31446 63880
rect 31114 46416 31170 46472
rect 30838 41520 30894 41576
rect 30562 31184 30618 31240
rect 30562 30912 30618 30968
rect 30838 32000 30894 32056
rect 31298 51176 31354 51232
rect 31298 50224 31354 50280
rect 31390 46416 31446 46472
rect 31390 37032 31446 37088
rect 31298 36080 31354 36136
rect 31482 30912 31538 30968
rect 31850 45056 31906 45112
rect 31850 37984 31906 38040
rect 31758 31864 31814 31920
rect 29826 6452 29882 6488
rect 29826 6432 29828 6452
rect 29828 6432 29880 6452
rect 29880 6432 29882 6452
rect 30102 6160 30158 6216
rect 29826 5364 29882 5400
rect 29826 5344 29828 5364
rect 29828 5344 29880 5364
rect 29880 5344 29882 5364
rect 28170 4800 28226 4856
rect 28722 4684 28778 4720
rect 28722 4664 28724 4684
rect 28724 4664 28776 4684
rect 28776 4664 28778 4684
rect 28170 3848 28226 3904
rect 29826 4020 29828 4040
rect 29828 4020 29880 4040
rect 29880 4020 29882 4040
rect 29826 3984 29882 4020
rect 28262 3476 28264 3496
rect 28264 3476 28316 3496
rect 28316 3476 28318 3496
rect 28262 3440 28318 3476
rect 2870 312 2926 368
rect 28722 1944 28778 2000
rect 28906 2896 28962 2952
rect 29734 2488 29790 2544
rect 28814 1536 28870 1592
rect 29642 992 29698 1048
rect 28722 584 28778 640
rect 28262 176 28318 232
<< metal3 >>
rect 0 79658 800 79688
rect 3785 79658 3851 79661
rect 0 79656 3851 79658
rect 0 79600 3790 79656
rect 3846 79600 3851 79656
rect 0 79598 3851 79600
rect 0 79568 800 79598
rect 3785 79595 3851 79598
rect 27889 79658 27955 79661
rect 31200 79658 32000 79688
rect 27889 79656 32000 79658
rect 27889 79600 27894 79656
rect 27950 79600 32000 79656
rect 27889 79598 32000 79600
rect 27889 79595 27955 79598
rect 31200 79568 32000 79598
rect 28809 79250 28875 79253
rect 31200 79250 32000 79280
rect 28809 79248 32000 79250
rect 28809 79192 28814 79248
rect 28870 79192 32000 79248
rect 28809 79190 32000 79192
rect 28809 79187 28875 79190
rect 31200 79160 32000 79190
rect 0 78978 800 79008
rect 2773 78978 2839 78981
rect 0 78976 2839 78978
rect 0 78920 2778 78976
rect 2834 78920 2839 78976
rect 0 78918 2839 78920
rect 0 78888 800 78918
rect 2773 78915 2839 78918
rect 28533 78706 28599 78709
rect 31200 78706 32000 78736
rect 28533 78704 32000 78706
rect 28533 78648 28538 78704
rect 28594 78648 32000 78704
rect 28533 78646 32000 78648
rect 28533 78643 28599 78646
rect 31200 78616 32000 78646
rect 0 78298 800 78328
rect 1301 78298 1367 78301
rect 0 78296 1367 78298
rect 0 78240 1306 78296
rect 1362 78240 1367 78296
rect 0 78238 1367 78240
rect 0 78208 800 78238
rect 1301 78235 1367 78238
rect 28165 78298 28231 78301
rect 31200 78298 32000 78328
rect 28165 78296 32000 78298
rect 28165 78240 28170 78296
rect 28226 78240 32000 78296
rect 28165 78238 32000 78240
rect 28165 78235 28231 78238
rect 31200 78208 32000 78238
rect 5909 77824 6229 77825
rect 5909 77760 5917 77824
rect 5981 77760 5997 77824
rect 6061 77760 6077 77824
rect 6141 77760 6157 77824
rect 6221 77760 6229 77824
rect 5909 77759 6229 77760
rect 15840 77824 16160 77825
rect 15840 77760 15848 77824
rect 15912 77760 15928 77824
rect 15992 77760 16008 77824
rect 16072 77760 16088 77824
rect 16152 77760 16160 77824
rect 15840 77759 16160 77760
rect 25770 77824 26090 77825
rect 25770 77760 25778 77824
rect 25842 77760 25858 77824
rect 25922 77760 25938 77824
rect 26002 77760 26018 77824
rect 26082 77760 26090 77824
rect 25770 77759 26090 77760
rect 29269 77754 29335 77757
rect 31200 77754 32000 77784
rect 29269 77752 32000 77754
rect 29269 77696 29274 77752
rect 29330 77696 32000 77752
rect 29269 77694 32000 77696
rect 29269 77691 29335 77694
rect 31200 77664 32000 77694
rect 0 77618 800 77648
rect 1393 77618 1459 77621
rect 0 77616 1459 77618
rect 0 77560 1398 77616
rect 1454 77560 1459 77616
rect 0 77558 1459 77560
rect 0 77528 800 77558
rect 1393 77555 1459 77558
rect 28901 77346 28967 77349
rect 31200 77346 32000 77376
rect 28901 77344 32000 77346
rect 28901 77288 28906 77344
rect 28962 77288 32000 77344
rect 28901 77286 32000 77288
rect 28901 77283 28967 77286
rect 10874 77280 11194 77281
rect 10874 77216 10882 77280
rect 10946 77216 10962 77280
rect 11026 77216 11042 77280
rect 11106 77216 11122 77280
rect 11186 77216 11194 77280
rect 10874 77215 11194 77216
rect 20805 77280 21125 77281
rect 20805 77216 20813 77280
rect 20877 77216 20893 77280
rect 20957 77216 20973 77280
rect 21037 77216 21053 77280
rect 21117 77216 21125 77280
rect 31200 77256 32000 77286
rect 20805 77215 21125 77216
rect 0 76938 800 76968
rect 1393 76938 1459 76941
rect 0 76936 1459 76938
rect 0 76880 1398 76936
rect 1454 76880 1459 76936
rect 0 76878 1459 76880
rect 0 76848 800 76878
rect 1393 76875 1459 76878
rect 30097 76802 30163 76805
rect 31200 76802 32000 76832
rect 30097 76800 32000 76802
rect 30097 76744 30102 76800
rect 30158 76744 32000 76800
rect 30097 76742 32000 76744
rect 30097 76739 30163 76742
rect 5909 76736 6229 76737
rect 5909 76672 5917 76736
rect 5981 76672 5997 76736
rect 6061 76672 6077 76736
rect 6141 76672 6157 76736
rect 6221 76672 6229 76736
rect 5909 76671 6229 76672
rect 15840 76736 16160 76737
rect 15840 76672 15848 76736
rect 15912 76672 15928 76736
rect 15992 76672 16008 76736
rect 16072 76672 16088 76736
rect 16152 76672 16160 76736
rect 15840 76671 16160 76672
rect 25770 76736 26090 76737
rect 25770 76672 25778 76736
rect 25842 76672 25858 76736
rect 25922 76672 25938 76736
rect 26002 76672 26018 76736
rect 26082 76672 26090 76736
rect 31200 76712 32000 76742
rect 25770 76671 26090 76672
rect 30005 76394 30071 76397
rect 31200 76394 32000 76424
rect 30005 76392 32000 76394
rect 30005 76336 30010 76392
rect 30066 76336 32000 76392
rect 30005 76334 32000 76336
rect 30005 76331 30071 76334
rect 31200 76304 32000 76334
rect 0 76258 800 76288
rect 2865 76258 2931 76261
rect 0 76256 2931 76258
rect 0 76200 2870 76256
rect 2926 76200 2931 76256
rect 0 76198 2931 76200
rect 0 76168 800 76198
rect 2865 76195 2931 76198
rect 10874 76192 11194 76193
rect 10874 76128 10882 76192
rect 10946 76128 10962 76192
rect 11026 76128 11042 76192
rect 11106 76128 11122 76192
rect 11186 76128 11194 76192
rect 10874 76127 11194 76128
rect 20805 76192 21125 76193
rect 20805 76128 20813 76192
rect 20877 76128 20893 76192
rect 20957 76128 20973 76192
rect 21037 76128 21053 76192
rect 21117 76128 21125 76192
rect 20805 76127 21125 76128
rect 29269 75850 29335 75853
rect 31200 75850 32000 75880
rect 29269 75848 32000 75850
rect 29269 75792 29274 75848
rect 29330 75792 32000 75848
rect 29269 75790 32000 75792
rect 29269 75787 29335 75790
rect 31200 75760 32000 75790
rect 5909 75648 6229 75649
rect 0 75578 800 75608
rect 5909 75584 5917 75648
rect 5981 75584 5997 75648
rect 6061 75584 6077 75648
rect 6141 75584 6157 75648
rect 6221 75584 6229 75648
rect 5909 75583 6229 75584
rect 15840 75648 16160 75649
rect 15840 75584 15848 75648
rect 15912 75584 15928 75648
rect 15992 75584 16008 75648
rect 16072 75584 16088 75648
rect 16152 75584 16160 75648
rect 15840 75583 16160 75584
rect 25770 75648 26090 75649
rect 25770 75584 25778 75648
rect 25842 75584 25858 75648
rect 25922 75584 25938 75648
rect 26002 75584 26018 75648
rect 26082 75584 26090 75648
rect 25770 75583 26090 75584
rect 1577 75578 1643 75581
rect 0 75576 1643 75578
rect 0 75520 1582 75576
rect 1638 75520 1643 75576
rect 0 75518 1643 75520
rect 0 75488 800 75518
rect 1577 75515 1643 75518
rect 30189 75442 30255 75445
rect 31200 75442 32000 75472
rect 30189 75440 32000 75442
rect 30189 75384 30194 75440
rect 30250 75384 32000 75440
rect 30189 75382 32000 75384
rect 30189 75379 30255 75382
rect 31200 75352 32000 75382
rect 10874 75104 11194 75105
rect 0 75034 800 75064
rect 10874 75040 10882 75104
rect 10946 75040 10962 75104
rect 11026 75040 11042 75104
rect 11106 75040 11122 75104
rect 11186 75040 11194 75104
rect 10874 75039 11194 75040
rect 20805 75104 21125 75105
rect 20805 75040 20813 75104
rect 20877 75040 20893 75104
rect 20957 75040 20973 75104
rect 21037 75040 21053 75104
rect 21117 75040 21125 75104
rect 20805 75039 21125 75040
rect 1577 75034 1643 75037
rect 0 75032 1643 75034
rect 0 74976 1582 75032
rect 1638 74976 1643 75032
rect 0 74974 1643 74976
rect 0 74944 800 74974
rect 1577 74971 1643 74974
rect 30005 74898 30071 74901
rect 31200 74898 32000 74928
rect 30005 74896 32000 74898
rect 30005 74840 30010 74896
rect 30066 74840 32000 74896
rect 30005 74838 32000 74840
rect 30005 74835 30071 74838
rect 31200 74808 32000 74838
rect 5909 74560 6229 74561
rect 5909 74496 5917 74560
rect 5981 74496 5997 74560
rect 6061 74496 6077 74560
rect 6141 74496 6157 74560
rect 6221 74496 6229 74560
rect 5909 74495 6229 74496
rect 15840 74560 16160 74561
rect 15840 74496 15848 74560
rect 15912 74496 15928 74560
rect 15992 74496 16008 74560
rect 16072 74496 16088 74560
rect 16152 74496 16160 74560
rect 15840 74495 16160 74496
rect 25770 74560 26090 74561
rect 25770 74496 25778 74560
rect 25842 74496 25858 74560
rect 25922 74496 25938 74560
rect 26002 74496 26018 74560
rect 26082 74496 26090 74560
rect 25770 74495 26090 74496
rect 30189 74490 30255 74493
rect 31200 74490 32000 74520
rect 30189 74488 32000 74490
rect 30189 74432 30194 74488
rect 30250 74432 32000 74488
rect 30189 74430 32000 74432
rect 30189 74427 30255 74430
rect 31200 74400 32000 74430
rect 0 74354 800 74384
rect 1577 74354 1643 74357
rect 0 74352 1643 74354
rect 0 74296 1582 74352
rect 1638 74296 1643 74352
rect 0 74294 1643 74296
rect 0 74264 800 74294
rect 1577 74291 1643 74294
rect 30005 74082 30071 74085
rect 31200 74082 32000 74112
rect 30005 74080 32000 74082
rect 30005 74024 30010 74080
rect 30066 74024 32000 74080
rect 30005 74022 32000 74024
rect 30005 74019 30071 74022
rect 10874 74016 11194 74017
rect 10874 73952 10882 74016
rect 10946 73952 10962 74016
rect 11026 73952 11042 74016
rect 11106 73952 11122 74016
rect 11186 73952 11194 74016
rect 10874 73951 11194 73952
rect 20805 74016 21125 74017
rect 20805 73952 20813 74016
rect 20877 73952 20893 74016
rect 20957 73952 20973 74016
rect 21037 73952 21053 74016
rect 21117 73952 21125 74016
rect 31200 73992 32000 74022
rect 20805 73951 21125 73952
rect 0 73674 800 73704
rect 1577 73674 1643 73677
rect 0 73672 1643 73674
rect 0 73616 1582 73672
rect 1638 73616 1643 73672
rect 0 73614 1643 73616
rect 0 73584 800 73614
rect 1577 73611 1643 73614
rect 30189 73538 30255 73541
rect 31200 73538 32000 73568
rect 30189 73536 32000 73538
rect 30189 73480 30194 73536
rect 30250 73480 32000 73536
rect 30189 73478 32000 73480
rect 30189 73475 30255 73478
rect 5909 73472 6229 73473
rect 5909 73408 5917 73472
rect 5981 73408 5997 73472
rect 6061 73408 6077 73472
rect 6141 73408 6157 73472
rect 6221 73408 6229 73472
rect 5909 73407 6229 73408
rect 15840 73472 16160 73473
rect 15840 73408 15848 73472
rect 15912 73408 15928 73472
rect 15992 73408 16008 73472
rect 16072 73408 16088 73472
rect 16152 73408 16160 73472
rect 15840 73407 16160 73408
rect 25770 73472 26090 73473
rect 25770 73408 25778 73472
rect 25842 73408 25858 73472
rect 25922 73408 25938 73472
rect 26002 73408 26018 73472
rect 26082 73408 26090 73472
rect 31200 73448 32000 73478
rect 25770 73407 26090 73408
rect 15837 73130 15903 73133
rect 17401 73130 17467 73133
rect 15837 73128 17467 73130
rect 15837 73072 15842 73128
rect 15898 73072 17406 73128
rect 17462 73072 17467 73128
rect 15837 73070 17467 73072
rect 15837 73067 15903 73070
rect 17401 73067 17467 73070
rect 30005 73130 30071 73133
rect 31200 73130 32000 73160
rect 30005 73128 32000 73130
rect 30005 73072 30010 73128
rect 30066 73072 32000 73128
rect 30005 73070 32000 73072
rect 30005 73067 30071 73070
rect 31200 73040 32000 73070
rect 0 72994 800 73024
rect 1577 72994 1643 72997
rect 0 72992 1643 72994
rect 0 72936 1582 72992
rect 1638 72936 1643 72992
rect 0 72934 1643 72936
rect 0 72904 800 72934
rect 1577 72931 1643 72934
rect 10874 72928 11194 72929
rect 10874 72864 10882 72928
rect 10946 72864 10962 72928
rect 11026 72864 11042 72928
rect 11106 72864 11122 72928
rect 11186 72864 11194 72928
rect 10874 72863 11194 72864
rect 20805 72928 21125 72929
rect 20805 72864 20813 72928
rect 20877 72864 20893 72928
rect 20957 72864 20973 72928
rect 21037 72864 21053 72928
rect 21117 72864 21125 72928
rect 20805 72863 21125 72864
rect 30005 72586 30071 72589
rect 31200 72586 32000 72616
rect 30005 72584 32000 72586
rect 30005 72528 30010 72584
rect 30066 72528 32000 72584
rect 30005 72526 32000 72528
rect 30005 72523 30071 72526
rect 31200 72496 32000 72526
rect 5909 72384 6229 72385
rect 0 72314 800 72344
rect 5909 72320 5917 72384
rect 5981 72320 5997 72384
rect 6061 72320 6077 72384
rect 6141 72320 6157 72384
rect 6221 72320 6229 72384
rect 5909 72319 6229 72320
rect 15840 72384 16160 72385
rect 15840 72320 15848 72384
rect 15912 72320 15928 72384
rect 15992 72320 16008 72384
rect 16072 72320 16088 72384
rect 16152 72320 16160 72384
rect 15840 72319 16160 72320
rect 25770 72384 26090 72385
rect 25770 72320 25778 72384
rect 25842 72320 25858 72384
rect 25922 72320 25938 72384
rect 26002 72320 26018 72384
rect 26082 72320 26090 72384
rect 25770 72319 26090 72320
rect 1577 72314 1643 72317
rect 0 72312 1643 72314
rect 0 72256 1582 72312
rect 1638 72256 1643 72312
rect 0 72254 1643 72256
rect 0 72224 800 72254
rect 1577 72251 1643 72254
rect 30005 72178 30071 72181
rect 31200 72178 32000 72208
rect 30005 72176 32000 72178
rect 30005 72120 30010 72176
rect 30066 72120 32000 72176
rect 30005 72118 32000 72120
rect 30005 72115 30071 72118
rect 31200 72088 32000 72118
rect 10874 71840 11194 71841
rect 10874 71776 10882 71840
rect 10946 71776 10962 71840
rect 11026 71776 11042 71840
rect 11106 71776 11122 71840
rect 11186 71776 11194 71840
rect 10874 71775 11194 71776
rect 20805 71840 21125 71841
rect 20805 71776 20813 71840
rect 20877 71776 20893 71840
rect 20957 71776 20973 71840
rect 21037 71776 21053 71840
rect 21117 71776 21125 71840
rect 20805 71775 21125 71776
rect 0 71634 800 71664
rect 1577 71634 1643 71637
rect 0 71632 1643 71634
rect 0 71576 1582 71632
rect 1638 71576 1643 71632
rect 0 71574 1643 71576
rect 0 71544 800 71574
rect 1577 71571 1643 71574
rect 30005 71634 30071 71637
rect 31200 71634 32000 71664
rect 30005 71632 32000 71634
rect 30005 71576 30010 71632
rect 30066 71576 32000 71632
rect 30005 71574 32000 71576
rect 30005 71571 30071 71574
rect 31200 71544 32000 71574
rect 17493 71498 17559 71501
rect 18413 71498 18479 71501
rect 17493 71496 18479 71498
rect 17493 71440 17498 71496
rect 17554 71440 18418 71496
rect 18474 71440 18479 71496
rect 17493 71438 18479 71440
rect 17493 71435 17559 71438
rect 18413 71435 18479 71438
rect 5909 71296 6229 71297
rect 5909 71232 5917 71296
rect 5981 71232 5997 71296
rect 6061 71232 6077 71296
rect 6141 71232 6157 71296
rect 6221 71232 6229 71296
rect 5909 71231 6229 71232
rect 15840 71296 16160 71297
rect 15840 71232 15848 71296
rect 15912 71232 15928 71296
rect 15992 71232 16008 71296
rect 16072 71232 16088 71296
rect 16152 71232 16160 71296
rect 15840 71231 16160 71232
rect 25770 71296 26090 71297
rect 25770 71232 25778 71296
rect 25842 71232 25858 71296
rect 25922 71232 25938 71296
rect 26002 71232 26018 71296
rect 26082 71232 26090 71296
rect 25770 71231 26090 71232
rect 30005 71226 30071 71229
rect 31200 71226 32000 71256
rect 30005 71224 32000 71226
rect 30005 71168 30010 71224
rect 30066 71168 32000 71224
rect 30005 71166 32000 71168
rect 30005 71163 30071 71166
rect 31200 71136 32000 71166
rect 0 70954 800 70984
rect 1393 70954 1459 70957
rect 0 70952 1459 70954
rect 0 70896 1398 70952
rect 1454 70896 1459 70952
rect 0 70894 1459 70896
rect 0 70864 800 70894
rect 1393 70891 1459 70894
rect 10874 70752 11194 70753
rect 10874 70688 10882 70752
rect 10946 70688 10962 70752
rect 11026 70688 11042 70752
rect 11106 70688 11122 70752
rect 11186 70688 11194 70752
rect 10874 70687 11194 70688
rect 20805 70752 21125 70753
rect 20805 70688 20813 70752
rect 20877 70688 20893 70752
rect 20957 70688 20973 70752
rect 21037 70688 21053 70752
rect 21117 70688 21125 70752
rect 20805 70687 21125 70688
rect 30005 70682 30071 70685
rect 31200 70682 32000 70712
rect 30005 70680 32000 70682
rect 30005 70624 30010 70680
rect 30066 70624 32000 70680
rect 30005 70622 32000 70624
rect 30005 70619 30071 70622
rect 31200 70592 32000 70622
rect 0 70410 800 70440
rect 1577 70410 1643 70413
rect 0 70408 1643 70410
rect 0 70352 1582 70408
rect 1638 70352 1643 70408
rect 0 70350 1643 70352
rect 0 70320 800 70350
rect 1577 70347 1643 70350
rect 30005 70274 30071 70277
rect 31200 70274 32000 70304
rect 30005 70272 32000 70274
rect 30005 70216 30010 70272
rect 30066 70216 32000 70272
rect 30005 70214 32000 70216
rect 30005 70211 30071 70214
rect 5909 70208 6229 70209
rect 5909 70144 5917 70208
rect 5981 70144 5997 70208
rect 6061 70144 6077 70208
rect 6141 70144 6157 70208
rect 6221 70144 6229 70208
rect 5909 70143 6229 70144
rect 15840 70208 16160 70209
rect 15840 70144 15848 70208
rect 15912 70144 15928 70208
rect 15992 70144 16008 70208
rect 16072 70144 16088 70208
rect 16152 70144 16160 70208
rect 15840 70143 16160 70144
rect 25770 70208 26090 70209
rect 25770 70144 25778 70208
rect 25842 70144 25858 70208
rect 25922 70144 25938 70208
rect 26002 70144 26018 70208
rect 26082 70144 26090 70208
rect 31200 70184 32000 70214
rect 25770 70143 26090 70144
rect 29177 70004 29243 70005
rect 29126 70002 29132 70004
rect 29086 69942 29132 70002
rect 29196 70000 29243 70004
rect 29238 69944 29243 70000
rect 29126 69940 29132 69942
rect 29196 69940 29243 69944
rect 29177 69939 29243 69940
rect 0 69730 800 69760
rect 1577 69730 1643 69733
rect 0 69728 1643 69730
rect 0 69672 1582 69728
rect 1638 69672 1643 69728
rect 0 69670 1643 69672
rect 0 69640 800 69670
rect 1577 69667 1643 69670
rect 30005 69730 30071 69733
rect 31200 69730 32000 69760
rect 30005 69728 32000 69730
rect 30005 69672 30010 69728
rect 30066 69672 32000 69728
rect 30005 69670 32000 69672
rect 30005 69667 30071 69670
rect 10874 69664 11194 69665
rect 10874 69600 10882 69664
rect 10946 69600 10962 69664
rect 11026 69600 11042 69664
rect 11106 69600 11122 69664
rect 11186 69600 11194 69664
rect 10874 69599 11194 69600
rect 20805 69664 21125 69665
rect 20805 69600 20813 69664
rect 20877 69600 20893 69664
rect 20957 69600 20973 69664
rect 21037 69600 21053 69664
rect 21117 69600 21125 69664
rect 31200 69640 32000 69670
rect 20805 69599 21125 69600
rect 29269 69322 29335 69325
rect 31200 69322 32000 69352
rect 29269 69320 32000 69322
rect 29269 69264 29274 69320
rect 29330 69264 32000 69320
rect 29269 69262 32000 69264
rect 29269 69259 29335 69262
rect 31200 69232 32000 69262
rect 5909 69120 6229 69121
rect 0 69050 800 69080
rect 5909 69056 5917 69120
rect 5981 69056 5997 69120
rect 6061 69056 6077 69120
rect 6141 69056 6157 69120
rect 6221 69056 6229 69120
rect 5909 69055 6229 69056
rect 15840 69120 16160 69121
rect 15840 69056 15848 69120
rect 15912 69056 15928 69120
rect 15992 69056 16008 69120
rect 16072 69056 16088 69120
rect 16152 69056 16160 69120
rect 15840 69055 16160 69056
rect 25770 69120 26090 69121
rect 25770 69056 25778 69120
rect 25842 69056 25858 69120
rect 25922 69056 25938 69120
rect 26002 69056 26018 69120
rect 26082 69056 26090 69120
rect 25770 69055 26090 69056
rect 1577 69050 1643 69053
rect 0 69048 1643 69050
rect 0 68992 1582 69048
rect 1638 68992 1643 69048
rect 0 68990 1643 68992
rect 0 68960 800 68990
rect 1577 68987 1643 68990
rect 20437 68914 20503 68917
rect 20437 68912 20546 68914
rect 20437 68856 20442 68912
rect 20498 68856 20546 68912
rect 20437 68851 20546 68856
rect 10874 68576 11194 68577
rect 10874 68512 10882 68576
rect 10946 68512 10962 68576
rect 11026 68512 11042 68576
rect 11106 68512 11122 68576
rect 11186 68512 11194 68576
rect 10874 68511 11194 68512
rect 0 68370 800 68400
rect 20486 68373 20546 68851
rect 28901 68778 28967 68781
rect 31200 68778 32000 68808
rect 28901 68776 32000 68778
rect 28901 68720 28906 68776
rect 28962 68720 32000 68776
rect 28901 68718 32000 68720
rect 28901 68715 28967 68718
rect 31200 68688 32000 68718
rect 20805 68576 21125 68577
rect 20805 68512 20813 68576
rect 20877 68512 20893 68576
rect 20957 68512 20973 68576
rect 21037 68512 21053 68576
rect 21117 68512 21125 68576
rect 20805 68511 21125 68512
rect 1577 68370 1643 68373
rect 0 68368 1643 68370
rect 0 68312 1582 68368
rect 1638 68312 1643 68368
rect 0 68310 1643 68312
rect 0 68280 800 68310
rect 1577 68307 1643 68310
rect 20437 68368 20546 68373
rect 20437 68312 20442 68368
rect 20498 68312 20546 68368
rect 20437 68310 20546 68312
rect 29913 68370 29979 68373
rect 31200 68370 32000 68400
rect 29913 68368 32000 68370
rect 29913 68312 29918 68368
rect 29974 68312 32000 68368
rect 29913 68310 32000 68312
rect 20437 68307 20503 68310
rect 29913 68307 29979 68310
rect 31200 68280 32000 68310
rect 25037 68234 25103 68237
rect 27521 68234 27587 68237
rect 25037 68232 27587 68234
rect 25037 68176 25042 68232
rect 25098 68176 27526 68232
rect 27582 68176 27587 68232
rect 25037 68174 27587 68176
rect 25037 68171 25103 68174
rect 27521 68171 27587 68174
rect 5909 68032 6229 68033
rect 5909 67968 5917 68032
rect 5981 67968 5997 68032
rect 6061 67968 6077 68032
rect 6141 67968 6157 68032
rect 6221 67968 6229 68032
rect 5909 67967 6229 67968
rect 15840 68032 16160 68033
rect 15840 67968 15848 68032
rect 15912 67968 15928 68032
rect 15992 67968 16008 68032
rect 16072 67968 16088 68032
rect 16152 67968 16160 68032
rect 15840 67967 16160 67968
rect 25770 68032 26090 68033
rect 25770 67968 25778 68032
rect 25842 67968 25858 68032
rect 25922 67968 25938 68032
rect 26002 67968 26018 68032
rect 26082 67968 26090 68032
rect 25770 67967 26090 67968
rect 30005 67962 30071 67965
rect 31200 67962 32000 67992
rect 30005 67960 32000 67962
rect 30005 67904 30010 67960
rect 30066 67904 32000 67960
rect 30005 67902 32000 67904
rect 30005 67899 30071 67902
rect 31200 67872 32000 67902
rect 26049 67826 26115 67829
rect 27521 67826 27587 67829
rect 26049 67824 27587 67826
rect 26049 67768 26054 67824
rect 26110 67768 27526 67824
rect 27582 67768 27587 67824
rect 26049 67766 27587 67768
rect 26049 67763 26115 67766
rect 27521 67763 27587 67766
rect 0 67690 800 67720
rect 1577 67690 1643 67693
rect 0 67688 1643 67690
rect 0 67632 1582 67688
rect 1638 67632 1643 67688
rect 0 67630 1643 67632
rect 0 67600 800 67630
rect 1577 67627 1643 67630
rect 25681 67690 25747 67693
rect 27797 67690 27863 67693
rect 25681 67688 27863 67690
rect 25681 67632 25686 67688
rect 25742 67632 27802 67688
rect 27858 67632 27863 67688
rect 25681 67630 27863 67632
rect 25681 67627 25747 67630
rect 27797 67627 27863 67630
rect 27102 67492 27108 67556
rect 27172 67554 27178 67556
rect 27797 67554 27863 67557
rect 27172 67552 27863 67554
rect 27172 67496 27802 67552
rect 27858 67496 27863 67552
rect 27172 67494 27863 67496
rect 27172 67492 27178 67494
rect 27797 67491 27863 67494
rect 10874 67488 11194 67489
rect 10874 67424 10882 67488
rect 10946 67424 10962 67488
rect 11026 67424 11042 67488
rect 11106 67424 11122 67488
rect 11186 67424 11194 67488
rect 10874 67423 11194 67424
rect 20805 67488 21125 67489
rect 20805 67424 20813 67488
rect 20877 67424 20893 67488
rect 20957 67424 20973 67488
rect 21037 67424 21053 67488
rect 21117 67424 21125 67488
rect 20805 67423 21125 67424
rect 28901 67418 28967 67421
rect 31200 67418 32000 67448
rect 28901 67416 32000 67418
rect 28901 67360 28906 67416
rect 28962 67360 32000 67416
rect 28901 67358 32000 67360
rect 28901 67355 28967 67358
rect 31200 67328 32000 67358
rect 27245 67282 27311 67285
rect 26374 67280 27311 67282
rect 26374 67224 27250 67280
rect 27306 67224 27311 67280
rect 26374 67222 27311 67224
rect 26233 67146 26299 67149
rect 26374 67146 26434 67222
rect 27245 67219 27311 67222
rect 26233 67144 26434 67146
rect 26233 67088 26238 67144
rect 26294 67088 26434 67144
rect 26233 67086 26434 67088
rect 26233 67083 26299 67086
rect 0 67010 800 67040
rect 1577 67010 1643 67013
rect 0 67008 1643 67010
rect 0 66952 1582 67008
rect 1638 66952 1643 67008
rect 0 66950 1643 66952
rect 0 66920 800 66950
rect 1577 66947 1643 66950
rect 29913 67010 29979 67013
rect 31200 67010 32000 67040
rect 29913 67008 32000 67010
rect 29913 66952 29918 67008
rect 29974 66952 32000 67008
rect 29913 66950 32000 66952
rect 29913 66947 29979 66950
rect 5909 66944 6229 66945
rect 5909 66880 5917 66944
rect 5981 66880 5997 66944
rect 6061 66880 6077 66944
rect 6141 66880 6157 66944
rect 6221 66880 6229 66944
rect 5909 66879 6229 66880
rect 15840 66944 16160 66945
rect 15840 66880 15848 66944
rect 15912 66880 15928 66944
rect 15992 66880 16008 66944
rect 16072 66880 16088 66944
rect 16152 66880 16160 66944
rect 15840 66879 16160 66880
rect 25770 66944 26090 66945
rect 25770 66880 25778 66944
rect 25842 66880 25858 66944
rect 25922 66880 25938 66944
rect 26002 66880 26018 66944
rect 26082 66880 26090 66944
rect 31200 66920 32000 66950
rect 25770 66879 26090 66880
rect 26366 66812 26372 66876
rect 26436 66874 26442 66876
rect 26877 66874 26943 66877
rect 26436 66872 26943 66874
rect 26436 66816 26882 66872
rect 26938 66816 26943 66872
rect 26436 66814 26943 66816
rect 26436 66812 26442 66814
rect 26877 66811 26943 66814
rect 28901 66466 28967 66469
rect 31200 66466 32000 66496
rect 28901 66464 32000 66466
rect 28901 66408 28906 66464
rect 28962 66408 32000 66464
rect 28901 66406 32000 66408
rect 28901 66403 28967 66406
rect 10874 66400 11194 66401
rect 0 66330 800 66360
rect 10874 66336 10882 66400
rect 10946 66336 10962 66400
rect 11026 66336 11042 66400
rect 11106 66336 11122 66400
rect 11186 66336 11194 66400
rect 10874 66335 11194 66336
rect 20805 66400 21125 66401
rect 20805 66336 20813 66400
rect 20877 66336 20893 66400
rect 20957 66336 20973 66400
rect 21037 66336 21053 66400
rect 21117 66336 21125 66400
rect 31200 66376 32000 66406
rect 20805 66335 21125 66336
rect 1577 66330 1643 66333
rect 0 66328 1643 66330
rect 0 66272 1582 66328
rect 1638 66272 1643 66328
rect 0 66270 1643 66272
rect 0 66240 800 66270
rect 1577 66267 1643 66270
rect 18505 66194 18571 66197
rect 22553 66194 22619 66197
rect 18505 66192 22619 66194
rect 18505 66136 18510 66192
rect 18566 66136 22558 66192
rect 22614 66136 22619 66192
rect 18505 66134 22619 66136
rect 18505 66131 18571 66134
rect 22553 66131 22619 66134
rect 22645 66058 22711 66061
rect 25078 66058 25084 66060
rect 22645 66056 25084 66058
rect 22645 66000 22650 66056
rect 22706 66000 25084 66056
rect 22645 65998 25084 66000
rect 22645 65995 22711 65998
rect 25078 65996 25084 65998
rect 25148 66058 25154 66060
rect 25405 66058 25471 66061
rect 25148 66056 25471 66058
rect 25148 66000 25410 66056
rect 25466 66000 25471 66056
rect 25148 65998 25471 66000
rect 25148 65996 25154 65998
rect 25405 65995 25471 65998
rect 30005 66058 30071 66061
rect 31200 66058 32000 66088
rect 30005 66056 32000 66058
rect 30005 66000 30010 66056
rect 30066 66000 32000 66056
rect 30005 65998 32000 66000
rect 30005 65995 30071 65998
rect 31200 65968 32000 65998
rect 5909 65856 6229 65857
rect 0 65786 800 65816
rect 5909 65792 5917 65856
rect 5981 65792 5997 65856
rect 6061 65792 6077 65856
rect 6141 65792 6157 65856
rect 6221 65792 6229 65856
rect 5909 65791 6229 65792
rect 15840 65856 16160 65857
rect 15840 65792 15848 65856
rect 15912 65792 15928 65856
rect 15992 65792 16008 65856
rect 16072 65792 16088 65856
rect 16152 65792 16160 65856
rect 15840 65791 16160 65792
rect 25770 65856 26090 65857
rect 25770 65792 25778 65856
rect 25842 65792 25858 65856
rect 25922 65792 25938 65856
rect 26002 65792 26018 65856
rect 26082 65792 26090 65856
rect 25770 65791 26090 65792
rect 1577 65786 1643 65789
rect 0 65784 1643 65786
rect 0 65728 1582 65784
rect 1638 65728 1643 65784
rect 0 65726 1643 65728
rect 0 65696 800 65726
rect 1577 65723 1643 65726
rect 27654 65588 27660 65652
rect 27724 65650 27730 65652
rect 27889 65650 27955 65653
rect 28441 65652 28507 65653
rect 28390 65650 28396 65652
rect 27724 65648 27955 65650
rect 27724 65592 27894 65648
rect 27950 65592 27955 65648
rect 27724 65590 27955 65592
rect 28350 65590 28396 65650
rect 28460 65648 28507 65652
rect 28502 65592 28507 65648
rect 27724 65588 27730 65590
rect 27889 65587 27955 65590
rect 28390 65588 28396 65590
rect 28460 65588 28507 65592
rect 28441 65587 28507 65588
rect 28073 65514 28139 65517
rect 31200 65514 32000 65544
rect 28073 65512 32000 65514
rect 28073 65456 28078 65512
rect 28134 65456 32000 65512
rect 28073 65454 32000 65456
rect 28073 65451 28139 65454
rect 31200 65424 32000 65454
rect 10874 65312 11194 65313
rect 10874 65248 10882 65312
rect 10946 65248 10962 65312
rect 11026 65248 11042 65312
rect 11106 65248 11122 65312
rect 11186 65248 11194 65312
rect 10874 65247 11194 65248
rect 20805 65312 21125 65313
rect 20805 65248 20813 65312
rect 20877 65248 20893 65312
rect 20957 65248 20973 65312
rect 21037 65248 21053 65312
rect 21117 65248 21125 65312
rect 20805 65247 21125 65248
rect 0 65106 800 65136
rect 1577 65106 1643 65109
rect 0 65104 1643 65106
rect 0 65048 1582 65104
rect 1638 65048 1643 65104
rect 0 65046 1643 65048
rect 0 65016 800 65046
rect 1577 65043 1643 65046
rect 29821 65106 29887 65109
rect 31200 65106 32000 65136
rect 29821 65104 32000 65106
rect 29821 65048 29826 65104
rect 29882 65048 32000 65104
rect 29821 65046 32000 65048
rect 29821 65043 29887 65046
rect 31200 65016 32000 65046
rect 28073 64970 28139 64973
rect 28758 64970 28764 64972
rect 28073 64968 28764 64970
rect 28073 64912 28078 64968
rect 28134 64912 28764 64968
rect 28073 64910 28764 64912
rect 28073 64907 28139 64910
rect 28758 64908 28764 64910
rect 28828 64908 28834 64972
rect 5909 64768 6229 64769
rect 5909 64704 5917 64768
rect 5981 64704 5997 64768
rect 6061 64704 6077 64768
rect 6141 64704 6157 64768
rect 6221 64704 6229 64768
rect 5909 64703 6229 64704
rect 15840 64768 16160 64769
rect 15840 64704 15848 64768
rect 15912 64704 15928 64768
rect 15992 64704 16008 64768
rect 16072 64704 16088 64768
rect 16152 64704 16160 64768
rect 15840 64703 16160 64704
rect 25770 64768 26090 64769
rect 25770 64704 25778 64768
rect 25842 64704 25858 64768
rect 25922 64704 25938 64768
rect 26002 64704 26018 64768
rect 26082 64704 26090 64768
rect 25770 64703 26090 64704
rect 28625 64562 28691 64565
rect 31200 64562 32000 64592
rect 28625 64560 32000 64562
rect 28625 64504 28630 64560
rect 28686 64504 32000 64560
rect 28625 64502 32000 64504
rect 28625 64499 28691 64502
rect 31200 64472 32000 64502
rect 0 64426 800 64456
rect 1577 64426 1643 64429
rect 0 64424 1643 64426
rect 0 64368 1582 64424
rect 1638 64368 1643 64424
rect 0 64366 1643 64368
rect 0 64336 800 64366
rect 1577 64363 1643 64366
rect 26325 64426 26391 64429
rect 27889 64426 27955 64429
rect 26325 64424 27955 64426
rect 26325 64368 26330 64424
rect 26386 64368 27894 64424
rect 27950 64368 27955 64424
rect 26325 64366 27955 64368
rect 26325 64363 26391 64366
rect 27889 64363 27955 64366
rect 10874 64224 11194 64225
rect 10874 64160 10882 64224
rect 10946 64160 10962 64224
rect 11026 64160 11042 64224
rect 11106 64160 11122 64224
rect 11186 64160 11194 64224
rect 10874 64159 11194 64160
rect 20805 64224 21125 64225
rect 20805 64160 20813 64224
rect 20877 64160 20893 64224
rect 20957 64160 20973 64224
rect 21037 64160 21053 64224
rect 21117 64160 21125 64224
rect 20805 64159 21125 64160
rect 27838 64092 27844 64156
rect 27908 64154 27914 64156
rect 28165 64154 28231 64157
rect 27908 64152 28231 64154
rect 27908 64096 28170 64152
rect 28226 64096 28231 64152
rect 27908 64094 28231 64096
rect 27908 64092 27914 64094
rect 28165 64091 28231 64094
rect 28809 64154 28875 64157
rect 31200 64154 32000 64184
rect 28809 64152 32000 64154
rect 28809 64096 28814 64152
rect 28870 64096 32000 64152
rect 28809 64094 32000 64096
rect 28809 64091 28875 64094
rect 31200 64064 32000 64094
rect 28257 64020 28323 64021
rect 28206 64018 28212 64020
rect 28166 63958 28212 64018
rect 28276 64016 28323 64020
rect 28318 63960 28323 64016
rect 28206 63956 28212 63958
rect 28276 63956 28323 63960
rect 28257 63955 28323 63956
rect 28073 63882 28139 63885
rect 31385 63882 31451 63885
rect 28073 63880 31451 63882
rect 28073 63824 28078 63880
rect 28134 63824 31390 63880
rect 31446 63824 31451 63880
rect 28073 63822 31451 63824
rect 28073 63819 28139 63822
rect 31385 63819 31451 63822
rect 0 63746 800 63776
rect 1577 63746 1643 63749
rect 0 63744 1643 63746
rect 0 63688 1582 63744
rect 1638 63688 1643 63744
rect 0 63686 1643 63688
rect 0 63656 800 63686
rect 1577 63683 1643 63686
rect 26550 63684 26556 63748
rect 26620 63746 26626 63748
rect 27429 63746 27495 63749
rect 26620 63744 27495 63746
rect 26620 63688 27434 63744
rect 27490 63688 27495 63744
rect 26620 63686 27495 63688
rect 26620 63684 26626 63686
rect 27429 63683 27495 63686
rect 5909 63680 6229 63681
rect 5909 63616 5917 63680
rect 5981 63616 5997 63680
rect 6061 63616 6077 63680
rect 6141 63616 6157 63680
rect 6221 63616 6229 63680
rect 5909 63615 6229 63616
rect 15840 63680 16160 63681
rect 15840 63616 15848 63680
rect 15912 63616 15928 63680
rect 15992 63616 16008 63680
rect 16072 63616 16088 63680
rect 16152 63616 16160 63680
rect 15840 63615 16160 63616
rect 25770 63680 26090 63681
rect 25770 63616 25778 63680
rect 25842 63616 25858 63680
rect 25922 63616 25938 63680
rect 26002 63616 26018 63680
rect 26082 63616 26090 63680
rect 25770 63615 26090 63616
rect 29913 63610 29979 63613
rect 31200 63610 32000 63640
rect 29913 63608 32000 63610
rect 29913 63552 29918 63608
rect 29974 63552 32000 63608
rect 29913 63550 32000 63552
rect 29913 63547 29979 63550
rect 31200 63520 32000 63550
rect 28533 63474 28599 63477
rect 28942 63474 28948 63476
rect 28533 63472 28948 63474
rect 28533 63416 28538 63472
rect 28594 63416 28948 63472
rect 28533 63414 28948 63416
rect 28533 63411 28599 63414
rect 28942 63412 28948 63414
rect 29012 63412 29018 63476
rect 27613 63202 27679 63205
rect 31200 63202 32000 63232
rect 27613 63200 32000 63202
rect 27613 63144 27618 63200
rect 27674 63144 32000 63200
rect 27613 63142 32000 63144
rect 27613 63139 27679 63142
rect 10874 63136 11194 63137
rect 0 63066 800 63096
rect 10874 63072 10882 63136
rect 10946 63072 10962 63136
rect 11026 63072 11042 63136
rect 11106 63072 11122 63136
rect 11186 63072 11194 63136
rect 10874 63071 11194 63072
rect 20805 63136 21125 63137
rect 20805 63072 20813 63136
rect 20877 63072 20893 63136
rect 20957 63072 20973 63136
rect 21037 63072 21053 63136
rect 21117 63072 21125 63136
rect 31200 63112 32000 63142
rect 20805 63071 21125 63072
rect 1577 63066 1643 63069
rect 0 63064 1643 63066
rect 0 63008 1582 63064
rect 1638 63008 1643 63064
rect 0 63006 1643 63008
rect 0 62976 800 63006
rect 1577 63003 1643 63006
rect 26509 63066 26575 63069
rect 28349 63068 28415 63069
rect 28533 63068 28599 63069
rect 28349 63066 28396 63068
rect 26509 63064 28136 63066
rect 26509 63008 26514 63064
rect 26570 63008 28136 63064
rect 26509 63006 28136 63008
rect 28304 63064 28396 63066
rect 28304 63008 28354 63064
rect 28304 63006 28396 63008
rect 26509 63003 26575 63006
rect 27521 62932 27587 62933
rect 27470 62930 27476 62932
rect 27430 62870 27476 62930
rect 27540 62928 27587 62932
rect 27582 62872 27587 62928
rect 27470 62868 27476 62870
rect 27540 62868 27587 62872
rect 28076 62930 28136 63006
rect 28349 63004 28396 63006
rect 28460 63004 28466 63068
rect 28533 63064 28580 63068
rect 28644 63066 28650 63068
rect 28533 63008 28538 63064
rect 28533 63004 28580 63008
rect 28644 63006 28690 63066
rect 28644 63004 28650 63006
rect 28349 63003 28415 63004
rect 28533 63003 28599 63004
rect 28533 62930 28599 62933
rect 28076 62928 28599 62930
rect 28076 62872 28538 62928
rect 28594 62872 28599 62928
rect 28076 62870 28599 62872
rect 27521 62867 27587 62868
rect 28533 62867 28599 62870
rect 27705 62794 27771 62797
rect 31200 62794 32000 62824
rect 27705 62792 32000 62794
rect 27705 62736 27710 62792
rect 27766 62736 32000 62792
rect 27705 62734 32000 62736
rect 27705 62731 27771 62734
rect 31200 62704 32000 62734
rect 5909 62592 6229 62593
rect 5909 62528 5917 62592
rect 5981 62528 5997 62592
rect 6061 62528 6077 62592
rect 6141 62528 6157 62592
rect 6221 62528 6229 62592
rect 5909 62527 6229 62528
rect 15840 62592 16160 62593
rect 15840 62528 15848 62592
rect 15912 62528 15928 62592
rect 15992 62528 16008 62592
rect 16072 62528 16088 62592
rect 16152 62528 16160 62592
rect 15840 62527 16160 62528
rect 25770 62592 26090 62593
rect 25770 62528 25778 62592
rect 25842 62528 25858 62592
rect 25922 62528 25938 62592
rect 26002 62528 26018 62592
rect 26082 62528 26090 62592
rect 25770 62527 26090 62528
rect 0 62386 800 62416
rect 1577 62386 1643 62389
rect 0 62384 1643 62386
rect 0 62328 1582 62384
rect 1638 62328 1643 62384
rect 0 62326 1643 62328
rect 0 62296 800 62326
rect 1577 62323 1643 62326
rect 17309 62386 17375 62389
rect 24853 62386 24919 62389
rect 25221 62388 25287 62389
rect 25221 62386 25268 62388
rect 17309 62384 24919 62386
rect 17309 62328 17314 62384
rect 17370 62328 24858 62384
rect 24914 62328 24919 62384
rect 17309 62326 24919 62328
rect 25176 62384 25268 62386
rect 25176 62328 25226 62384
rect 25176 62326 25268 62328
rect 17309 62323 17375 62326
rect 24853 62323 24919 62326
rect 25221 62324 25268 62326
rect 25332 62324 25338 62388
rect 26182 62324 26188 62388
rect 26252 62386 26258 62388
rect 27245 62386 27311 62389
rect 26252 62384 27311 62386
rect 26252 62328 27250 62384
rect 27306 62328 27311 62384
rect 26252 62326 27311 62328
rect 26252 62324 26258 62326
rect 25221 62323 25287 62324
rect 27245 62323 27311 62326
rect 27613 62250 27679 62253
rect 31200 62250 32000 62280
rect 27613 62248 32000 62250
rect 27613 62192 27618 62248
rect 27674 62192 32000 62248
rect 27613 62190 32000 62192
rect 27613 62187 27679 62190
rect 31200 62160 32000 62190
rect 24761 62114 24827 62117
rect 27429 62114 27495 62117
rect 24761 62112 27495 62114
rect 24761 62056 24766 62112
rect 24822 62056 27434 62112
rect 27490 62056 27495 62112
rect 24761 62054 27495 62056
rect 24761 62051 24827 62054
rect 27429 62051 27495 62054
rect 27889 62114 27955 62117
rect 28390 62114 28396 62116
rect 27889 62112 28396 62114
rect 27889 62056 27894 62112
rect 27950 62056 28396 62112
rect 27889 62054 28396 62056
rect 27889 62051 27955 62054
rect 28390 62052 28396 62054
rect 28460 62052 28466 62116
rect 10874 62048 11194 62049
rect 10874 61984 10882 62048
rect 10946 61984 10962 62048
rect 11026 61984 11042 62048
rect 11106 61984 11122 62048
rect 11186 61984 11194 62048
rect 10874 61983 11194 61984
rect 20805 62048 21125 62049
rect 20805 61984 20813 62048
rect 20877 61984 20893 62048
rect 20957 61984 20973 62048
rect 21037 61984 21053 62048
rect 21117 61984 21125 62048
rect 20805 61983 21125 61984
rect 28625 61842 28691 61845
rect 31200 61842 32000 61872
rect 28625 61840 32000 61842
rect 28625 61784 28630 61840
rect 28686 61784 32000 61840
rect 28625 61782 32000 61784
rect 28625 61779 28691 61782
rect 31200 61752 32000 61782
rect 0 61706 800 61736
rect 1577 61706 1643 61709
rect 0 61704 1643 61706
rect 0 61648 1582 61704
rect 1638 61648 1643 61704
rect 0 61646 1643 61648
rect 0 61616 800 61646
rect 1577 61643 1643 61646
rect 24853 61706 24919 61709
rect 25037 61706 25103 61709
rect 28625 61708 28691 61709
rect 28574 61706 28580 61708
rect 24853 61704 25103 61706
rect 24853 61648 24858 61704
rect 24914 61648 25042 61704
rect 25098 61648 25103 61704
rect 24853 61646 25103 61648
rect 28534 61646 28580 61706
rect 28644 61704 28691 61708
rect 28686 61648 28691 61704
rect 24853 61643 24919 61646
rect 25037 61643 25103 61646
rect 28574 61644 28580 61646
rect 28644 61644 28691 61648
rect 28625 61643 28691 61644
rect 28717 61572 28783 61573
rect 28717 61570 28764 61572
rect 28672 61568 28764 61570
rect 28672 61512 28722 61568
rect 28672 61510 28764 61512
rect 28717 61508 28764 61510
rect 28828 61508 28834 61572
rect 28717 61507 28783 61508
rect 5909 61504 6229 61505
rect 5909 61440 5917 61504
rect 5981 61440 5997 61504
rect 6061 61440 6077 61504
rect 6141 61440 6157 61504
rect 6221 61440 6229 61504
rect 5909 61439 6229 61440
rect 15840 61504 16160 61505
rect 15840 61440 15848 61504
rect 15912 61440 15928 61504
rect 15992 61440 16008 61504
rect 16072 61440 16088 61504
rect 16152 61440 16160 61504
rect 15840 61439 16160 61440
rect 25770 61504 26090 61505
rect 25770 61440 25778 61504
rect 25842 61440 25858 61504
rect 25922 61440 25938 61504
rect 26002 61440 26018 61504
rect 26082 61440 26090 61504
rect 25770 61439 26090 61440
rect 26785 61434 26851 61437
rect 26918 61434 26924 61436
rect 26785 61432 26924 61434
rect 26785 61376 26790 61432
rect 26846 61376 26924 61432
rect 26785 61374 26924 61376
rect 26785 61371 26851 61374
rect 26918 61372 26924 61374
rect 26988 61372 26994 61436
rect 28809 61434 28875 61437
rect 29310 61434 29316 61436
rect 28809 61432 29316 61434
rect 28809 61376 28814 61432
rect 28870 61376 29316 61432
rect 28809 61374 29316 61376
rect 28809 61371 28875 61374
rect 29310 61372 29316 61374
rect 29380 61372 29386 61436
rect 26601 61298 26667 61301
rect 26734 61298 26740 61300
rect 26601 61296 26740 61298
rect 26601 61240 26606 61296
rect 26662 61240 26740 61296
rect 26601 61238 26740 61240
rect 26601 61235 26667 61238
rect 26734 61236 26740 61238
rect 26804 61236 26810 61300
rect 28441 61298 28507 61301
rect 28574 61298 28580 61300
rect 28441 61296 28580 61298
rect 28441 61240 28446 61296
rect 28502 61240 28580 61296
rect 28441 61238 28580 61240
rect 28441 61235 28507 61238
rect 28574 61236 28580 61238
rect 28644 61236 28650 61300
rect 28809 61298 28875 61301
rect 29126 61298 29132 61300
rect 28809 61296 29132 61298
rect 28809 61240 28814 61296
rect 28870 61240 29132 61296
rect 28809 61238 29132 61240
rect 28809 61235 28875 61238
rect 29126 61236 29132 61238
rect 29196 61236 29202 61300
rect 29729 61298 29795 61301
rect 31200 61298 32000 61328
rect 29729 61296 32000 61298
rect 29729 61240 29734 61296
rect 29790 61240 32000 61296
rect 29729 61238 32000 61240
rect 29729 61235 29795 61238
rect 31200 61208 32000 61238
rect 0 61162 800 61192
rect 1577 61162 1643 61165
rect 0 61160 1643 61162
rect 0 61104 1582 61160
rect 1638 61104 1643 61160
rect 0 61102 1643 61104
rect 0 61072 800 61102
rect 1577 61099 1643 61102
rect 18965 61162 19031 61165
rect 25773 61162 25839 61165
rect 18965 61160 25839 61162
rect 18965 61104 18970 61160
rect 19026 61104 25778 61160
rect 25834 61104 25839 61160
rect 18965 61102 25839 61104
rect 18965 61099 19031 61102
rect 25773 61099 25839 61102
rect 26233 61162 26299 61165
rect 27705 61162 27771 61165
rect 28206 61162 28212 61164
rect 26233 61160 26986 61162
rect 26233 61104 26238 61160
rect 26294 61104 26986 61160
rect 26233 61102 26986 61104
rect 26233 61099 26299 61102
rect 26926 61029 26986 61102
rect 27705 61160 28212 61162
rect 27705 61104 27710 61160
rect 27766 61104 28212 61160
rect 27705 61102 28212 61104
rect 27705 61099 27771 61102
rect 28206 61100 28212 61102
rect 28276 61100 28282 61164
rect 28809 61160 28875 61165
rect 28809 61104 28814 61160
rect 28870 61104 28875 61160
rect 28809 61099 28875 61104
rect 29085 61162 29151 61165
rect 29085 61160 29194 61162
rect 29085 61104 29090 61160
rect 29146 61104 29194 61160
rect 29085 61099 29194 61104
rect 29494 61100 29500 61164
rect 29564 61162 29570 61164
rect 29637 61162 29703 61165
rect 29564 61160 29703 61162
rect 29564 61104 29642 61160
rect 29698 61104 29703 61160
rect 29564 61102 29703 61104
rect 29564 61100 29570 61102
rect 29637 61099 29703 61102
rect 26417 61026 26483 61029
rect 26550 61026 26556 61028
rect 26417 61024 26556 61026
rect 26417 60968 26422 61024
rect 26478 60968 26556 61024
rect 26417 60966 26556 60968
rect 26417 60963 26483 60966
rect 26550 60964 26556 60966
rect 26620 60964 26626 61028
rect 26926 61024 27035 61029
rect 26926 60968 26974 61024
rect 27030 60968 27035 61024
rect 26926 60966 27035 60968
rect 26969 60963 27035 60966
rect 27153 61024 27219 61029
rect 27337 61026 27403 61029
rect 27153 60968 27158 61024
rect 27214 60968 27219 61024
rect 27153 60963 27219 60968
rect 27294 61024 27403 61026
rect 27294 60968 27342 61024
rect 27398 60968 27403 61024
rect 27294 60963 27403 60968
rect 27889 61026 27955 61029
rect 28073 61026 28139 61029
rect 27889 61024 28139 61026
rect 27889 60968 27894 61024
rect 27950 60968 28078 61024
rect 28134 60968 28139 61024
rect 27889 60966 28139 60968
rect 27889 60963 27955 60966
rect 28073 60963 28139 60966
rect 28206 60964 28212 61028
rect 28276 61026 28282 61028
rect 28533 61026 28599 61029
rect 28812 61026 28872 61099
rect 28276 61024 28599 61026
rect 28276 60968 28538 61024
rect 28594 60968 28599 61024
rect 28276 60966 28599 60968
rect 28276 60964 28282 60966
rect 28533 60963 28599 60966
rect 28766 60966 28872 61026
rect 29134 61026 29194 61099
rect 30005 61026 30071 61029
rect 29134 61024 30071 61026
rect 29134 60968 30010 61024
rect 30066 60968 30071 61024
rect 29134 60966 30071 60968
rect 10874 60960 11194 60961
rect 10874 60896 10882 60960
rect 10946 60896 10962 60960
rect 11026 60896 11042 60960
rect 11106 60896 11122 60960
rect 11186 60896 11194 60960
rect 10874 60895 11194 60896
rect 20805 60960 21125 60961
rect 20805 60896 20813 60960
rect 20877 60896 20893 60960
rect 20957 60896 20973 60960
rect 21037 60896 21053 60960
rect 21117 60896 21125 60960
rect 20805 60895 21125 60896
rect 25313 60892 25379 60893
rect 25262 60890 25268 60892
rect 25222 60830 25268 60890
rect 25332 60888 25379 60892
rect 25374 60832 25379 60888
rect 25262 60828 25268 60830
rect 25332 60828 25379 60832
rect 25313 60827 25379 60828
rect 25589 60890 25655 60893
rect 26366 60890 26372 60892
rect 25589 60888 26372 60890
rect 25589 60832 25594 60888
rect 25650 60832 26372 60888
rect 25589 60830 26372 60832
rect 25589 60827 25655 60830
rect 26366 60828 26372 60830
rect 26436 60828 26442 60892
rect 20805 60754 20871 60757
rect 22369 60754 22435 60757
rect 25865 60754 25931 60757
rect 20805 60752 22435 60754
rect 20805 60696 20810 60752
rect 20866 60696 22374 60752
rect 22430 60696 22435 60752
rect 20805 60694 22435 60696
rect 20805 60691 20871 60694
rect 22369 60691 22435 60694
rect 25224 60752 25931 60754
rect 25224 60696 25870 60752
rect 25926 60696 25931 60752
rect 25224 60694 25931 60696
rect 0 60482 800 60512
rect 1577 60482 1643 60485
rect 0 60480 1643 60482
rect 0 60424 1582 60480
rect 1638 60424 1643 60480
rect 0 60422 1643 60424
rect 0 60392 800 60422
rect 1577 60419 1643 60422
rect 24577 60482 24643 60485
rect 25037 60482 25103 60485
rect 24577 60480 25103 60482
rect 24577 60424 24582 60480
rect 24638 60424 25042 60480
rect 25098 60424 25103 60480
rect 24577 60422 25103 60424
rect 24577 60419 24643 60422
rect 25037 60419 25103 60422
rect 5909 60416 6229 60417
rect 5909 60352 5917 60416
rect 5981 60352 5997 60416
rect 6061 60352 6077 60416
rect 6141 60352 6157 60416
rect 6221 60352 6229 60416
rect 5909 60351 6229 60352
rect 15840 60416 16160 60417
rect 15840 60352 15848 60416
rect 15912 60352 15928 60416
rect 15992 60352 16008 60416
rect 16072 60352 16088 60416
rect 16152 60352 16160 60416
rect 15840 60351 16160 60352
rect 24577 60346 24643 60349
rect 25224 60346 25284 60694
rect 25865 60691 25931 60694
rect 25957 60618 26023 60621
rect 24577 60344 25284 60346
rect 24577 60288 24582 60344
rect 24638 60288 25284 60344
rect 24577 60286 25284 60288
rect 25638 60616 26023 60618
rect 25638 60560 25962 60616
rect 26018 60560 26023 60616
rect 25638 60558 26023 60560
rect 24577 60283 24643 60286
rect 19333 60210 19399 60213
rect 19885 60210 19951 60213
rect 19333 60208 19951 60210
rect 19333 60152 19338 60208
rect 19394 60152 19890 60208
rect 19946 60152 19951 60208
rect 19333 60150 19951 60152
rect 25638 60210 25698 60558
rect 25957 60555 26023 60558
rect 26969 60618 27035 60621
rect 27156 60618 27216 60963
rect 27294 60620 27354 60963
rect 28766 60890 28826 60966
rect 27432 60830 28826 60890
rect 26969 60616 27216 60618
rect 26969 60560 26974 60616
rect 27030 60560 27216 60616
rect 26969 60558 27216 60560
rect 26969 60555 27035 60558
rect 27286 60556 27292 60620
rect 27356 60556 27362 60620
rect 26734 60420 26740 60484
rect 26804 60482 26810 60484
rect 27432 60482 27492 60830
rect 29134 60757 29194 60966
rect 30005 60963 30071 60966
rect 29269 60890 29335 60893
rect 29821 60890 29887 60893
rect 31200 60890 32000 60920
rect 29269 60888 29378 60890
rect 29269 60832 29274 60888
rect 29330 60832 29378 60888
rect 29269 60827 29378 60832
rect 29821 60888 32000 60890
rect 29821 60832 29826 60888
rect 29882 60832 32000 60888
rect 29821 60830 32000 60832
rect 29821 60827 29887 60830
rect 29134 60752 29243 60757
rect 29134 60696 29182 60752
rect 29238 60696 29243 60752
rect 29134 60694 29243 60696
rect 29177 60691 29243 60694
rect 28809 60618 28875 60621
rect 26804 60422 27492 60482
rect 27892 60616 28875 60618
rect 27892 60560 28814 60616
rect 28870 60560 28875 60616
rect 27892 60558 28875 60560
rect 26804 60420 26810 60422
rect 25770 60416 26090 60417
rect 25770 60352 25778 60416
rect 25842 60352 25858 60416
rect 25922 60352 25938 60416
rect 26002 60352 26018 60416
rect 26082 60352 26090 60416
rect 25770 60351 26090 60352
rect 26918 60284 26924 60348
rect 26988 60346 26994 60348
rect 27061 60346 27127 60349
rect 26988 60344 27127 60346
rect 26988 60288 27066 60344
rect 27122 60288 27127 60344
rect 26988 60286 27127 60288
rect 27892 60346 27952 60558
rect 28809 60555 28875 60558
rect 29085 60618 29151 60621
rect 29318 60618 29378 60827
rect 31200 60800 32000 60830
rect 29085 60616 29378 60618
rect 29085 60560 29090 60616
rect 29146 60560 29378 60616
rect 29085 60558 29378 60560
rect 29085 60555 29151 60558
rect 29361 60484 29427 60485
rect 29310 60482 29316 60484
rect 29270 60422 29316 60482
rect 29380 60480 29427 60484
rect 29422 60424 29427 60480
rect 29310 60420 29316 60422
rect 29380 60420 29427 60424
rect 29361 60419 29427 60420
rect 28022 60346 28028 60348
rect 27892 60286 28028 60346
rect 26988 60284 26994 60286
rect 27061 60283 27127 60286
rect 28022 60284 28028 60286
rect 28092 60284 28098 60348
rect 28533 60346 28599 60349
rect 31200 60346 32000 60376
rect 28533 60344 32000 60346
rect 28533 60288 28538 60344
rect 28594 60288 32000 60344
rect 28533 60286 32000 60288
rect 28533 60283 28599 60286
rect 31200 60256 32000 60286
rect 25773 60210 25839 60213
rect 26141 60212 26207 60213
rect 26141 60210 26188 60212
rect 25638 60208 25839 60210
rect 25638 60152 25778 60208
rect 25834 60152 25839 60208
rect 25638 60150 25839 60152
rect 26096 60208 26188 60210
rect 26096 60152 26146 60208
rect 26096 60150 26188 60152
rect 19333 60147 19399 60150
rect 19885 60147 19951 60150
rect 25773 60147 25839 60150
rect 26141 60148 26188 60150
rect 26252 60148 26258 60212
rect 27153 60210 27219 60213
rect 27838 60210 27844 60212
rect 27153 60208 27844 60210
rect 27153 60152 27158 60208
rect 27214 60152 27844 60208
rect 27153 60150 27844 60152
rect 26141 60147 26207 60148
rect 27153 60147 27219 60150
rect 27838 60148 27844 60150
rect 27908 60210 27914 60212
rect 28073 60210 28139 60213
rect 27908 60208 28139 60210
rect 27908 60152 28078 60208
rect 28134 60152 28139 60208
rect 27908 60150 28139 60152
rect 27908 60148 27914 60150
rect 28073 60147 28139 60150
rect 28574 60148 28580 60212
rect 28644 60210 28650 60212
rect 29361 60210 29427 60213
rect 28644 60208 29427 60210
rect 28644 60152 29366 60208
rect 29422 60152 29427 60208
rect 28644 60150 29427 60152
rect 28644 60148 28650 60150
rect 29361 60147 29427 60150
rect 18965 60074 19031 60077
rect 24669 60074 24735 60077
rect 18965 60072 24735 60074
rect 18965 60016 18970 60072
rect 19026 60016 24674 60072
rect 24730 60016 24735 60072
rect 18965 60014 24735 60016
rect 18965 60011 19031 60014
rect 24669 60011 24735 60014
rect 26601 60072 26667 60077
rect 26601 60016 26606 60072
rect 26662 60016 26667 60072
rect 26601 60011 26667 60016
rect 26785 60074 26851 60077
rect 28206 60074 28212 60076
rect 26785 60072 28212 60074
rect 26785 60016 26790 60072
rect 26846 60016 28212 60072
rect 26785 60014 28212 60016
rect 26785 60011 26851 60014
rect 28206 60012 28212 60014
rect 28276 60012 28282 60076
rect 28809 60074 28875 60077
rect 28942 60074 28948 60076
rect 28809 60072 28948 60074
rect 28809 60016 28814 60072
rect 28870 60016 28948 60072
rect 28809 60014 28948 60016
rect 28809 60011 28875 60014
rect 28942 60012 28948 60014
rect 29012 60012 29018 60076
rect 25262 59876 25268 59940
rect 25332 59938 25338 59940
rect 25865 59938 25931 59941
rect 25332 59936 25931 59938
rect 25332 59880 25870 59936
rect 25926 59880 25931 59936
rect 25332 59878 25931 59880
rect 26604 59938 26664 60011
rect 31200 59938 32000 59968
rect 26604 59878 32000 59938
rect 25332 59876 25338 59878
rect 25865 59875 25931 59878
rect 10874 59872 11194 59873
rect 0 59802 800 59832
rect 10874 59808 10882 59872
rect 10946 59808 10962 59872
rect 11026 59808 11042 59872
rect 11106 59808 11122 59872
rect 11186 59808 11194 59872
rect 10874 59807 11194 59808
rect 20805 59872 21125 59873
rect 20805 59808 20813 59872
rect 20877 59808 20893 59872
rect 20957 59808 20973 59872
rect 21037 59808 21053 59872
rect 21117 59808 21125 59872
rect 31200 59848 32000 59878
rect 20805 59807 21125 59808
rect 1577 59802 1643 59805
rect 0 59800 1643 59802
rect 0 59744 1582 59800
rect 1638 59744 1643 59800
rect 0 59742 1643 59744
rect 0 59712 800 59742
rect 1577 59739 1643 59742
rect 27654 59740 27660 59804
rect 27724 59802 27730 59804
rect 29678 59802 29684 59804
rect 27724 59742 29684 59802
rect 27724 59740 27730 59742
rect 29678 59740 29684 59742
rect 29748 59802 29754 59804
rect 29821 59802 29887 59805
rect 29748 59800 29887 59802
rect 29748 59744 29826 59800
rect 29882 59744 29887 59800
rect 29748 59742 29887 59744
rect 29748 59740 29754 59742
rect 29821 59739 29887 59742
rect 25630 59604 25636 59668
rect 25700 59666 25706 59668
rect 25865 59666 25931 59669
rect 25700 59664 25931 59666
rect 25700 59608 25870 59664
rect 25926 59608 25931 59664
rect 25700 59606 25931 59608
rect 25700 59604 25706 59606
rect 25865 59603 25931 59606
rect 26049 59666 26115 59669
rect 28073 59666 28139 59669
rect 26049 59664 28139 59666
rect 26049 59608 26054 59664
rect 26110 59608 28078 59664
rect 28134 59608 28139 59664
rect 26049 59606 28139 59608
rect 26049 59603 26115 59606
rect 28073 59603 28139 59606
rect 26550 59468 26556 59532
rect 26620 59530 26626 59532
rect 26969 59530 27035 59533
rect 26620 59528 27035 59530
rect 26620 59472 26974 59528
rect 27030 59472 27035 59528
rect 26620 59470 27035 59472
rect 26620 59468 26626 59470
rect 26969 59467 27035 59470
rect 28073 59530 28139 59533
rect 28390 59530 28396 59532
rect 28073 59528 28396 59530
rect 28073 59472 28078 59528
rect 28134 59472 28396 59528
rect 28073 59470 28396 59472
rect 28073 59467 28139 59470
rect 28390 59468 28396 59470
rect 28460 59468 28466 59532
rect 28901 59394 28967 59397
rect 31200 59394 32000 59424
rect 28901 59392 32000 59394
rect 28901 59336 28906 59392
rect 28962 59336 32000 59392
rect 28901 59334 32000 59336
rect 28901 59331 28967 59334
rect 5909 59328 6229 59329
rect 5909 59264 5917 59328
rect 5981 59264 5997 59328
rect 6061 59264 6077 59328
rect 6141 59264 6157 59328
rect 6221 59264 6229 59328
rect 5909 59263 6229 59264
rect 15840 59328 16160 59329
rect 15840 59264 15848 59328
rect 15912 59264 15928 59328
rect 15992 59264 16008 59328
rect 16072 59264 16088 59328
rect 16152 59264 16160 59328
rect 15840 59263 16160 59264
rect 25770 59328 26090 59329
rect 25770 59264 25778 59328
rect 25842 59264 25858 59328
rect 25922 59264 25938 59328
rect 26002 59264 26018 59328
rect 26082 59264 26090 59328
rect 31200 59304 32000 59334
rect 25770 59263 26090 59264
rect 27102 59196 27108 59260
rect 27172 59258 27178 59260
rect 28625 59258 28691 59261
rect 27172 59256 28691 59258
rect 27172 59200 28630 59256
rect 28686 59200 28691 59256
rect 27172 59198 28691 59200
rect 27172 59196 27178 59198
rect 0 59122 800 59152
rect 1577 59122 1643 59125
rect 0 59120 1643 59122
rect 0 59064 1582 59120
rect 1638 59064 1643 59120
rect 0 59062 1643 59064
rect 0 59032 800 59062
rect 1577 59059 1643 59062
rect 24117 59122 24183 59125
rect 27110 59122 27170 59196
rect 28625 59195 28691 59198
rect 24117 59120 27170 59122
rect 24117 59064 24122 59120
rect 24178 59064 27170 59120
rect 24117 59062 27170 59064
rect 24117 59059 24183 59062
rect 28625 58986 28691 58989
rect 31200 58986 32000 59016
rect 28625 58984 32000 58986
rect 28625 58928 28630 58984
rect 28686 58928 32000 58984
rect 28625 58926 32000 58928
rect 28625 58923 28691 58926
rect 31200 58896 32000 58926
rect 27153 58850 27219 58853
rect 28758 58850 28764 58852
rect 27153 58848 28764 58850
rect 27153 58792 27158 58848
rect 27214 58792 28764 58848
rect 27153 58790 28764 58792
rect 27153 58787 27219 58790
rect 28758 58788 28764 58790
rect 28828 58850 28834 58852
rect 28901 58850 28967 58853
rect 28828 58848 28967 58850
rect 28828 58792 28906 58848
rect 28962 58792 28967 58848
rect 28828 58790 28967 58792
rect 28828 58788 28834 58790
rect 28901 58787 28967 58790
rect 10874 58784 11194 58785
rect 10874 58720 10882 58784
rect 10946 58720 10962 58784
rect 11026 58720 11042 58784
rect 11106 58720 11122 58784
rect 11186 58720 11194 58784
rect 10874 58719 11194 58720
rect 20805 58784 21125 58785
rect 20805 58720 20813 58784
rect 20877 58720 20893 58784
rect 20957 58720 20973 58784
rect 21037 58720 21053 58784
rect 21117 58720 21125 58784
rect 20805 58719 21125 58720
rect 28625 58714 28691 58717
rect 28758 58714 28764 58716
rect 28625 58712 28764 58714
rect 28625 58656 28630 58712
rect 28686 58656 28764 58712
rect 28625 58654 28764 58656
rect 28625 58651 28691 58654
rect 28758 58652 28764 58654
rect 28828 58652 28834 58716
rect 26325 58576 26391 58581
rect 26325 58520 26330 58576
rect 26386 58520 26391 58576
rect 26325 58515 26391 58520
rect 27613 58578 27679 58581
rect 27838 58578 27844 58580
rect 27613 58576 27844 58578
rect 27613 58520 27618 58576
rect 27674 58520 27844 58576
rect 27613 58518 27844 58520
rect 27613 58515 27679 58518
rect 27838 58516 27844 58518
rect 27908 58516 27914 58580
rect 0 58442 800 58472
rect 1577 58442 1643 58445
rect 0 58440 1643 58442
rect 0 58384 1582 58440
rect 1638 58384 1643 58440
rect 0 58382 1643 58384
rect 0 58352 800 58382
rect 1577 58379 1643 58382
rect 5909 58240 6229 58241
rect 5909 58176 5917 58240
rect 5981 58176 5997 58240
rect 6061 58176 6077 58240
rect 6141 58176 6157 58240
rect 6221 58176 6229 58240
rect 5909 58175 6229 58176
rect 15840 58240 16160 58241
rect 15840 58176 15848 58240
rect 15912 58176 15928 58240
rect 15992 58176 16008 58240
rect 16072 58176 16088 58240
rect 16152 58176 16160 58240
rect 15840 58175 16160 58176
rect 25770 58240 26090 58241
rect 25770 58176 25778 58240
rect 25842 58176 25858 58240
rect 25922 58176 25938 58240
rect 26002 58176 26018 58240
rect 26082 58176 26090 58240
rect 25770 58175 26090 58176
rect 25957 58034 26023 58037
rect 26328 58034 26388 58515
rect 29821 58442 29887 58445
rect 31200 58442 32000 58472
rect 29821 58440 32000 58442
rect 29821 58384 29826 58440
rect 29882 58384 32000 58440
rect 29821 58382 32000 58384
rect 29821 58379 29887 58382
rect 31200 58352 32000 58382
rect 25957 58032 26388 58034
rect 25957 57976 25962 58032
rect 26018 57976 26388 58032
rect 25957 57974 26388 57976
rect 29729 58034 29795 58037
rect 31200 58034 32000 58064
rect 29729 58032 32000 58034
rect 29729 57976 29734 58032
rect 29790 57976 32000 58032
rect 29729 57974 32000 57976
rect 25957 57971 26023 57974
rect 29729 57971 29795 57974
rect 31200 57944 32000 57974
rect 27470 57836 27476 57900
rect 27540 57898 27546 57900
rect 29729 57898 29795 57901
rect 29862 57898 29868 57900
rect 27540 57896 29868 57898
rect 27540 57840 29734 57896
rect 29790 57840 29868 57896
rect 27540 57838 29868 57840
rect 27540 57836 27546 57838
rect 29729 57835 29795 57838
rect 29862 57836 29868 57838
rect 29932 57836 29938 57900
rect 0 57762 800 57792
rect 1577 57762 1643 57765
rect 27429 57764 27495 57765
rect 27429 57762 27476 57764
rect 0 57760 1643 57762
rect 0 57704 1582 57760
rect 1638 57704 1643 57760
rect 0 57702 1643 57704
rect 27384 57760 27476 57762
rect 27384 57704 27434 57760
rect 27384 57702 27476 57704
rect 0 57672 800 57702
rect 1577 57699 1643 57702
rect 27429 57700 27476 57702
rect 27540 57700 27546 57764
rect 27429 57699 27495 57700
rect 10874 57696 11194 57697
rect 10874 57632 10882 57696
rect 10946 57632 10962 57696
rect 11026 57632 11042 57696
rect 11106 57632 11122 57696
rect 11186 57632 11194 57696
rect 10874 57631 11194 57632
rect 20805 57696 21125 57697
rect 20805 57632 20813 57696
rect 20877 57632 20893 57696
rect 20957 57632 20973 57696
rect 21037 57632 21053 57696
rect 21117 57632 21125 57696
rect 20805 57631 21125 57632
rect 26182 57564 26188 57628
rect 26252 57626 26258 57628
rect 26325 57626 26391 57629
rect 26252 57624 26391 57626
rect 26252 57568 26330 57624
rect 26386 57568 26391 57624
rect 26252 57566 26391 57568
rect 26252 57564 26258 57566
rect 26325 57563 26391 57566
rect 26601 57626 26667 57629
rect 26918 57626 26924 57628
rect 26601 57624 26924 57626
rect 26601 57568 26606 57624
rect 26662 57568 26924 57624
rect 26601 57566 26924 57568
rect 26601 57563 26667 57566
rect 26918 57564 26924 57566
rect 26988 57564 26994 57628
rect 19793 57490 19859 57493
rect 20805 57490 20871 57493
rect 19793 57488 20871 57490
rect 19793 57432 19798 57488
rect 19854 57432 20810 57488
rect 20866 57432 20871 57488
rect 19793 57430 20871 57432
rect 19793 57427 19859 57430
rect 20805 57427 20871 57430
rect 26049 57490 26115 57493
rect 27429 57490 27495 57493
rect 26049 57488 27495 57490
rect 26049 57432 26054 57488
rect 26110 57432 27434 57488
rect 27490 57432 27495 57488
rect 26049 57430 27495 57432
rect 26049 57427 26115 57430
rect 27429 57427 27495 57430
rect 29729 57490 29795 57493
rect 31200 57490 32000 57520
rect 29729 57488 32000 57490
rect 29729 57432 29734 57488
rect 29790 57432 32000 57488
rect 29729 57430 32000 57432
rect 29729 57427 29795 57430
rect 31200 57400 32000 57430
rect 23974 57292 23980 57356
rect 24044 57354 24050 57356
rect 24117 57354 24183 57357
rect 24044 57352 24183 57354
rect 24044 57296 24122 57352
rect 24178 57296 24183 57352
rect 24044 57294 24183 57296
rect 24044 57292 24050 57294
rect 24117 57291 24183 57294
rect 25957 57354 26023 57357
rect 26366 57354 26372 57356
rect 25957 57352 26372 57354
rect 25957 57296 25962 57352
rect 26018 57296 26372 57352
rect 25957 57294 26372 57296
rect 25957 57291 26023 57294
rect 26366 57292 26372 57294
rect 26436 57292 26442 57356
rect 27337 57218 27403 57221
rect 27654 57218 27660 57220
rect 27337 57216 27660 57218
rect 27337 57160 27342 57216
rect 27398 57160 27660 57216
rect 27337 57158 27660 57160
rect 27337 57155 27403 57158
rect 27654 57156 27660 57158
rect 27724 57156 27730 57220
rect 28717 57216 28783 57221
rect 28717 57160 28722 57216
rect 28778 57160 28783 57216
rect 28717 57155 28783 57160
rect 29729 57218 29795 57221
rect 30649 57220 30715 57221
rect 30046 57218 30052 57220
rect 29729 57216 30052 57218
rect 29729 57160 29734 57216
rect 29790 57160 30052 57216
rect 29729 57158 30052 57160
rect 29729 57155 29795 57158
rect 30046 57156 30052 57158
rect 30116 57156 30122 57220
rect 30598 57156 30604 57220
rect 30668 57218 30715 57220
rect 30668 57216 30760 57218
rect 30710 57160 30760 57216
rect 30668 57158 30760 57160
rect 30668 57156 30715 57158
rect 30649 57155 30715 57156
rect 5909 57152 6229 57153
rect 0 57082 800 57112
rect 5909 57088 5917 57152
rect 5981 57088 5997 57152
rect 6061 57088 6077 57152
rect 6141 57088 6157 57152
rect 6221 57088 6229 57152
rect 5909 57087 6229 57088
rect 15840 57152 16160 57153
rect 15840 57088 15848 57152
rect 15912 57088 15928 57152
rect 15992 57088 16008 57152
rect 16072 57088 16088 57152
rect 16152 57088 16160 57152
rect 15840 57087 16160 57088
rect 25770 57152 26090 57153
rect 25770 57088 25778 57152
rect 25842 57088 25858 57152
rect 25922 57088 25938 57152
rect 26002 57088 26018 57152
rect 26082 57088 26090 57152
rect 25770 57087 26090 57088
rect 1577 57082 1643 57085
rect 0 57080 1643 57082
rect 0 57024 1582 57080
rect 1638 57024 1643 57080
rect 0 57022 1643 57024
rect 0 56992 800 57022
rect 1577 57019 1643 57022
rect 23473 57082 23539 57085
rect 27337 57082 27403 57085
rect 28165 57082 28231 57085
rect 23473 57080 25698 57082
rect 23473 57024 23478 57080
rect 23534 57024 25698 57080
rect 23473 57022 25698 57024
rect 23473 57019 23539 57022
rect 23422 56884 23428 56948
rect 23492 56946 23498 56948
rect 24577 56946 24643 56949
rect 23492 56944 24643 56946
rect 23492 56888 24582 56944
rect 24638 56888 24643 56944
rect 23492 56886 24643 56888
rect 25638 56946 25698 57022
rect 27337 57080 28231 57082
rect 27337 57024 27342 57080
rect 27398 57024 28170 57080
rect 28226 57024 28231 57080
rect 27337 57022 28231 57024
rect 28720 57082 28780 57155
rect 31200 57082 32000 57112
rect 28720 57022 32000 57082
rect 27337 57019 27403 57022
rect 28165 57019 28231 57022
rect 31200 56992 32000 57022
rect 26049 56946 26115 56949
rect 25638 56944 26115 56946
rect 25638 56888 26054 56944
rect 26110 56888 26115 56944
rect 25638 56886 26115 56888
rect 23492 56884 23498 56886
rect 24577 56883 24643 56886
rect 26049 56883 26115 56886
rect 28717 56946 28783 56949
rect 29494 56946 29500 56948
rect 28717 56944 29500 56946
rect 28717 56888 28722 56944
rect 28778 56888 29500 56944
rect 28717 56886 29500 56888
rect 28717 56883 28783 56886
rect 29494 56884 29500 56886
rect 29564 56884 29570 56948
rect 17350 56748 17356 56812
rect 17420 56810 17426 56812
rect 24393 56810 24459 56813
rect 17420 56808 24459 56810
rect 17420 56752 24398 56808
rect 24454 56752 24459 56808
rect 17420 56750 24459 56752
rect 17420 56748 17426 56750
rect 24393 56747 24459 56750
rect 28349 56810 28415 56813
rect 29126 56810 29132 56812
rect 28349 56808 29132 56810
rect 28349 56752 28354 56808
rect 28410 56752 29132 56808
rect 28349 56750 29132 56752
rect 28349 56747 28415 56750
rect 29126 56748 29132 56750
rect 29196 56748 29202 56812
rect 23565 56676 23631 56677
rect 23565 56674 23612 56676
rect 23520 56672 23612 56674
rect 23520 56616 23570 56672
rect 23520 56614 23612 56616
rect 23565 56612 23612 56614
rect 23676 56612 23682 56676
rect 25078 56612 25084 56676
rect 25148 56674 25154 56676
rect 25221 56674 25287 56677
rect 25148 56672 25287 56674
rect 25148 56616 25226 56672
rect 25282 56616 25287 56672
rect 25148 56614 25287 56616
rect 25148 56612 25154 56614
rect 23565 56611 23631 56612
rect 25221 56611 25287 56614
rect 28165 56674 28231 56677
rect 29361 56674 29427 56677
rect 28165 56672 29427 56674
rect 28165 56616 28170 56672
rect 28226 56616 29366 56672
rect 29422 56616 29427 56672
rect 28165 56614 29427 56616
rect 28165 56611 28231 56614
rect 29361 56611 29427 56614
rect 29913 56674 29979 56677
rect 31200 56674 32000 56704
rect 29913 56672 32000 56674
rect 29913 56616 29918 56672
rect 29974 56616 32000 56672
rect 29913 56614 32000 56616
rect 29913 56611 29979 56614
rect 10874 56608 11194 56609
rect 0 56538 800 56568
rect 10874 56544 10882 56608
rect 10946 56544 10962 56608
rect 11026 56544 11042 56608
rect 11106 56544 11122 56608
rect 11186 56544 11194 56608
rect 10874 56543 11194 56544
rect 20805 56608 21125 56609
rect 20805 56544 20813 56608
rect 20877 56544 20893 56608
rect 20957 56544 20973 56608
rect 21037 56544 21053 56608
rect 21117 56544 21125 56608
rect 31200 56584 32000 56614
rect 20805 56543 21125 56544
rect 1577 56538 1643 56541
rect 0 56536 1643 56538
rect 0 56480 1582 56536
rect 1638 56480 1643 56536
rect 0 56478 1643 56480
rect 0 56448 800 56478
rect 1577 56475 1643 56478
rect 23289 56538 23355 56541
rect 28165 56538 28231 56541
rect 23289 56536 28231 56538
rect 23289 56480 23294 56536
rect 23350 56480 28170 56536
rect 28226 56480 28231 56536
rect 23289 56478 28231 56480
rect 23289 56475 23355 56478
rect 28165 56475 28231 56478
rect 28625 56130 28691 56133
rect 31200 56130 32000 56160
rect 28625 56128 32000 56130
rect 28625 56072 28630 56128
rect 28686 56072 32000 56128
rect 28625 56070 32000 56072
rect 28625 56067 28691 56070
rect 5909 56064 6229 56065
rect 5909 56000 5917 56064
rect 5981 56000 5997 56064
rect 6061 56000 6077 56064
rect 6141 56000 6157 56064
rect 6221 56000 6229 56064
rect 5909 55999 6229 56000
rect 15840 56064 16160 56065
rect 15840 56000 15848 56064
rect 15912 56000 15928 56064
rect 15992 56000 16008 56064
rect 16072 56000 16088 56064
rect 16152 56000 16160 56064
rect 15840 55999 16160 56000
rect 25770 56064 26090 56065
rect 25770 56000 25778 56064
rect 25842 56000 25858 56064
rect 25922 56000 25938 56064
rect 26002 56000 26018 56064
rect 26082 56000 26090 56064
rect 31200 56040 32000 56070
rect 25770 55999 26090 56000
rect 26785 55994 26851 55997
rect 26785 55992 26986 55994
rect 26785 55936 26790 55992
rect 26846 55936 26986 55992
rect 26785 55934 26986 55936
rect 26785 55931 26851 55934
rect 0 55858 800 55888
rect 1577 55858 1643 55861
rect 23841 55860 23907 55861
rect 23790 55858 23796 55860
rect 0 55856 1643 55858
rect 0 55800 1582 55856
rect 1638 55800 1643 55856
rect 0 55798 1643 55800
rect 23750 55798 23796 55858
rect 23860 55856 23907 55860
rect 23902 55800 23907 55856
rect 0 55768 800 55798
rect 1577 55795 1643 55798
rect 23790 55796 23796 55798
rect 23860 55796 23907 55800
rect 24894 55796 24900 55860
rect 24964 55858 24970 55860
rect 25129 55858 25195 55861
rect 24964 55856 25195 55858
rect 24964 55800 25134 55856
rect 25190 55800 25195 55856
rect 24964 55798 25195 55800
rect 24964 55796 24970 55798
rect 23841 55795 23907 55796
rect 25129 55795 25195 55798
rect 25497 55858 25563 55861
rect 25957 55858 26023 55861
rect 25497 55856 26023 55858
rect 25497 55800 25502 55856
rect 25558 55800 25962 55856
rect 26018 55800 26023 55856
rect 25497 55798 26023 55800
rect 25497 55795 25563 55798
rect 25957 55795 26023 55798
rect 26926 55586 26986 55934
rect 30782 55660 30788 55724
rect 30852 55722 30858 55724
rect 31200 55722 32000 55752
rect 30852 55662 32000 55722
rect 30852 55660 30858 55662
rect 31200 55632 32000 55662
rect 27429 55586 27495 55589
rect 26926 55584 27495 55586
rect 26926 55528 27434 55584
rect 27490 55528 27495 55584
rect 26926 55526 27495 55528
rect 27429 55523 27495 55526
rect 28809 55586 28875 55589
rect 29177 55586 29243 55589
rect 28809 55584 29010 55586
rect 28809 55528 28814 55584
rect 28870 55528 29010 55584
rect 28809 55526 29010 55528
rect 28809 55523 28875 55526
rect 10874 55520 11194 55521
rect 10874 55456 10882 55520
rect 10946 55456 10962 55520
rect 11026 55456 11042 55520
rect 11106 55456 11122 55520
rect 11186 55456 11194 55520
rect 10874 55455 11194 55456
rect 20805 55520 21125 55521
rect 20805 55456 20813 55520
rect 20877 55456 20893 55520
rect 20957 55456 20973 55520
rect 21037 55456 21053 55520
rect 21117 55456 21125 55520
rect 20805 55455 21125 55456
rect 24209 55450 24275 55453
rect 25037 55450 25103 55453
rect 25865 55450 25931 55453
rect 24209 55448 25931 55450
rect 24209 55392 24214 55448
rect 24270 55392 25042 55448
rect 25098 55392 25870 55448
rect 25926 55392 25931 55448
rect 24209 55390 25931 55392
rect 24209 55387 24275 55390
rect 25037 55387 25103 55390
rect 25865 55387 25931 55390
rect 27286 55388 27292 55452
rect 27356 55450 27362 55452
rect 28717 55450 28783 55453
rect 27356 55448 28783 55450
rect 27356 55392 28722 55448
rect 28778 55392 28783 55448
rect 27356 55390 28783 55392
rect 27356 55388 27362 55390
rect 28717 55387 28783 55390
rect 9489 55314 9555 55317
rect 22829 55314 22895 55317
rect 23197 55314 23263 55317
rect 9489 55312 23263 55314
rect 9489 55256 9494 55312
rect 9550 55256 22834 55312
rect 22890 55256 23202 55312
rect 23258 55256 23263 55312
rect 9489 55254 23263 55256
rect 9489 55251 9555 55254
rect 22829 55251 22895 55254
rect 23197 55251 23263 55254
rect 25773 55314 25839 55317
rect 25773 55312 26250 55314
rect 25773 55256 25778 55312
rect 25834 55256 26250 55312
rect 25773 55254 26250 55256
rect 25773 55251 25839 55254
rect 0 55178 800 55208
rect 1577 55178 1643 55181
rect 0 55176 1643 55178
rect 0 55120 1582 55176
rect 1638 55120 1643 55176
rect 0 55118 1643 55120
rect 0 55088 800 55118
rect 1577 55115 1643 55118
rect 23197 55178 23263 55181
rect 23841 55178 23907 55181
rect 23197 55176 23907 55178
rect 23197 55120 23202 55176
rect 23258 55120 23846 55176
rect 23902 55120 23907 55176
rect 23197 55118 23907 55120
rect 23197 55115 23263 55118
rect 23841 55115 23907 55118
rect 24945 55178 25011 55181
rect 25957 55178 26023 55181
rect 24945 55176 26023 55178
rect 24945 55120 24950 55176
rect 25006 55120 25962 55176
rect 26018 55120 26023 55176
rect 24945 55118 26023 55120
rect 24945 55115 25011 55118
rect 25957 55115 26023 55118
rect 24577 55042 24643 55045
rect 25078 55042 25084 55044
rect 24577 55040 25084 55042
rect 24577 54984 24582 55040
rect 24638 54984 25084 55040
rect 24577 54982 25084 54984
rect 24577 54979 24643 54982
rect 25078 54980 25084 54982
rect 25148 54980 25154 55044
rect 5909 54976 6229 54977
rect 5909 54912 5917 54976
rect 5981 54912 5997 54976
rect 6061 54912 6077 54976
rect 6141 54912 6157 54976
rect 6221 54912 6229 54976
rect 5909 54911 6229 54912
rect 15840 54976 16160 54977
rect 15840 54912 15848 54976
rect 15912 54912 15928 54976
rect 15992 54912 16008 54976
rect 16072 54912 16088 54976
rect 16152 54912 16160 54976
rect 15840 54911 16160 54912
rect 25770 54976 26090 54977
rect 25770 54912 25778 54976
rect 25842 54912 25858 54976
rect 25922 54912 25938 54976
rect 26002 54912 26018 54976
rect 26082 54912 26090 54976
rect 25770 54911 26090 54912
rect 24209 54906 24275 54909
rect 24526 54906 24532 54908
rect 24209 54904 24532 54906
rect 24209 54848 24214 54904
rect 24270 54848 24532 54904
rect 24209 54846 24532 54848
rect 24209 54843 24275 54846
rect 24526 54844 24532 54846
rect 24596 54844 24602 54908
rect 24710 54844 24716 54908
rect 24780 54906 24786 54908
rect 25037 54906 25103 54909
rect 24780 54904 25103 54906
rect 24780 54848 25042 54904
rect 25098 54848 25103 54904
rect 24780 54846 25103 54848
rect 24780 54844 24786 54846
rect 25037 54843 25103 54846
rect 26190 54773 26250 55254
rect 28206 55252 28212 55316
rect 28276 55314 28282 55316
rect 28809 55314 28875 55317
rect 28276 55312 28875 55314
rect 28276 55256 28814 55312
rect 28870 55256 28875 55312
rect 28276 55254 28875 55256
rect 28276 55252 28282 55254
rect 28809 55251 28875 55254
rect 28809 55178 28875 55181
rect 28950 55178 29010 55526
rect 28809 55176 29010 55178
rect 28809 55120 28814 55176
rect 28870 55120 29010 55176
rect 28809 55118 29010 55120
rect 29134 55584 29243 55586
rect 29134 55528 29182 55584
rect 29238 55528 29243 55584
rect 29134 55523 29243 55528
rect 28809 55115 28875 55118
rect 26141 54768 26250 54773
rect 26141 54712 26146 54768
rect 26202 54712 26250 54768
rect 26141 54710 26250 54712
rect 26969 54770 27035 54773
rect 27102 54770 27108 54772
rect 26969 54768 27108 54770
rect 26969 54712 26974 54768
rect 27030 54712 27108 54768
rect 26969 54710 27108 54712
rect 26141 54707 26207 54710
rect 26969 54707 27035 54710
rect 27102 54708 27108 54710
rect 27172 54708 27178 54772
rect 27429 54634 27495 54637
rect 28574 54634 28580 54636
rect 27429 54632 28580 54634
rect 27429 54576 27434 54632
rect 27490 54576 28580 54632
rect 27429 54574 28580 54576
rect 27429 54571 27495 54574
rect 28574 54572 28580 54574
rect 28644 54572 28650 54636
rect 0 54498 800 54528
rect 1577 54498 1643 54501
rect 0 54496 1643 54498
rect 0 54440 1582 54496
rect 1638 54440 1643 54496
rect 0 54438 1643 54440
rect 0 54408 800 54438
rect 1577 54435 1643 54438
rect 27429 54498 27495 54501
rect 29134 54498 29194 55523
rect 29913 55314 29979 55317
rect 30281 55314 30347 55317
rect 29913 55312 30347 55314
rect 29913 55256 29918 55312
rect 29974 55256 30286 55312
rect 30342 55256 30347 55312
rect 29913 55254 30347 55256
rect 29913 55251 29979 55254
rect 30281 55251 30347 55254
rect 29729 55178 29795 55181
rect 31200 55178 32000 55208
rect 29729 55176 32000 55178
rect 29729 55120 29734 55176
rect 29790 55120 32000 55176
rect 29729 55118 32000 55120
rect 29729 55115 29795 55118
rect 31200 55088 32000 55118
rect 30046 54980 30052 55044
rect 30116 55042 30122 55044
rect 30925 55042 30991 55045
rect 30116 55040 30991 55042
rect 30116 54984 30930 55040
rect 30986 54984 30991 55040
rect 30116 54982 30991 54984
rect 30116 54980 30122 54982
rect 30925 54979 30991 54982
rect 29729 54770 29795 54773
rect 31200 54770 32000 54800
rect 29729 54768 32000 54770
rect 29729 54712 29734 54768
rect 29790 54712 32000 54768
rect 29729 54710 32000 54712
rect 29729 54707 29795 54710
rect 31200 54680 32000 54710
rect 27429 54496 29194 54498
rect 27429 54440 27434 54496
rect 27490 54440 29194 54496
rect 27429 54438 29194 54440
rect 30281 54498 30347 54501
rect 31518 54498 31524 54500
rect 30281 54496 31524 54498
rect 30281 54440 30286 54496
rect 30342 54440 31524 54496
rect 30281 54438 31524 54440
rect 27429 54435 27495 54438
rect 30281 54435 30347 54438
rect 31518 54436 31524 54438
rect 31588 54436 31594 54500
rect 10874 54432 11194 54433
rect 10874 54368 10882 54432
rect 10946 54368 10962 54432
rect 11026 54368 11042 54432
rect 11106 54368 11122 54432
rect 11186 54368 11194 54432
rect 10874 54367 11194 54368
rect 20805 54432 21125 54433
rect 20805 54368 20813 54432
rect 20877 54368 20893 54432
rect 20957 54368 20973 54432
rect 21037 54368 21053 54432
rect 21117 54368 21125 54432
rect 20805 54367 21125 54368
rect 26141 54362 26207 54365
rect 26366 54362 26372 54364
rect 26141 54360 26372 54362
rect 26141 54304 26146 54360
rect 26202 54304 26372 54360
rect 26141 54302 26372 54304
rect 26141 54299 26207 54302
rect 26366 54300 26372 54302
rect 26436 54300 26442 54364
rect 26049 54226 26115 54229
rect 26366 54226 26372 54228
rect 26049 54224 26372 54226
rect 26049 54168 26054 54224
rect 26110 54168 26372 54224
rect 26049 54166 26372 54168
rect 26049 54163 26115 54166
rect 26366 54164 26372 54166
rect 26436 54164 26442 54228
rect 28625 54226 28691 54229
rect 31200 54226 32000 54256
rect 28625 54224 32000 54226
rect 28625 54168 28630 54224
rect 28686 54168 32000 54224
rect 28625 54166 32000 54168
rect 28625 54163 28691 54166
rect 31200 54136 32000 54166
rect 25221 54092 25287 54093
rect 25221 54090 25268 54092
rect 25176 54088 25268 54090
rect 25176 54032 25226 54088
rect 25176 54030 25268 54032
rect 25221 54028 25268 54030
rect 25332 54028 25338 54092
rect 28758 54028 28764 54092
rect 28828 54090 28834 54092
rect 29453 54090 29519 54093
rect 28828 54088 29519 54090
rect 28828 54032 29458 54088
rect 29514 54032 29519 54088
rect 28828 54030 29519 54032
rect 28828 54028 28834 54030
rect 25221 54027 25287 54028
rect 29453 54027 29519 54030
rect 5909 53888 6229 53889
rect 0 53818 800 53848
rect 5909 53824 5917 53888
rect 5981 53824 5997 53888
rect 6061 53824 6077 53888
rect 6141 53824 6157 53888
rect 6221 53824 6229 53888
rect 5909 53823 6229 53824
rect 15840 53888 16160 53889
rect 15840 53824 15848 53888
rect 15912 53824 15928 53888
rect 15992 53824 16008 53888
rect 16072 53824 16088 53888
rect 16152 53824 16160 53888
rect 15840 53823 16160 53824
rect 25770 53888 26090 53889
rect 25770 53824 25778 53888
rect 25842 53824 25858 53888
rect 25922 53824 25938 53888
rect 26002 53824 26018 53888
rect 26082 53824 26090 53888
rect 25770 53823 26090 53824
rect 1577 53818 1643 53821
rect 27889 53820 27955 53821
rect 0 53816 1643 53818
rect 0 53760 1582 53816
rect 1638 53760 1643 53816
rect 0 53758 1643 53760
rect 0 53728 800 53758
rect 1577 53755 1643 53758
rect 19190 53756 19196 53820
rect 19260 53818 19266 53820
rect 23606 53818 23612 53820
rect 19260 53758 23612 53818
rect 19260 53756 19266 53758
rect 23606 53756 23612 53758
rect 23676 53756 23682 53820
rect 27838 53818 27844 53820
rect 27798 53758 27844 53818
rect 27908 53816 27955 53820
rect 27950 53760 27955 53816
rect 27838 53756 27844 53758
rect 27908 53756 27955 53760
rect 27889 53755 27955 53756
rect 29729 53818 29795 53821
rect 31200 53818 32000 53848
rect 29729 53816 32000 53818
rect 29729 53760 29734 53816
rect 29790 53760 32000 53816
rect 29729 53758 32000 53760
rect 29729 53755 29795 53758
rect 31200 53728 32000 53758
rect 17534 53620 17540 53684
rect 17604 53682 17610 53684
rect 23841 53682 23907 53685
rect 17604 53680 23907 53682
rect 17604 53624 23846 53680
rect 23902 53624 23907 53680
rect 17604 53622 23907 53624
rect 17604 53620 17610 53622
rect 23841 53619 23907 53622
rect 29494 53620 29500 53684
rect 29564 53682 29570 53684
rect 29637 53682 29703 53685
rect 29564 53680 29703 53682
rect 29564 53624 29642 53680
rect 29698 53624 29703 53680
rect 29564 53622 29703 53624
rect 29564 53620 29570 53622
rect 29637 53619 29703 53622
rect 29177 53546 29243 53549
rect 30230 53546 30236 53548
rect 29177 53544 30236 53546
rect 29177 53488 29182 53544
rect 29238 53488 30236 53544
rect 29177 53486 30236 53488
rect 29177 53483 29243 53486
rect 30230 53484 30236 53486
rect 30300 53484 30306 53548
rect 24025 53410 24091 53413
rect 28390 53410 28396 53412
rect 24025 53408 28396 53410
rect 24025 53352 24030 53408
rect 24086 53352 28396 53408
rect 24025 53350 28396 53352
rect 24025 53347 24091 53350
rect 28390 53348 28396 53350
rect 28460 53348 28466 53412
rect 28942 53348 28948 53412
rect 29012 53410 29018 53412
rect 29085 53410 29151 53413
rect 29012 53408 29151 53410
rect 29012 53352 29090 53408
rect 29146 53352 29151 53408
rect 29012 53350 29151 53352
rect 29012 53348 29018 53350
rect 29085 53347 29151 53350
rect 10874 53344 11194 53345
rect 10874 53280 10882 53344
rect 10946 53280 10962 53344
rect 11026 53280 11042 53344
rect 11106 53280 11122 53344
rect 11186 53280 11194 53344
rect 10874 53279 11194 53280
rect 20805 53344 21125 53345
rect 20805 53280 20813 53344
rect 20877 53280 20893 53344
rect 20957 53280 20973 53344
rect 21037 53280 21053 53344
rect 21117 53280 21125 53344
rect 20805 53279 21125 53280
rect 27705 53274 27771 53277
rect 31200 53274 32000 53304
rect 27705 53272 32000 53274
rect 27705 53216 27710 53272
rect 27766 53216 32000 53272
rect 27705 53214 32000 53216
rect 27705 53211 27771 53214
rect 31200 53184 32000 53214
rect 0 53138 800 53168
rect 1577 53138 1643 53141
rect 0 53136 1643 53138
rect 0 53080 1582 53136
rect 1638 53080 1643 53136
rect 0 53078 1643 53080
rect 0 53048 800 53078
rect 1577 53075 1643 53078
rect 25957 53138 26023 53141
rect 29269 53140 29335 53141
rect 28758 53138 28764 53140
rect 25957 53136 28764 53138
rect 25957 53080 25962 53136
rect 26018 53080 28764 53136
rect 25957 53078 28764 53080
rect 25957 53075 26023 53078
rect 28758 53076 28764 53078
rect 28828 53076 28834 53140
rect 29269 53136 29316 53140
rect 29380 53138 29386 53140
rect 30005 53138 30071 53141
rect 30782 53138 30788 53140
rect 29269 53080 29274 53136
rect 29269 53076 29316 53080
rect 29380 53078 29426 53138
rect 30005 53136 30788 53138
rect 30005 53080 30010 53136
rect 30066 53080 30788 53136
rect 30005 53078 30788 53080
rect 29380 53076 29386 53078
rect 29269 53075 29335 53076
rect 30005 53075 30071 53078
rect 30782 53076 30788 53078
rect 30852 53076 30858 53140
rect 23657 53002 23723 53005
rect 24158 53002 24164 53004
rect 23657 53000 24164 53002
rect 23657 52944 23662 53000
rect 23718 52944 24164 53000
rect 23657 52942 24164 52944
rect 23657 52939 23723 52942
rect 24158 52940 24164 52942
rect 24228 52940 24234 53004
rect 26325 53002 26391 53005
rect 27102 53002 27108 53004
rect 26325 53000 27108 53002
rect 26325 52944 26330 53000
rect 26386 52944 27108 53000
rect 26325 52942 27108 52944
rect 26325 52939 26391 52942
rect 27102 52940 27108 52942
rect 27172 52940 27178 53004
rect 28022 52940 28028 53004
rect 28092 53002 28098 53004
rect 28901 53002 28967 53005
rect 29637 53002 29703 53005
rect 28092 53000 29703 53002
rect 28092 52944 28906 53000
rect 28962 52944 29642 53000
rect 29698 52944 29703 53000
rect 28092 52942 29703 52944
rect 28092 52940 28098 52942
rect 28901 52939 28967 52942
rect 29637 52939 29703 52942
rect 23238 52804 23244 52868
rect 23308 52866 23314 52868
rect 23657 52866 23723 52869
rect 23308 52864 23723 52866
rect 23308 52808 23662 52864
rect 23718 52808 23723 52864
rect 23308 52806 23723 52808
rect 23308 52804 23314 52806
rect 23657 52803 23723 52806
rect 27981 52866 28047 52869
rect 31200 52866 32000 52896
rect 27981 52864 32000 52866
rect 27981 52808 27986 52864
rect 28042 52808 32000 52864
rect 27981 52806 32000 52808
rect 27981 52803 28047 52806
rect 5909 52800 6229 52801
rect 5909 52736 5917 52800
rect 5981 52736 5997 52800
rect 6061 52736 6077 52800
rect 6141 52736 6157 52800
rect 6221 52736 6229 52800
rect 5909 52735 6229 52736
rect 15840 52800 16160 52801
rect 15840 52736 15848 52800
rect 15912 52736 15928 52800
rect 15992 52736 16008 52800
rect 16072 52736 16088 52800
rect 16152 52736 16160 52800
rect 15840 52735 16160 52736
rect 25770 52800 26090 52801
rect 25770 52736 25778 52800
rect 25842 52736 25858 52800
rect 25922 52736 25938 52800
rect 26002 52736 26018 52800
rect 26082 52736 26090 52800
rect 31200 52776 32000 52806
rect 25770 52735 26090 52736
rect 27981 52732 28047 52733
rect 27981 52728 28028 52732
rect 28092 52730 28098 52732
rect 27981 52672 27986 52728
rect 27981 52668 28028 52672
rect 28092 52670 28138 52730
rect 28092 52668 28098 52670
rect 28390 52668 28396 52732
rect 28460 52730 28466 52732
rect 28625 52730 28691 52733
rect 28460 52728 28691 52730
rect 28460 52672 28630 52728
rect 28686 52672 28691 52728
rect 28460 52670 28691 52672
rect 28460 52668 28466 52670
rect 27981 52667 28047 52668
rect 28625 52667 28691 52670
rect 29269 52730 29335 52733
rect 30414 52730 30420 52732
rect 29269 52728 30420 52730
rect 29269 52672 29274 52728
rect 29330 52672 30420 52728
rect 29269 52670 30420 52672
rect 29269 52667 29335 52670
rect 30414 52668 30420 52670
rect 30484 52668 30490 52732
rect 27613 52594 27679 52597
rect 29361 52596 29427 52597
rect 29310 52594 29316 52596
rect 27613 52592 28458 52594
rect 27613 52536 27618 52592
rect 27674 52536 28458 52592
rect 27613 52534 28458 52536
rect 29270 52534 29316 52594
rect 29380 52592 29427 52596
rect 29422 52536 29427 52592
rect 27613 52531 27679 52534
rect 0 52458 800 52488
rect 2037 52458 2103 52461
rect 0 52456 2103 52458
rect 0 52400 2042 52456
rect 2098 52400 2103 52456
rect 0 52398 2103 52400
rect 0 52368 800 52398
rect 2037 52395 2103 52398
rect 23606 52396 23612 52460
rect 23676 52458 23682 52460
rect 27613 52458 27679 52461
rect 23676 52456 27679 52458
rect 23676 52400 27618 52456
rect 27674 52400 27679 52456
rect 23676 52398 27679 52400
rect 23676 52396 23682 52398
rect 27613 52395 27679 52398
rect 23933 52322 23999 52325
rect 26550 52322 26556 52324
rect 23933 52320 26556 52322
rect 23933 52264 23938 52320
rect 23994 52264 26556 52320
rect 23933 52262 26556 52264
rect 23933 52259 23999 52262
rect 26550 52260 26556 52262
rect 26620 52260 26626 52324
rect 10874 52256 11194 52257
rect 10874 52192 10882 52256
rect 10946 52192 10962 52256
rect 11026 52192 11042 52256
rect 11106 52192 11122 52256
rect 11186 52192 11194 52256
rect 10874 52191 11194 52192
rect 20805 52256 21125 52257
rect 20805 52192 20813 52256
rect 20877 52192 20893 52256
rect 20957 52192 20973 52256
rect 21037 52192 21053 52256
rect 21117 52192 21125 52256
rect 20805 52191 21125 52192
rect 26550 52124 26556 52188
rect 26620 52186 26626 52188
rect 27286 52186 27292 52188
rect 26620 52126 27292 52186
rect 26620 52124 26626 52126
rect 27286 52124 27292 52126
rect 27356 52124 27362 52188
rect 26601 52048 26667 52053
rect 26601 51992 26606 52048
rect 26662 51992 26667 52048
rect 26601 51987 26667 51992
rect 27286 51988 27292 52052
rect 27356 52050 27362 52052
rect 27654 52050 27660 52052
rect 27356 51990 27660 52050
rect 27356 51988 27362 51990
rect 27654 51988 27660 51990
rect 27724 51988 27730 52052
rect 0 51914 800 51944
rect 1577 51914 1643 51917
rect 0 51912 1643 51914
rect 0 51856 1582 51912
rect 1638 51856 1643 51912
rect 0 51854 1643 51856
rect 0 51824 800 51854
rect 1577 51851 1643 51854
rect 26604 51778 26664 51987
rect 28398 51917 28458 52534
rect 29310 52532 29316 52534
rect 29380 52532 29427 52536
rect 29361 52531 29427 52532
rect 28758 52396 28764 52460
rect 28828 52458 28834 52460
rect 29453 52458 29519 52461
rect 28828 52456 29519 52458
rect 28828 52400 29458 52456
rect 29514 52400 29519 52456
rect 28828 52398 29519 52400
rect 28828 52396 28834 52398
rect 29453 52395 29519 52398
rect 28717 52322 28783 52325
rect 31200 52322 32000 52352
rect 28717 52320 32000 52322
rect 28717 52264 28722 52320
rect 28778 52264 32000 52320
rect 28717 52262 32000 52264
rect 28717 52259 28783 52262
rect 31200 52232 32000 52262
rect 28625 52186 28691 52189
rect 28942 52186 28948 52188
rect 28625 52184 28948 52186
rect 28625 52128 28630 52184
rect 28686 52128 28948 52184
rect 28625 52126 28948 52128
rect 28625 52123 28691 52126
rect 28942 52124 28948 52126
rect 29012 52124 29018 52188
rect 29177 52186 29243 52189
rect 30230 52186 30236 52188
rect 29177 52184 30236 52186
rect 29177 52128 29182 52184
rect 29238 52128 30236 52184
rect 29177 52126 30236 52128
rect 29177 52123 29243 52126
rect 30230 52124 30236 52126
rect 30300 52124 30306 52188
rect 30465 52184 30531 52189
rect 30465 52128 30470 52184
rect 30526 52128 30531 52184
rect 30465 52123 30531 52128
rect 28717 52050 28783 52053
rect 28582 52048 28783 52050
rect 28582 51992 28722 52048
rect 28778 51992 28783 52048
rect 28582 51990 28783 51992
rect 26918 51852 26924 51916
rect 26988 51914 26994 51916
rect 27654 51914 27660 51916
rect 26988 51854 27660 51914
rect 26988 51852 26994 51854
rect 27654 51852 27660 51854
rect 27724 51852 27730 51916
rect 28398 51912 28507 51917
rect 28398 51856 28446 51912
rect 28502 51856 28507 51912
rect 28398 51854 28507 51856
rect 28441 51851 28507 51854
rect 28582 51778 28642 51990
rect 28717 51987 28783 51990
rect 29085 52050 29151 52053
rect 30468 52050 30528 52123
rect 29085 52048 30528 52050
rect 29085 51992 29090 52048
rect 29146 51992 30528 52048
rect 29085 51990 30528 51992
rect 29085 51987 29151 51990
rect 28717 51914 28783 51917
rect 31200 51914 32000 51944
rect 28717 51912 32000 51914
rect 28717 51856 28722 51912
rect 28778 51856 32000 51912
rect 28717 51854 32000 51856
rect 28717 51851 28783 51854
rect 31200 51824 32000 51854
rect 26604 51718 28642 51778
rect 29545 51778 29611 51781
rect 29862 51778 29868 51780
rect 29545 51776 29868 51778
rect 29545 51720 29550 51776
rect 29606 51720 29868 51776
rect 29545 51718 29868 51720
rect 29545 51715 29611 51718
rect 29862 51716 29868 51718
rect 29932 51716 29938 51780
rect 5909 51712 6229 51713
rect 5909 51648 5917 51712
rect 5981 51648 5997 51712
rect 6061 51648 6077 51712
rect 6141 51648 6157 51712
rect 6221 51648 6229 51712
rect 5909 51647 6229 51648
rect 15840 51712 16160 51713
rect 15840 51648 15848 51712
rect 15912 51648 15928 51712
rect 15992 51648 16008 51712
rect 16072 51648 16088 51712
rect 16152 51648 16160 51712
rect 15840 51647 16160 51648
rect 25770 51712 26090 51713
rect 25770 51648 25778 51712
rect 25842 51648 25858 51712
rect 25922 51648 25938 51712
rect 26002 51648 26018 51712
rect 26082 51648 26090 51712
rect 25770 51647 26090 51648
rect 24342 51580 24348 51644
rect 24412 51642 24418 51644
rect 24945 51642 25011 51645
rect 29913 51644 29979 51645
rect 29862 51642 29868 51644
rect 24412 51640 25011 51642
rect 24412 51584 24950 51640
rect 25006 51584 25011 51640
rect 24412 51582 25011 51584
rect 29822 51582 29868 51642
rect 29932 51640 29979 51644
rect 29974 51584 29979 51640
rect 24412 51580 24418 51582
rect 24945 51579 25011 51582
rect 29862 51580 29868 51582
rect 29932 51580 29979 51584
rect 29913 51579 29979 51580
rect 23841 51506 23907 51509
rect 23974 51506 23980 51508
rect 23841 51504 23980 51506
rect 23841 51448 23846 51504
rect 23902 51448 23980 51504
rect 23841 51446 23980 51448
rect 23841 51443 23907 51446
rect 23974 51444 23980 51446
rect 24044 51444 24050 51508
rect 29729 51506 29795 51509
rect 31200 51506 32000 51536
rect 29729 51504 32000 51506
rect 29729 51448 29734 51504
rect 29790 51448 32000 51504
rect 29729 51446 32000 51448
rect 29729 51443 29795 51446
rect 31200 51416 32000 51446
rect 14549 51370 14615 51373
rect 15101 51370 15167 51373
rect 23473 51372 23539 51373
rect 23422 51370 23428 51372
rect 14549 51368 15167 51370
rect 14549 51312 14554 51368
rect 14610 51312 15106 51368
rect 15162 51312 15167 51368
rect 14549 51310 15167 51312
rect 23382 51310 23428 51370
rect 23492 51368 23539 51372
rect 23534 51312 23539 51368
rect 14549 51307 14615 51310
rect 15101 51307 15167 51310
rect 23422 51308 23428 51310
rect 23492 51308 23539 51312
rect 23606 51308 23612 51372
rect 23676 51370 23682 51372
rect 24577 51370 24643 51373
rect 26366 51370 26372 51372
rect 23676 51368 24643 51370
rect 23676 51312 24582 51368
rect 24638 51312 24643 51368
rect 23676 51310 24643 51312
rect 23676 51308 23682 51310
rect 23473 51307 23539 51308
rect 24577 51307 24643 51310
rect 25822 51310 26372 51370
rect 0 51234 800 51264
rect 2221 51234 2287 51237
rect 25630 51234 25636 51236
rect 0 51232 2287 51234
rect 0 51176 2226 51232
rect 2282 51176 2287 51232
rect 0 51174 2287 51176
rect 0 51144 800 51174
rect 2221 51171 2287 51174
rect 25454 51174 25636 51234
rect 10874 51168 11194 51169
rect 10874 51104 10882 51168
rect 10946 51104 10962 51168
rect 11026 51104 11042 51168
rect 11106 51104 11122 51168
rect 11186 51104 11194 51168
rect 10874 51103 11194 51104
rect 20805 51168 21125 51169
rect 20805 51104 20813 51168
rect 20877 51104 20893 51168
rect 20957 51104 20973 51168
rect 21037 51104 21053 51168
rect 21117 51104 21125 51168
rect 20805 51103 21125 51104
rect 24485 51100 24551 51101
rect 24485 51096 24532 51100
rect 24596 51098 24602 51100
rect 25129 51098 25195 51101
rect 25454 51098 25514 51174
rect 25630 51172 25636 51174
rect 25700 51172 25706 51236
rect 25822 51101 25882 51310
rect 26366 51308 26372 51310
rect 26436 51308 26442 51372
rect 27102 51308 27108 51372
rect 27172 51370 27178 51372
rect 28625 51370 28691 51373
rect 29361 51372 29427 51373
rect 27172 51368 28691 51370
rect 27172 51312 28630 51368
rect 28686 51312 28691 51368
rect 27172 51310 28691 51312
rect 27172 51308 27178 51310
rect 28625 51307 28691 51310
rect 29310 51308 29316 51372
rect 29380 51370 29427 51372
rect 29637 51372 29703 51373
rect 29380 51368 29472 51370
rect 29422 51312 29472 51368
rect 29380 51310 29472 51312
rect 29637 51368 29684 51372
rect 29748 51370 29754 51372
rect 29637 51312 29642 51368
rect 29380 51308 29427 51310
rect 29361 51307 29427 51308
rect 29637 51308 29684 51312
rect 29748 51310 29794 51370
rect 29748 51308 29754 51310
rect 29637 51307 29703 51308
rect 26417 51236 26483 51237
rect 26366 51234 26372 51236
rect 26326 51174 26372 51234
rect 26436 51232 26483 51236
rect 27797 51236 27863 51237
rect 27797 51234 27844 51236
rect 26478 51176 26483 51232
rect 26366 51172 26372 51174
rect 26436 51172 26483 51176
rect 27752 51232 27844 51234
rect 27752 51176 27802 51232
rect 27752 51174 27844 51176
rect 26417 51171 26483 51172
rect 27797 51172 27844 51174
rect 27908 51172 27914 51236
rect 28390 51172 28396 51236
rect 28460 51234 28466 51236
rect 28901 51234 28967 51237
rect 28460 51232 28967 51234
rect 28460 51176 28906 51232
rect 28962 51176 28967 51232
rect 28460 51174 28967 51176
rect 28460 51172 28466 51174
rect 27797 51171 27863 51172
rect 28901 51171 28967 51174
rect 29177 51234 29243 51237
rect 30046 51234 30052 51236
rect 29177 51232 30052 51234
rect 29177 51176 29182 51232
rect 29238 51176 30052 51232
rect 29177 51174 30052 51176
rect 29177 51171 29243 51174
rect 30046 51172 30052 51174
rect 30116 51172 30122 51236
rect 30782 51172 30788 51236
rect 30852 51234 30858 51236
rect 30925 51234 30991 51237
rect 30852 51232 30991 51234
rect 30852 51176 30930 51232
rect 30986 51176 30991 51232
rect 30852 51174 30991 51176
rect 30852 51172 30858 51174
rect 30925 51171 30991 51174
rect 31150 51172 31156 51236
rect 31220 51234 31226 51236
rect 31293 51234 31359 51237
rect 31220 51232 31359 51234
rect 31220 51176 31298 51232
rect 31354 51176 31359 51232
rect 31220 51174 31359 51176
rect 31220 51172 31226 51174
rect 31293 51171 31359 51174
rect 21541 51090 21607 51093
rect 21406 51088 21607 51090
rect 21406 51032 21546 51088
rect 21602 51032 21607 51088
rect 24485 51040 24490 51096
rect 24485 51036 24532 51040
rect 24596 51038 24642 51098
rect 25129 51096 25514 51098
rect 25129 51040 25134 51096
rect 25190 51040 25514 51096
rect 25129 51038 25514 51040
rect 25773 51096 25882 51101
rect 25773 51040 25778 51096
rect 25834 51040 25882 51096
rect 25773 51038 25882 51040
rect 27705 51098 27771 51101
rect 28165 51098 28231 51101
rect 29085 51100 29151 51101
rect 29085 51098 29132 51100
rect 27705 51096 28231 51098
rect 27705 51040 27710 51096
rect 27766 51040 28170 51096
rect 28226 51040 28231 51096
rect 27705 51038 28231 51040
rect 29040 51096 29132 51098
rect 29040 51040 29090 51096
rect 29040 51038 29132 51040
rect 24596 51036 24602 51038
rect 24485 51035 24551 51036
rect 25129 51035 25195 51038
rect 25773 51035 25839 51038
rect 27705 51035 27771 51038
rect 28165 51035 28231 51038
rect 29085 51036 29132 51038
rect 29196 51036 29202 51100
rect 29085 51035 29151 51036
rect 21406 51030 21607 51032
rect 21081 50962 21147 50965
rect 21406 50964 21466 51030
rect 21541 51027 21607 51030
rect 21398 50962 21404 50964
rect 21081 50960 21404 50962
rect 21081 50904 21086 50960
rect 21142 50904 21404 50960
rect 21081 50902 21404 50904
rect 21081 50899 21147 50902
rect 21398 50900 21404 50902
rect 21468 50900 21474 50964
rect 21541 50962 21607 50965
rect 22001 50962 22067 50965
rect 21541 50960 22067 50962
rect 21541 50904 21546 50960
rect 21602 50904 22006 50960
rect 22062 50904 22067 50960
rect 21541 50902 22067 50904
rect 21541 50899 21607 50902
rect 22001 50899 22067 50902
rect 23749 50962 23815 50965
rect 24158 50962 24164 50964
rect 23749 50960 24164 50962
rect 23749 50904 23754 50960
rect 23810 50904 24164 50960
rect 23749 50902 24164 50904
rect 23749 50899 23815 50902
rect 24158 50900 24164 50902
rect 24228 50900 24234 50964
rect 24526 50900 24532 50964
rect 24596 50962 24602 50964
rect 24853 50962 24919 50965
rect 24596 50960 24919 50962
rect 24596 50904 24858 50960
rect 24914 50904 24919 50960
rect 24596 50902 24919 50904
rect 24596 50900 24602 50902
rect 24853 50899 24919 50902
rect 27654 50900 27660 50964
rect 27724 50962 27730 50964
rect 27981 50962 28047 50965
rect 30465 50964 30531 50965
rect 30414 50962 30420 50964
rect 27724 50960 28047 50962
rect 27724 50904 27986 50960
rect 28042 50904 28047 50960
rect 27724 50902 28047 50904
rect 30374 50902 30420 50962
rect 30484 50960 30531 50964
rect 30526 50904 30531 50960
rect 27724 50900 27730 50902
rect 27981 50899 28047 50902
rect 30414 50900 30420 50902
rect 30484 50900 30531 50904
rect 30465 50899 30531 50900
rect 30925 50964 30991 50965
rect 30925 50960 30972 50964
rect 31036 50962 31042 50964
rect 31200 50962 32000 50992
rect 30925 50904 30930 50960
rect 30925 50900 30972 50904
rect 31036 50902 31082 50962
rect 31036 50900 31042 50902
rect 30925 50899 30991 50900
rect 31158 50872 32000 50962
rect 17718 50764 17724 50828
rect 17788 50826 17794 50828
rect 25773 50826 25839 50829
rect 17788 50824 25839 50826
rect 17788 50768 25778 50824
rect 25834 50768 25839 50824
rect 17788 50766 25839 50768
rect 17788 50764 17794 50766
rect 25773 50763 25839 50766
rect 29913 50826 29979 50829
rect 31158 50826 31218 50872
rect 29913 50824 31218 50826
rect 29913 50768 29918 50824
rect 29974 50768 31218 50824
rect 29913 50766 31218 50768
rect 29913 50763 29979 50766
rect 24710 50628 24716 50692
rect 24780 50690 24786 50692
rect 24853 50690 24919 50693
rect 29821 50692 29887 50693
rect 29821 50690 29868 50692
rect 24780 50688 24919 50690
rect 24780 50632 24858 50688
rect 24914 50632 24919 50688
rect 24780 50630 24919 50632
rect 29776 50688 29868 50690
rect 29776 50632 29826 50688
rect 29776 50630 29868 50632
rect 24780 50628 24786 50630
rect 24853 50627 24919 50630
rect 29821 50628 29868 50630
rect 29932 50628 29938 50692
rect 30465 50690 30531 50693
rect 30782 50690 30788 50692
rect 30465 50688 30788 50690
rect 30465 50632 30470 50688
rect 30526 50632 30788 50688
rect 30465 50630 30788 50632
rect 29821 50627 29887 50628
rect 30465 50627 30531 50630
rect 30782 50628 30788 50630
rect 30852 50628 30858 50692
rect 5909 50624 6229 50625
rect 0 50554 800 50584
rect 5909 50560 5917 50624
rect 5981 50560 5997 50624
rect 6061 50560 6077 50624
rect 6141 50560 6157 50624
rect 6221 50560 6229 50624
rect 5909 50559 6229 50560
rect 15840 50624 16160 50625
rect 15840 50560 15848 50624
rect 15912 50560 15928 50624
rect 15992 50560 16008 50624
rect 16072 50560 16088 50624
rect 16152 50560 16160 50624
rect 15840 50559 16160 50560
rect 25770 50624 26090 50625
rect 25770 50560 25778 50624
rect 25842 50560 25858 50624
rect 25922 50560 25938 50624
rect 26002 50560 26018 50624
rect 26082 50560 26090 50624
rect 25770 50559 26090 50560
rect 1393 50554 1459 50557
rect 0 50552 1459 50554
rect 0 50496 1398 50552
rect 1454 50496 1459 50552
rect 0 50494 1459 50496
rect 0 50464 800 50494
rect 1393 50491 1459 50494
rect 24526 50492 24532 50556
rect 24596 50554 24602 50556
rect 24853 50554 24919 50557
rect 24596 50552 24919 50554
rect 24596 50496 24858 50552
rect 24914 50496 24919 50552
rect 24596 50494 24919 50496
rect 24596 50492 24602 50494
rect 24853 50491 24919 50494
rect 30925 50554 30991 50557
rect 31200 50554 32000 50584
rect 30925 50552 32000 50554
rect 30925 50496 30930 50552
rect 30986 50496 32000 50552
rect 30925 50494 32000 50496
rect 30925 50491 30991 50494
rect 31200 50464 32000 50494
rect 20529 50418 20595 50421
rect 20529 50416 22892 50418
rect 20529 50360 20534 50416
rect 20590 50360 22892 50416
rect 20529 50358 22892 50360
rect 20529 50355 20595 50358
rect 22645 50282 22711 50285
rect 22832 50282 22892 50358
rect 23606 50356 23612 50420
rect 23676 50418 23682 50420
rect 23749 50418 23815 50421
rect 23676 50416 23815 50418
rect 23676 50360 23754 50416
rect 23810 50360 23815 50416
rect 23676 50358 23815 50360
rect 23676 50356 23682 50358
rect 23749 50355 23815 50358
rect 25446 50356 25452 50420
rect 25516 50418 25522 50420
rect 28993 50418 29059 50421
rect 25516 50416 29059 50418
rect 25516 50360 28998 50416
rect 29054 50360 29059 50416
rect 25516 50358 29059 50360
rect 25516 50356 25522 50358
rect 28993 50355 29059 50358
rect 29729 50418 29795 50421
rect 30046 50418 30052 50420
rect 29729 50416 30052 50418
rect 29729 50360 29734 50416
rect 29790 50360 30052 50416
rect 29729 50358 30052 50360
rect 29729 50355 29795 50358
rect 30046 50356 30052 50358
rect 30116 50356 30122 50420
rect 25865 50282 25931 50285
rect 22645 50280 22754 50282
rect 22645 50224 22650 50280
rect 22706 50224 22754 50280
rect 22645 50219 22754 50224
rect 22832 50280 25931 50282
rect 22832 50224 25870 50280
rect 25926 50224 25931 50280
rect 22832 50222 25931 50224
rect 25865 50219 25931 50222
rect 30598 50220 30604 50284
rect 30668 50282 30674 50284
rect 31293 50282 31359 50285
rect 30668 50280 31359 50282
rect 30668 50224 31298 50280
rect 31354 50224 31359 50280
rect 30668 50222 31359 50224
rect 30668 50220 30674 50222
rect 31293 50219 31359 50222
rect 10874 50080 11194 50081
rect 10874 50016 10882 50080
rect 10946 50016 10962 50080
rect 11026 50016 11042 50080
rect 11106 50016 11122 50080
rect 11186 50016 11194 50080
rect 10874 50015 11194 50016
rect 20805 50080 21125 50081
rect 20805 50016 20813 50080
rect 20877 50016 20893 50080
rect 20957 50016 20973 50080
rect 21037 50016 21053 50080
rect 21117 50016 21125 50080
rect 20805 50015 21125 50016
rect 22694 50010 22754 50219
rect 27654 50084 27660 50148
rect 27724 50146 27730 50148
rect 29821 50146 29887 50149
rect 27724 50144 29887 50146
rect 27724 50088 29826 50144
rect 29882 50088 29887 50144
rect 27724 50086 29887 50088
rect 27724 50084 27730 50086
rect 29821 50083 29887 50086
rect 22829 50010 22895 50013
rect 22694 50008 22895 50010
rect 22694 49952 22834 50008
rect 22890 49952 22895 50008
rect 22694 49950 22895 49952
rect 22829 49947 22895 49950
rect 23657 50010 23723 50013
rect 23933 50012 23999 50013
rect 24761 50012 24827 50013
rect 23790 50010 23796 50012
rect 23657 50008 23796 50010
rect 23657 49952 23662 50008
rect 23718 49952 23796 50008
rect 23657 49950 23796 49952
rect 23657 49947 23723 49950
rect 23790 49948 23796 49950
rect 23860 49948 23866 50012
rect 23933 50008 23980 50012
rect 24044 50010 24050 50012
rect 23933 49952 23938 50008
rect 23933 49948 23980 49952
rect 24044 49950 24090 50010
rect 24044 49948 24050 49950
rect 24710 49948 24716 50012
rect 24780 50010 24827 50012
rect 25773 50010 25839 50013
rect 26918 50010 26924 50012
rect 24780 50008 24872 50010
rect 24822 49952 24872 50008
rect 24780 49950 24872 49952
rect 25773 50008 26924 50010
rect 25773 49952 25778 50008
rect 25834 49952 26924 50008
rect 25773 49950 26924 49952
rect 24780 49948 24827 49950
rect 23933 49947 23999 49948
rect 24761 49947 24827 49948
rect 25773 49947 25839 49950
rect 26918 49948 26924 49950
rect 26988 49948 26994 50012
rect 29729 50010 29795 50013
rect 31200 50010 32000 50040
rect 29729 50008 32000 50010
rect 29729 49952 29734 50008
rect 29790 49952 32000 50008
rect 29729 49950 32000 49952
rect 29729 49947 29795 49950
rect 31200 49920 32000 49950
rect 0 49874 800 49904
rect 1577 49874 1643 49877
rect 0 49872 1643 49874
rect 0 49816 1582 49872
rect 1638 49816 1643 49872
rect 0 49814 1643 49816
rect 0 49784 800 49814
rect 1577 49811 1643 49814
rect 23013 49874 23079 49877
rect 23238 49874 23244 49876
rect 23013 49872 23244 49874
rect 23013 49816 23018 49872
rect 23074 49816 23244 49872
rect 23013 49814 23244 49816
rect 23013 49811 23079 49814
rect 23238 49812 23244 49814
rect 23308 49812 23314 49876
rect 23381 49874 23447 49877
rect 28717 49874 28783 49877
rect 23381 49872 28783 49874
rect 23381 49816 23386 49872
rect 23442 49816 28722 49872
rect 28778 49816 28783 49872
rect 23381 49814 28783 49816
rect 23381 49811 23447 49814
rect 28717 49811 28783 49814
rect 24342 49676 24348 49740
rect 24412 49738 24418 49740
rect 24945 49738 25011 49741
rect 27429 49738 27495 49741
rect 24412 49736 25011 49738
rect 24412 49680 24950 49736
rect 25006 49680 25011 49736
rect 24412 49678 25011 49680
rect 24412 49676 24418 49678
rect 24945 49675 25011 49678
rect 25224 49736 27495 49738
rect 25224 49680 27434 49736
rect 27490 49680 27495 49736
rect 25224 49678 27495 49680
rect 21909 49602 21975 49605
rect 25224 49602 25284 49678
rect 27429 49675 27495 49678
rect 21909 49600 25284 49602
rect 21909 49544 21914 49600
rect 21970 49544 25284 49600
rect 21909 49542 25284 49544
rect 26877 49602 26943 49605
rect 27981 49602 28047 49605
rect 31200 49602 32000 49632
rect 26877 49600 27906 49602
rect 26877 49544 26882 49600
rect 26938 49544 27906 49600
rect 26877 49542 27906 49544
rect 21909 49539 21975 49542
rect 26877 49539 26943 49542
rect 5909 49536 6229 49537
rect 5909 49472 5917 49536
rect 5981 49472 5997 49536
rect 6061 49472 6077 49536
rect 6141 49472 6157 49536
rect 6221 49472 6229 49536
rect 5909 49471 6229 49472
rect 15840 49536 16160 49537
rect 15840 49472 15848 49536
rect 15912 49472 15928 49536
rect 15992 49472 16008 49536
rect 16072 49472 16088 49536
rect 16152 49472 16160 49536
rect 15840 49471 16160 49472
rect 25770 49536 26090 49537
rect 25770 49472 25778 49536
rect 25842 49472 25858 49536
rect 25922 49472 25938 49536
rect 26002 49472 26018 49536
rect 26082 49472 26090 49536
rect 25770 49471 26090 49472
rect 26969 49468 27035 49469
rect 26918 49466 26924 49468
rect 26878 49406 26924 49466
rect 26988 49464 27035 49468
rect 27429 49468 27495 49469
rect 27429 49466 27476 49468
rect 27030 49408 27035 49464
rect 26918 49404 26924 49406
rect 26988 49404 27035 49408
rect 27384 49464 27476 49466
rect 27384 49408 27434 49464
rect 27384 49406 27476 49408
rect 26969 49403 27035 49404
rect 27429 49404 27476 49406
rect 27540 49404 27546 49468
rect 27429 49403 27495 49404
rect 0 49194 800 49224
rect 2773 49194 2839 49197
rect 0 49192 2839 49194
rect 0 49136 2778 49192
rect 2834 49136 2839 49192
rect 0 49134 2839 49136
rect 0 49104 800 49134
rect 2773 49131 2839 49134
rect 26785 49192 26851 49197
rect 27061 49194 27127 49197
rect 26785 49136 26790 49192
rect 26846 49136 26851 49192
rect 26785 49131 26851 49136
rect 26926 49192 27127 49194
rect 26926 49136 27066 49192
rect 27122 49136 27127 49192
rect 26926 49134 27127 49136
rect 10874 48992 11194 48993
rect 10874 48928 10882 48992
rect 10946 48928 10962 48992
rect 11026 48928 11042 48992
rect 11106 48928 11122 48992
rect 11186 48928 11194 48992
rect 10874 48927 11194 48928
rect 20805 48992 21125 48993
rect 20805 48928 20813 48992
rect 20877 48928 20893 48992
rect 20957 48928 20973 48992
rect 21037 48928 21053 48992
rect 21117 48928 21125 48992
rect 20805 48927 21125 48928
rect 24526 48860 24532 48924
rect 24596 48922 24602 48924
rect 25497 48922 25563 48925
rect 24596 48920 25563 48922
rect 24596 48864 25502 48920
rect 25558 48864 25563 48920
rect 24596 48862 25563 48864
rect 24596 48860 24602 48862
rect 25497 48859 25563 48862
rect 24158 48724 24164 48788
rect 24228 48786 24234 48788
rect 24485 48786 24551 48789
rect 24228 48784 24551 48786
rect 24228 48728 24490 48784
rect 24546 48728 24551 48784
rect 24228 48726 24551 48728
rect 24228 48724 24234 48726
rect 24485 48723 24551 48726
rect 26141 48784 26207 48789
rect 26141 48728 26146 48784
rect 26202 48728 26207 48784
rect 26141 48723 26207 48728
rect 26325 48784 26391 48789
rect 26325 48728 26330 48784
rect 26386 48728 26391 48784
rect 26325 48723 26391 48728
rect 21725 48650 21791 48653
rect 25957 48650 26023 48653
rect 21725 48648 26023 48650
rect 21725 48592 21730 48648
rect 21786 48592 25962 48648
rect 26018 48592 26023 48648
rect 21725 48590 26023 48592
rect 26144 48650 26204 48723
rect 26144 48590 26250 48650
rect 21725 48587 21791 48590
rect 25957 48587 26023 48590
rect 0 48514 800 48544
rect 3417 48514 3483 48517
rect 0 48512 3483 48514
rect 0 48456 3422 48512
rect 3478 48456 3483 48512
rect 0 48454 3483 48456
rect 0 48424 800 48454
rect 3417 48451 3483 48454
rect 24577 48514 24643 48517
rect 24894 48514 24900 48516
rect 24577 48512 24900 48514
rect 24577 48456 24582 48512
rect 24638 48456 24900 48512
rect 24577 48454 24900 48456
rect 24577 48451 24643 48454
rect 24894 48452 24900 48454
rect 24964 48452 24970 48516
rect 5909 48448 6229 48449
rect 5909 48384 5917 48448
rect 5981 48384 5997 48448
rect 6061 48384 6077 48448
rect 6141 48384 6157 48448
rect 6221 48384 6229 48448
rect 5909 48383 6229 48384
rect 15840 48448 16160 48449
rect 15840 48384 15848 48448
rect 15912 48384 15928 48448
rect 15992 48384 16008 48448
rect 16072 48384 16088 48448
rect 16152 48384 16160 48448
rect 15840 48383 16160 48384
rect 25770 48448 26090 48449
rect 25770 48384 25778 48448
rect 25842 48384 25858 48448
rect 25922 48384 25938 48448
rect 26002 48384 26018 48448
rect 26082 48384 26090 48448
rect 25770 48383 26090 48384
rect 26190 48242 26250 48590
rect 26328 48378 26388 48723
rect 26788 48517 26848 49131
rect 26785 48512 26851 48517
rect 26785 48456 26790 48512
rect 26846 48456 26851 48512
rect 26785 48451 26851 48456
rect 26926 48514 26986 49134
rect 27061 49131 27127 49134
rect 27337 49056 27403 49061
rect 27337 49000 27342 49056
rect 27398 49000 27403 49056
rect 27337 48995 27403 49000
rect 27846 49058 27906 49542
rect 27981 49600 32000 49602
rect 27981 49544 27986 49600
rect 28042 49544 32000 49600
rect 27981 49542 32000 49544
rect 27981 49539 28047 49542
rect 31200 49512 32000 49542
rect 29729 49466 29795 49469
rect 30414 49466 30420 49468
rect 29729 49464 30420 49466
rect 29729 49408 29734 49464
rect 29790 49408 30420 49464
rect 29729 49406 30420 49408
rect 29729 49403 29795 49406
rect 30414 49404 30420 49406
rect 30484 49404 30490 49468
rect 30925 49330 30991 49333
rect 31150 49330 31156 49332
rect 30925 49328 31156 49330
rect 30925 49272 30930 49328
rect 30986 49272 31156 49328
rect 30925 49270 31156 49272
rect 30925 49267 30991 49270
rect 31150 49268 31156 49270
rect 31220 49268 31226 49332
rect 28809 49058 28875 49061
rect 31200 49058 32000 49088
rect 27846 48998 28458 49058
rect 27340 48786 27400 48995
rect 27470 48860 27476 48924
rect 27540 48922 27546 48924
rect 28257 48922 28323 48925
rect 27540 48920 28323 48922
rect 27540 48864 28262 48920
rect 28318 48864 28323 48920
rect 27540 48862 28323 48864
rect 27540 48860 27546 48862
rect 28257 48859 28323 48862
rect 27470 48786 27476 48788
rect 27340 48726 27476 48786
rect 27470 48724 27476 48726
rect 27540 48724 27546 48788
rect 27613 48786 27679 48789
rect 28257 48786 28323 48789
rect 28398 48786 28458 48998
rect 28809 49056 32000 49058
rect 28809 49000 28814 49056
rect 28870 49000 32000 49056
rect 28809 48998 32000 49000
rect 28809 48995 28875 48998
rect 31200 48968 32000 48998
rect 27613 48784 28044 48786
rect 27613 48728 27618 48784
rect 27674 48728 28044 48784
rect 27613 48726 28044 48728
rect 27613 48723 27679 48726
rect 27061 48650 27127 48653
rect 27838 48650 27844 48652
rect 27061 48648 27844 48650
rect 27061 48592 27066 48648
rect 27122 48592 27844 48648
rect 27061 48590 27844 48592
rect 27061 48587 27127 48590
rect 27838 48588 27844 48590
rect 27908 48588 27914 48652
rect 27984 48650 28044 48726
rect 28257 48784 28458 48786
rect 28257 48728 28262 48784
rect 28318 48728 28458 48784
rect 28257 48726 28458 48728
rect 28257 48723 28323 48726
rect 28809 48650 28875 48653
rect 31200 48650 32000 48680
rect 27984 48590 28228 48650
rect 27061 48514 27127 48517
rect 26926 48512 27127 48514
rect 26926 48456 27066 48512
rect 27122 48456 27127 48512
rect 26926 48454 27127 48456
rect 27061 48451 27127 48454
rect 27429 48514 27495 48517
rect 28022 48514 28028 48516
rect 27429 48512 28028 48514
rect 27429 48456 27434 48512
rect 27490 48456 28028 48512
rect 27429 48454 28028 48456
rect 27429 48451 27495 48454
rect 28022 48452 28028 48454
rect 28092 48452 28098 48516
rect 26328 48318 26572 48378
rect 26918 48333 26924 48380
rect 26325 48242 26391 48245
rect 26190 48240 26391 48242
rect 26190 48184 26330 48240
rect 26386 48184 26391 48240
rect 26190 48182 26391 48184
rect 26325 48179 26391 48182
rect 20345 48106 20411 48109
rect 25262 48106 25268 48108
rect 20345 48104 25268 48106
rect 20345 48048 20350 48104
rect 20406 48048 25268 48104
rect 20345 48046 25268 48048
rect 20345 48043 20411 48046
rect 25262 48044 25268 48046
rect 25332 48044 25338 48108
rect 26233 48106 26299 48109
rect 26512 48106 26572 48318
rect 26877 48328 26924 48333
rect 26877 48272 26882 48328
rect 26988 48316 26994 48380
rect 28168 48378 28228 48590
rect 28809 48648 32000 48650
rect 28809 48592 28814 48648
rect 28870 48592 32000 48648
rect 28809 48590 32000 48592
rect 28809 48587 28875 48590
rect 31200 48560 32000 48590
rect 28942 48452 28948 48516
rect 29012 48514 29018 48516
rect 29678 48514 29684 48516
rect 29012 48454 29684 48514
rect 29012 48452 29018 48454
rect 29678 48452 29684 48454
rect 29748 48452 29754 48516
rect 27616 48333 28228 48378
rect 27613 48328 28228 48333
rect 26938 48272 26986 48316
rect 26877 48270 26986 48272
rect 27613 48272 27618 48328
rect 27674 48318 28228 48328
rect 27674 48272 27679 48318
rect 28758 48316 28764 48380
rect 28828 48378 28834 48380
rect 28828 48318 29240 48378
rect 28828 48316 28834 48318
rect 26877 48267 26943 48270
rect 27613 48267 27679 48272
rect 28717 48242 28783 48245
rect 28582 48240 28783 48242
rect 28582 48184 28722 48240
rect 28778 48184 28783 48240
rect 28582 48182 28783 48184
rect 29180 48242 29240 48318
rect 29310 48316 29316 48380
rect 29380 48378 29386 48380
rect 29545 48378 29611 48381
rect 29380 48376 29611 48378
rect 29380 48320 29550 48376
rect 29606 48320 29611 48376
rect 29380 48318 29611 48320
rect 29380 48316 29386 48318
rect 29545 48315 29611 48318
rect 30097 48378 30163 48381
rect 31518 48378 31524 48380
rect 30097 48376 31524 48378
rect 30097 48320 30102 48376
rect 30158 48320 31524 48376
rect 30097 48318 31524 48320
rect 30097 48315 30163 48318
rect 31518 48316 31524 48318
rect 31588 48316 31594 48380
rect 29545 48242 29611 48245
rect 29180 48240 29611 48242
rect 29180 48184 29550 48240
rect 29606 48184 29611 48240
rect 29180 48182 29611 48184
rect 26233 48104 26572 48106
rect 26233 48048 26238 48104
rect 26294 48048 26572 48104
rect 26233 48046 26572 48048
rect 27245 48108 27311 48109
rect 27245 48104 27292 48108
rect 27356 48106 27362 48108
rect 27245 48048 27250 48104
rect 26233 48043 26299 48046
rect 27245 48044 27292 48048
rect 27356 48046 27402 48106
rect 27356 48044 27362 48046
rect 27245 48043 27311 48044
rect 27337 47970 27403 47973
rect 27470 47970 27476 47972
rect 27337 47968 27476 47970
rect 27337 47912 27342 47968
rect 27398 47912 27476 47968
rect 27337 47910 27476 47912
rect 27337 47907 27403 47910
rect 27470 47908 27476 47910
rect 27540 47908 27546 47972
rect 10874 47904 11194 47905
rect 0 47834 800 47864
rect 10874 47840 10882 47904
rect 10946 47840 10962 47904
rect 11026 47840 11042 47904
rect 11106 47840 11122 47904
rect 11186 47840 11194 47904
rect 10874 47839 11194 47840
rect 20805 47904 21125 47905
rect 20805 47840 20813 47904
rect 20877 47840 20893 47904
rect 20957 47840 20973 47904
rect 21037 47840 21053 47904
rect 21117 47840 21125 47904
rect 20805 47839 21125 47840
rect 2221 47834 2287 47837
rect 0 47832 2287 47834
rect 0 47776 2226 47832
rect 2282 47776 2287 47832
rect 0 47774 2287 47776
rect 0 47744 800 47774
rect 2221 47771 2287 47774
rect 16849 47834 16915 47837
rect 17861 47834 17927 47837
rect 16849 47832 17927 47834
rect 16849 47776 16854 47832
rect 16910 47776 17866 47832
rect 17922 47776 17927 47832
rect 16849 47774 17927 47776
rect 16849 47771 16915 47774
rect 17861 47771 17927 47774
rect 25957 47834 26023 47837
rect 26182 47834 26188 47836
rect 25957 47832 26188 47834
rect 25957 47776 25962 47832
rect 26018 47776 26188 47832
rect 25957 47774 26188 47776
rect 25957 47771 26023 47774
rect 26182 47772 26188 47774
rect 26252 47772 26258 47836
rect 28582 47698 28642 48182
rect 28717 48179 28783 48182
rect 29545 48179 29611 48182
rect 28717 48106 28783 48109
rect 31200 48106 32000 48136
rect 28717 48104 32000 48106
rect 28717 48048 28722 48104
rect 28778 48048 32000 48104
rect 28717 48046 32000 48048
rect 28717 48043 28783 48046
rect 31200 48016 32000 48046
rect 28758 47908 28764 47972
rect 28828 47970 28834 47972
rect 28993 47970 29059 47973
rect 28828 47968 29059 47970
rect 28828 47912 28998 47968
rect 29054 47912 29059 47968
rect 28828 47910 29059 47912
rect 28828 47908 28834 47910
rect 28993 47907 29059 47910
rect 31200 47698 32000 47728
rect 28582 47638 32000 47698
rect 31200 47608 32000 47638
rect 30046 47364 30052 47428
rect 30116 47426 30122 47428
rect 31886 47426 31892 47428
rect 30116 47366 31892 47426
rect 30116 47364 30122 47366
rect 31886 47364 31892 47366
rect 31956 47364 31962 47428
rect 5909 47360 6229 47361
rect 0 47290 800 47320
rect 5909 47296 5917 47360
rect 5981 47296 5997 47360
rect 6061 47296 6077 47360
rect 6141 47296 6157 47360
rect 6221 47296 6229 47360
rect 5909 47295 6229 47296
rect 15840 47360 16160 47361
rect 15840 47296 15848 47360
rect 15912 47296 15928 47360
rect 15992 47296 16008 47360
rect 16072 47296 16088 47360
rect 16152 47296 16160 47360
rect 15840 47295 16160 47296
rect 25770 47360 26090 47361
rect 25770 47296 25778 47360
rect 25842 47296 25858 47360
rect 25922 47296 25938 47360
rect 26002 47296 26018 47360
rect 26082 47296 26090 47360
rect 25770 47295 26090 47296
rect 1577 47290 1643 47293
rect 0 47288 1643 47290
rect 0 47232 1582 47288
rect 1638 47232 1643 47288
rect 0 47230 1643 47232
rect 0 47200 800 47230
rect 1577 47227 1643 47230
rect 30782 47228 30788 47292
rect 30852 47290 30858 47292
rect 30925 47290 30991 47293
rect 30852 47288 30991 47290
rect 30852 47232 30930 47288
rect 30986 47232 30991 47288
rect 30852 47230 30991 47232
rect 30852 47228 30858 47230
rect 30925 47227 30991 47230
rect 17309 47154 17375 47157
rect 19149 47154 19215 47157
rect 17309 47152 19215 47154
rect 17309 47096 17314 47152
rect 17370 47096 19154 47152
rect 19210 47096 19215 47152
rect 17309 47094 19215 47096
rect 17309 47091 17375 47094
rect 19149 47091 19215 47094
rect 29729 47154 29795 47157
rect 31200 47154 32000 47184
rect 29729 47152 32000 47154
rect 29729 47096 29734 47152
rect 29790 47096 32000 47152
rect 29729 47094 32000 47096
rect 29729 47091 29795 47094
rect 31200 47064 32000 47094
rect 26366 46820 26372 46884
rect 26436 46882 26442 46884
rect 26509 46882 26575 46885
rect 26436 46880 26575 46882
rect 26436 46824 26514 46880
rect 26570 46824 26575 46880
rect 26436 46822 26575 46824
rect 26436 46820 26442 46822
rect 26509 46819 26575 46822
rect 10874 46816 11194 46817
rect 10874 46752 10882 46816
rect 10946 46752 10962 46816
rect 11026 46752 11042 46816
rect 11106 46752 11122 46816
rect 11186 46752 11194 46816
rect 10874 46751 11194 46752
rect 20805 46816 21125 46817
rect 20805 46752 20813 46816
rect 20877 46752 20893 46816
rect 20957 46752 20973 46816
rect 21037 46752 21053 46816
rect 21117 46752 21125 46816
rect 20805 46751 21125 46752
rect 25262 46684 25268 46748
rect 25332 46684 25338 46748
rect 29729 46746 29795 46749
rect 31200 46746 32000 46776
rect 29729 46744 32000 46746
rect 29729 46688 29734 46744
rect 29790 46688 32000 46744
rect 29729 46686 32000 46688
rect 0 46610 800 46640
rect 1577 46610 1643 46613
rect 0 46608 1643 46610
rect 0 46552 1582 46608
rect 1638 46552 1643 46608
rect 0 46550 1643 46552
rect 0 46520 800 46550
rect 1577 46547 1643 46550
rect 22185 46474 22251 46477
rect 23238 46474 23244 46476
rect 22185 46472 23244 46474
rect 22185 46416 22190 46472
rect 22246 46416 23244 46472
rect 22185 46414 23244 46416
rect 22185 46411 22251 46414
rect 23238 46412 23244 46414
rect 23308 46412 23314 46476
rect 24894 46412 24900 46476
rect 24964 46474 24970 46476
rect 25270 46474 25330 46684
rect 29729 46683 29795 46686
rect 31200 46656 32000 46686
rect 25497 46474 25563 46477
rect 24964 46472 25563 46474
rect 24964 46416 25502 46472
rect 25558 46416 25563 46472
rect 24964 46414 25563 46416
rect 24964 46412 24970 46414
rect 25497 46411 25563 46414
rect 25773 46474 25839 46477
rect 26182 46474 26188 46476
rect 25773 46472 26188 46474
rect 25773 46416 25778 46472
rect 25834 46416 26188 46472
rect 25773 46414 26188 46416
rect 25773 46411 25839 46414
rect 26182 46412 26188 46414
rect 26252 46412 26258 46476
rect 30598 46412 30604 46476
rect 30668 46474 30674 46476
rect 31109 46474 31175 46477
rect 30668 46472 31175 46474
rect 30668 46416 31114 46472
rect 31170 46416 31175 46472
rect 30668 46414 31175 46416
rect 30668 46412 30674 46414
rect 31109 46411 31175 46414
rect 31385 46474 31451 46477
rect 31518 46474 31524 46476
rect 31385 46472 31524 46474
rect 31385 46416 31390 46472
rect 31446 46416 31524 46472
rect 31385 46414 31524 46416
rect 31385 46411 31451 46414
rect 31518 46412 31524 46414
rect 31588 46412 31594 46476
rect 5909 46272 6229 46273
rect 5909 46208 5917 46272
rect 5981 46208 5997 46272
rect 6061 46208 6077 46272
rect 6141 46208 6157 46272
rect 6221 46208 6229 46272
rect 5909 46207 6229 46208
rect 15840 46272 16160 46273
rect 15840 46208 15848 46272
rect 15912 46208 15928 46272
rect 15992 46208 16008 46272
rect 16072 46208 16088 46272
rect 16152 46208 16160 46272
rect 15840 46207 16160 46208
rect 25770 46272 26090 46273
rect 25770 46208 25778 46272
rect 25842 46208 25858 46272
rect 25922 46208 25938 46272
rect 26002 46208 26018 46272
rect 26082 46208 26090 46272
rect 25770 46207 26090 46208
rect 25078 46140 25084 46204
rect 25148 46202 25154 46204
rect 25221 46202 25287 46205
rect 25148 46200 25287 46202
rect 25148 46144 25226 46200
rect 25282 46144 25287 46200
rect 25148 46142 25287 46144
rect 25148 46140 25154 46142
rect 25221 46139 25287 46142
rect 27838 46140 27844 46204
rect 27908 46202 27914 46204
rect 28942 46202 28948 46204
rect 27908 46142 28948 46202
rect 27908 46140 27914 46142
rect 28942 46140 28948 46142
rect 29012 46140 29018 46204
rect 29729 46202 29795 46205
rect 31200 46202 32000 46232
rect 29729 46200 32000 46202
rect 29729 46144 29734 46200
rect 29790 46144 32000 46200
rect 29729 46142 32000 46144
rect 29729 46139 29795 46142
rect 31200 46112 32000 46142
rect 29729 46066 29795 46069
rect 30230 46066 30236 46068
rect 29729 46064 30236 46066
rect 29729 46008 29734 46064
rect 29790 46008 30236 46064
rect 29729 46006 30236 46008
rect 29729 46003 29795 46006
rect 30230 46004 30236 46006
rect 30300 46004 30306 46068
rect 0 45930 800 45960
rect 1393 45930 1459 45933
rect 0 45928 1459 45930
rect 0 45872 1398 45928
rect 1454 45872 1459 45928
rect 0 45870 1459 45872
rect 0 45840 800 45870
rect 1393 45867 1459 45870
rect 28206 45868 28212 45932
rect 28276 45930 28282 45932
rect 28901 45930 28967 45933
rect 28276 45928 28967 45930
rect 28276 45872 28906 45928
rect 28962 45872 28967 45928
rect 28276 45870 28967 45872
rect 28276 45868 28282 45870
rect 28901 45867 28967 45870
rect 10874 45728 11194 45729
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 45663 11194 45664
rect 20805 45728 21125 45729
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 31200 45704 32000 45824
rect 20805 45663 21125 45664
rect 28942 45596 28948 45660
rect 29012 45658 29018 45660
rect 29085 45658 29151 45661
rect 29637 45658 29703 45661
rect 29012 45656 29151 45658
rect 29012 45600 29090 45656
rect 29146 45600 29151 45656
rect 29012 45598 29151 45600
rect 29012 45596 29018 45598
rect 29085 45595 29151 45598
rect 29318 45656 29703 45658
rect 29318 45600 29642 45656
rect 29698 45600 29703 45656
rect 29318 45598 29703 45600
rect 26918 45460 26924 45524
rect 26988 45522 26994 45524
rect 28533 45522 28599 45525
rect 26988 45520 28599 45522
rect 26988 45464 28538 45520
rect 28594 45464 28599 45520
rect 26988 45462 28599 45464
rect 26988 45460 26994 45462
rect 28533 45459 28599 45462
rect 29085 45522 29151 45525
rect 29318 45522 29378 45598
rect 29637 45595 29703 45598
rect 29085 45520 29378 45522
rect 29085 45464 29090 45520
rect 29146 45464 29378 45520
rect 29085 45462 29378 45464
rect 29085 45459 29151 45462
rect 31200 45296 32000 45416
rect 0 45250 800 45280
rect 1485 45250 1551 45253
rect 0 45248 1551 45250
rect 0 45192 1490 45248
rect 1546 45192 1551 45248
rect 0 45190 1551 45192
rect 0 45160 800 45190
rect 1485 45187 1551 45190
rect 5909 45184 6229 45185
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6229 45184
rect 5909 45119 6229 45120
rect 15840 45184 16160 45185
rect 15840 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15840 45119 16160 45120
rect 25770 45184 26090 45185
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26090 45184
rect 25770 45119 26090 45120
rect 24342 45052 24348 45116
rect 24412 45114 24418 45116
rect 24669 45114 24735 45117
rect 24412 45112 24735 45114
rect 24412 45056 24674 45112
rect 24730 45056 24735 45112
rect 24412 45054 24735 45056
rect 24412 45052 24418 45054
rect 24669 45051 24735 45054
rect 26325 45116 26391 45117
rect 26325 45112 26372 45116
rect 26436 45114 26442 45116
rect 26325 45056 26330 45112
rect 26325 45052 26372 45056
rect 26436 45054 26482 45114
rect 26436 45052 26442 45054
rect 31518 45052 31524 45116
rect 31588 45114 31594 45116
rect 31845 45114 31911 45117
rect 31588 45112 31911 45114
rect 31588 45056 31850 45112
rect 31906 45056 31911 45112
rect 31588 45054 31911 45056
rect 31588 45052 31594 45054
rect 26325 45051 26391 45052
rect 31845 45051 31911 45054
rect 28809 44842 28875 44845
rect 31200 44842 32000 44872
rect 28809 44840 32000 44842
rect 28809 44784 28814 44840
rect 28870 44784 32000 44840
rect 28809 44782 32000 44784
rect 28809 44779 28875 44782
rect 31200 44752 32000 44782
rect 27470 44644 27476 44708
rect 27540 44706 27546 44708
rect 27797 44706 27863 44709
rect 27540 44704 27863 44706
rect 27540 44648 27802 44704
rect 27858 44648 27863 44704
rect 27540 44646 27863 44648
rect 27540 44644 27546 44646
rect 27797 44643 27863 44646
rect 10874 44640 11194 44641
rect 0 44570 800 44600
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 44575 11194 44576
rect 20805 44640 21125 44641
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 44575 21125 44576
rect 1577 44570 1643 44573
rect 0 44568 1643 44570
rect 0 44512 1582 44568
rect 1638 44512 1643 44568
rect 0 44510 1643 44512
rect 0 44480 800 44510
rect 1577 44507 1643 44510
rect 27286 44508 27292 44572
rect 27356 44570 27362 44572
rect 27981 44570 28047 44573
rect 28758 44570 28764 44572
rect 27356 44568 28047 44570
rect 27356 44512 27986 44568
rect 28042 44512 28047 44568
rect 27356 44510 28047 44512
rect 27356 44508 27362 44510
rect 27981 44507 28047 44510
rect 28582 44510 28764 44570
rect 12341 44434 12407 44437
rect 12893 44434 12959 44437
rect 12341 44432 12959 44434
rect 12341 44376 12346 44432
rect 12402 44376 12898 44432
rect 12954 44376 12959 44432
rect 12341 44374 12959 44376
rect 12341 44371 12407 44374
rect 12893 44371 12959 44374
rect 27429 44434 27495 44437
rect 27654 44434 27660 44436
rect 27429 44432 27660 44434
rect 27429 44376 27434 44432
rect 27490 44376 27660 44432
rect 27429 44374 27660 44376
rect 27429 44371 27495 44374
rect 27654 44372 27660 44374
rect 27724 44372 27730 44436
rect 11605 44298 11671 44301
rect 18597 44298 18663 44301
rect 11605 44296 18663 44298
rect 11605 44240 11610 44296
rect 11666 44240 18602 44296
rect 18658 44240 18663 44296
rect 11605 44238 18663 44240
rect 11605 44235 11671 44238
rect 18597 44235 18663 44238
rect 28582 44162 28642 44510
rect 28758 44508 28764 44510
rect 28828 44508 28834 44572
rect 30005 44570 30071 44573
rect 30230 44570 30236 44572
rect 30005 44568 30236 44570
rect 30005 44512 30010 44568
rect 30066 44512 30236 44568
rect 30005 44510 30236 44512
rect 30005 44507 30071 44510
rect 30230 44508 30236 44510
rect 30300 44508 30306 44572
rect 28717 44434 28783 44437
rect 31200 44434 32000 44464
rect 28717 44432 32000 44434
rect 28717 44376 28722 44432
rect 28778 44376 32000 44432
rect 28717 44374 32000 44376
rect 28717 44371 28783 44374
rect 31200 44344 32000 44374
rect 28758 44236 28764 44300
rect 28828 44298 28834 44300
rect 28901 44298 28967 44301
rect 28828 44296 28967 44298
rect 28828 44240 28906 44296
rect 28962 44240 28967 44296
rect 28828 44238 28967 44240
rect 28828 44236 28834 44238
rect 28901 44235 28967 44238
rect 29678 44236 29684 44300
rect 29748 44298 29754 44300
rect 30005 44298 30071 44301
rect 29748 44296 30071 44298
rect 29748 44240 30010 44296
rect 30066 44240 30071 44296
rect 29748 44238 30071 44240
rect 29748 44236 29754 44238
rect 30005 44235 30071 44238
rect 28901 44162 28967 44165
rect 28582 44160 28967 44162
rect 28582 44104 28906 44160
rect 28962 44104 28967 44160
rect 28582 44102 28967 44104
rect 28901 44099 28967 44102
rect 30649 44162 30715 44165
rect 31702 44162 31708 44164
rect 30649 44160 31708 44162
rect 30649 44104 30654 44160
rect 30710 44104 31708 44160
rect 30649 44102 31708 44104
rect 30649 44099 30715 44102
rect 31702 44100 31708 44102
rect 31772 44100 31778 44164
rect 5909 44096 6229 44097
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6229 44096
rect 5909 44031 6229 44032
rect 15840 44096 16160 44097
rect 15840 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15840 44031 16160 44032
rect 25770 44096 26090 44097
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26090 44096
rect 25770 44031 26090 44032
rect 24485 44024 24551 44029
rect 24485 43968 24490 44024
rect 24546 43968 24551 44024
rect 24485 43963 24551 43968
rect 0 43890 800 43920
rect 2773 43890 2839 43893
rect 0 43888 2839 43890
rect 0 43832 2778 43888
rect 2834 43832 2839 43888
rect 0 43830 2839 43832
rect 0 43800 800 43830
rect 2773 43827 2839 43830
rect 9397 43754 9463 43757
rect 13077 43754 13143 43757
rect 9397 43752 13143 43754
rect 9397 43696 9402 43752
rect 9458 43696 13082 43752
rect 13138 43696 13143 43752
rect 9397 43694 13143 43696
rect 9397 43691 9463 43694
rect 13077 43691 13143 43694
rect 23749 43754 23815 43757
rect 24301 43754 24367 43757
rect 24488 43754 24548 43963
rect 29821 43890 29887 43893
rect 31200 43890 32000 43920
rect 29821 43888 32000 43890
rect 29821 43832 29826 43888
rect 29882 43832 32000 43888
rect 29821 43830 32000 43832
rect 29821 43827 29887 43830
rect 31200 43800 32000 43830
rect 23749 43752 24548 43754
rect 23749 43696 23754 43752
rect 23810 43696 24306 43752
rect 24362 43696 24548 43752
rect 23749 43694 24548 43696
rect 23749 43691 23815 43694
rect 24301 43691 24367 43694
rect 29913 43618 29979 43621
rect 30966 43618 30972 43620
rect 29913 43616 30972 43618
rect 29913 43560 29918 43616
rect 29974 43560 30972 43616
rect 29913 43558 30972 43560
rect 29913 43555 29979 43558
rect 30966 43556 30972 43558
rect 31036 43556 31042 43620
rect 10874 43552 11194 43553
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 43487 11194 43488
rect 20805 43552 21125 43553
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 43487 21125 43488
rect 29821 43482 29887 43485
rect 31200 43482 32000 43512
rect 29821 43480 32000 43482
rect 29821 43424 29826 43480
rect 29882 43424 32000 43480
rect 29821 43422 32000 43424
rect 29821 43419 29887 43422
rect 31200 43392 32000 43422
rect 21398 43284 21404 43348
rect 21468 43346 21474 43348
rect 22001 43346 22067 43349
rect 28993 43346 29059 43349
rect 21468 43344 22067 43346
rect 21468 43288 22006 43344
rect 22062 43288 22067 43344
rect 21468 43286 22067 43288
rect 21468 43284 21474 43286
rect 22001 43283 22067 43286
rect 28950 43344 29059 43346
rect 28950 43288 28998 43344
rect 29054 43288 29059 43344
rect 28950 43283 29059 43288
rect 29361 43346 29427 43349
rect 29361 43344 30298 43346
rect 29361 43288 29366 43344
rect 29422 43288 30298 43344
rect 29361 43286 30298 43288
rect 29361 43283 29427 43286
rect 0 43210 800 43240
rect 2221 43210 2287 43213
rect 0 43208 2287 43210
rect 0 43152 2226 43208
rect 2282 43152 2287 43208
rect 0 43150 2287 43152
rect 0 43120 800 43150
rect 2221 43147 2287 43150
rect 23289 43208 23355 43213
rect 24025 43212 24091 43213
rect 24761 43212 24827 43213
rect 23289 43152 23294 43208
rect 23350 43152 23355 43208
rect 23289 43147 23355 43152
rect 23974 43148 23980 43212
rect 24044 43210 24091 43212
rect 24710 43210 24716 43212
rect 24044 43208 24136 43210
rect 24086 43152 24136 43208
rect 24044 43150 24136 43152
rect 24670 43150 24716 43210
rect 24780 43208 24827 43212
rect 24822 43152 24827 43208
rect 24044 43148 24091 43150
rect 24710 43148 24716 43150
rect 24780 43148 24827 43152
rect 27654 43148 27660 43212
rect 27724 43210 27730 43212
rect 27981 43210 28047 43213
rect 27724 43208 28047 43210
rect 27724 43152 27986 43208
rect 28042 43152 28047 43208
rect 27724 43150 28047 43152
rect 27724 43148 27730 43150
rect 24025 43147 24091 43148
rect 24761 43147 24827 43148
rect 27981 43147 28047 43150
rect 23292 43074 23352 43147
rect 24025 43074 24091 43077
rect 23292 43072 24091 43074
rect 23292 43016 24030 43072
rect 24086 43016 24091 43072
rect 23292 43014 24091 43016
rect 24025 43011 24091 43014
rect 24485 43074 24551 43077
rect 25129 43074 25195 43077
rect 24485 43072 25195 43074
rect 24485 43016 24490 43072
rect 24546 43016 25134 43072
rect 25190 43016 25195 43072
rect 24485 43014 25195 43016
rect 24485 43011 24551 43014
rect 25129 43011 25195 43014
rect 5909 43008 6229 43009
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6229 43008
rect 5909 42943 6229 42944
rect 15840 43008 16160 43009
rect 15840 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15840 42943 16160 42944
rect 25770 43008 26090 43009
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26090 43008
rect 25770 42943 26090 42944
rect 24761 42938 24827 42941
rect 25262 42938 25268 42940
rect 24761 42936 25268 42938
rect 24761 42880 24766 42936
rect 24822 42880 25268 42936
rect 24761 42878 25268 42880
rect 24761 42875 24827 42878
rect 25262 42876 25268 42878
rect 25332 42876 25338 42940
rect 25865 42802 25931 42805
rect 26182 42802 26188 42804
rect 25865 42800 26188 42802
rect 25865 42744 25870 42800
rect 25926 42744 26188 42800
rect 25865 42742 26188 42744
rect 25865 42739 25931 42742
rect 26182 42740 26188 42742
rect 26252 42740 26258 42804
rect 0 42666 800 42696
rect 1577 42666 1643 42669
rect 0 42664 1643 42666
rect 0 42608 1582 42664
rect 1638 42608 1643 42664
rect 0 42606 1643 42608
rect 0 42576 800 42606
rect 1577 42603 1643 42606
rect 24669 42666 24735 42669
rect 24853 42666 24919 42669
rect 24669 42664 24919 42666
rect 24669 42608 24674 42664
rect 24730 42608 24858 42664
rect 24914 42608 24919 42664
rect 24669 42606 24919 42608
rect 24669 42603 24735 42606
rect 24853 42603 24919 42606
rect 25262 42604 25268 42668
rect 25332 42666 25338 42668
rect 27102 42666 27108 42668
rect 25332 42606 27108 42666
rect 25332 42604 25338 42606
rect 27102 42604 27108 42606
rect 27172 42604 27178 42668
rect 27705 42666 27771 42669
rect 27705 42664 28228 42666
rect 27705 42608 27710 42664
rect 27766 42608 28228 42664
rect 27705 42606 28228 42608
rect 27705 42603 27771 42606
rect 22277 42530 22343 42533
rect 25773 42530 25839 42533
rect 22277 42528 25839 42530
rect 22277 42472 22282 42528
rect 22338 42472 25778 42528
rect 25834 42472 25839 42528
rect 22277 42470 25839 42472
rect 22277 42467 22343 42470
rect 25773 42467 25839 42470
rect 10874 42464 11194 42465
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 42399 11194 42400
rect 20805 42464 21125 42465
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 20805 42399 21125 42400
rect 23289 42396 23355 42397
rect 23238 42332 23244 42396
rect 23308 42394 23355 42396
rect 25313 42394 25379 42397
rect 26182 42394 26188 42396
rect 23308 42392 23400 42394
rect 23350 42336 23400 42392
rect 23308 42334 23400 42336
rect 25313 42392 26188 42394
rect 25313 42336 25318 42392
rect 25374 42336 26188 42392
rect 25313 42334 26188 42336
rect 23308 42332 23355 42334
rect 23289 42331 23355 42332
rect 25313 42331 25379 42334
rect 26182 42332 26188 42334
rect 26252 42332 26258 42396
rect 27429 42394 27495 42397
rect 26742 42392 27495 42394
rect 26742 42336 27434 42392
rect 27490 42336 27495 42392
rect 26742 42334 27495 42336
rect 24025 42258 24091 42261
rect 24710 42258 24716 42260
rect 24025 42256 24716 42258
rect 24025 42200 24030 42256
rect 24086 42200 24716 42256
rect 24025 42198 24716 42200
rect 24025 42195 24091 42198
rect 24710 42196 24716 42198
rect 24780 42258 24786 42260
rect 25865 42258 25931 42261
rect 24780 42256 25931 42258
rect 24780 42200 25870 42256
rect 25926 42200 25931 42256
rect 24780 42198 25931 42200
rect 24780 42196 24786 42198
rect 25865 42195 25931 42198
rect 0 41986 800 42016
rect 26742 41989 26802 42334
rect 27429 42331 27495 42334
rect 27613 42256 27679 42261
rect 27613 42200 27618 42256
rect 27674 42200 27679 42256
rect 27613 42195 27679 42200
rect 1577 41986 1643 41989
rect 0 41984 1643 41986
rect 0 41928 1582 41984
rect 1638 41928 1643 41984
rect 0 41926 1643 41928
rect 0 41896 800 41926
rect 1577 41923 1643 41926
rect 26693 41984 26802 41989
rect 26693 41928 26698 41984
rect 26754 41928 26802 41984
rect 26693 41926 26802 41928
rect 26693 41923 26759 41926
rect 5909 41920 6229 41921
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6229 41920
rect 5909 41855 6229 41856
rect 15840 41920 16160 41921
rect 15840 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15840 41855 16160 41856
rect 25770 41920 26090 41921
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26090 41920
rect 25770 41855 26090 41856
rect 27616 41850 27676 42195
rect 27797 41986 27863 41989
rect 28168 41986 28228 42606
rect 27797 41984 28228 41986
rect 27797 41928 27802 41984
rect 27858 41928 28228 41984
rect 27797 41926 28228 41928
rect 28950 41986 29010 43283
rect 29269 43210 29335 43213
rect 29134 43208 29335 43210
rect 29134 43152 29274 43208
rect 29330 43152 29335 43208
rect 29134 43150 29335 43152
rect 29134 42666 29194 43150
rect 29269 43147 29335 43150
rect 29862 43012 29868 43076
rect 29932 43074 29938 43076
rect 30046 43074 30052 43076
rect 29932 43014 30052 43074
rect 29932 43012 29938 43014
rect 30046 43012 30052 43014
rect 30116 43012 30122 43076
rect 30238 43074 30298 43286
rect 30414 43284 30420 43348
rect 30484 43346 30490 43348
rect 30649 43346 30715 43349
rect 30484 43344 30715 43346
rect 30484 43288 30654 43344
rect 30710 43288 30715 43344
rect 30484 43286 30715 43288
rect 30484 43284 30490 43286
rect 30649 43283 30715 43286
rect 30782 43148 30788 43212
rect 30852 43210 30858 43212
rect 31334 43210 31340 43212
rect 30852 43150 31340 43210
rect 30852 43148 30858 43150
rect 31334 43148 31340 43150
rect 31404 43148 31410 43212
rect 30414 43074 30420 43076
rect 30238 43014 30420 43074
rect 30414 43012 30420 43014
rect 30484 43012 30490 43076
rect 29269 42938 29335 42941
rect 31200 42938 32000 42968
rect 29269 42936 32000 42938
rect 29269 42880 29274 42936
rect 29330 42880 32000 42936
rect 29269 42878 32000 42880
rect 29269 42875 29335 42878
rect 31200 42848 32000 42878
rect 29862 42740 29868 42804
rect 29932 42802 29938 42804
rect 30005 42802 30071 42805
rect 29932 42800 30071 42802
rect 29932 42744 30010 42800
rect 30066 42744 30071 42800
rect 29932 42742 30071 42744
rect 29932 42740 29938 42742
rect 30005 42739 30071 42742
rect 29361 42666 29427 42669
rect 29134 42664 29427 42666
rect 29134 42608 29366 42664
rect 29422 42608 29427 42664
rect 29134 42606 29427 42608
rect 29361 42603 29427 42606
rect 29637 42666 29703 42669
rect 30966 42666 30972 42668
rect 29637 42664 30972 42666
rect 29637 42608 29642 42664
rect 29698 42608 30972 42664
rect 29637 42606 30972 42608
rect 29637 42603 29703 42606
rect 30966 42604 30972 42606
rect 31036 42604 31042 42668
rect 29913 42530 29979 42533
rect 31200 42530 32000 42560
rect 29913 42528 32000 42530
rect 29913 42472 29918 42528
rect 29974 42472 32000 42528
rect 29913 42470 32000 42472
rect 29913 42467 29979 42470
rect 31200 42440 32000 42470
rect 29126 42332 29132 42396
rect 29196 42394 29202 42396
rect 29545 42394 29611 42397
rect 29196 42392 29611 42394
rect 29196 42336 29550 42392
rect 29606 42336 29611 42392
rect 29196 42334 29611 42336
rect 29196 42332 29202 42334
rect 29545 42331 29611 42334
rect 29177 42260 29243 42261
rect 29126 42196 29132 42260
rect 29196 42258 29243 42260
rect 29729 42258 29795 42261
rect 30557 42258 30623 42261
rect 29196 42256 29288 42258
rect 29238 42200 29288 42256
rect 29196 42198 29288 42200
rect 29729 42256 30623 42258
rect 29729 42200 29734 42256
rect 29790 42200 30562 42256
rect 30618 42200 30623 42256
rect 29729 42198 30623 42200
rect 29196 42196 29243 42198
rect 29177 42195 29243 42196
rect 29729 42195 29795 42198
rect 30557 42195 30623 42198
rect 29453 42120 29519 42125
rect 29453 42064 29458 42120
rect 29514 42064 29519 42120
rect 29453 42059 29519 42064
rect 30005 42120 30071 42125
rect 30005 42064 30010 42120
rect 30066 42064 30071 42120
rect 30005 42059 30071 42064
rect 29085 41986 29151 41989
rect 28950 41984 29151 41986
rect 28950 41928 29090 41984
rect 29146 41928 29151 41984
rect 28950 41926 29151 41928
rect 27797 41923 27863 41926
rect 29085 41923 29151 41926
rect 29456 41850 29516 42059
rect 30008 41986 30068 42059
rect 31200 41986 32000 42016
rect 30008 41926 32000 41986
rect 31200 41896 32000 41926
rect 22326 41790 23536 41850
rect 27616 41790 27722 41850
rect 29456 41790 31034 41850
rect 22093 41714 22159 41717
rect 22326 41714 22386 41790
rect 22093 41712 22386 41714
rect 22093 41656 22098 41712
rect 22154 41656 22386 41712
rect 22093 41654 22386 41656
rect 23013 41712 23079 41717
rect 23013 41656 23018 41712
rect 23074 41656 23079 41712
rect 22093 41651 22159 41654
rect 23013 41651 23079 41656
rect 23476 41714 23536 41790
rect 27521 41714 27587 41717
rect 23476 41654 26572 41714
rect 10874 41376 11194 41377
rect 0 41306 800 41336
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 41311 11194 41312
rect 20805 41376 21125 41377
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 41311 21125 41312
rect 1577 41306 1643 41309
rect 0 41304 1643 41306
rect 0 41248 1582 41304
rect 1638 41248 1643 41304
rect 0 41246 1643 41248
rect 23016 41306 23076 41651
rect 23473 41578 23539 41581
rect 25313 41580 25379 41581
rect 24158 41578 24164 41580
rect 23473 41576 24164 41578
rect 23473 41520 23478 41576
rect 23534 41520 24164 41576
rect 23473 41518 24164 41520
rect 23473 41515 23539 41518
rect 24158 41516 24164 41518
rect 24228 41516 24234 41580
rect 25262 41516 25268 41580
rect 25332 41578 25379 41580
rect 25681 41578 25747 41581
rect 26366 41578 26372 41580
rect 25332 41576 25424 41578
rect 25374 41520 25424 41576
rect 25332 41518 25424 41520
rect 25681 41576 26372 41578
rect 25681 41520 25686 41576
rect 25742 41520 26372 41576
rect 25681 41518 26372 41520
rect 25332 41516 25379 41518
rect 25313 41515 25379 41516
rect 25681 41515 25747 41518
rect 26366 41516 26372 41518
rect 26436 41516 26442 41580
rect 26512 41445 26572 41654
rect 27294 41712 27587 41714
rect 27294 41656 27526 41712
rect 27582 41656 27587 41712
rect 27294 41654 27587 41656
rect 26877 41580 26943 41581
rect 26877 41578 26924 41580
rect 26832 41576 26924 41578
rect 26832 41520 26882 41576
rect 26832 41518 26924 41520
rect 26877 41516 26924 41518
rect 26988 41516 26994 41580
rect 26877 41515 26943 41516
rect 24342 41380 24348 41444
rect 24412 41442 24418 41444
rect 25497 41442 25563 41445
rect 24412 41440 25563 41442
rect 24412 41384 25502 41440
rect 25558 41384 25563 41440
rect 24412 41382 25563 41384
rect 24412 41380 24418 41382
rect 25497 41379 25563 41382
rect 26141 41442 26207 41445
rect 26366 41442 26372 41444
rect 26141 41440 26372 41442
rect 26141 41384 26146 41440
rect 26202 41384 26372 41440
rect 26141 41382 26372 41384
rect 26141 41379 26207 41382
rect 26366 41380 26372 41382
rect 26436 41380 26442 41444
rect 26509 41442 26575 41445
rect 26734 41442 26740 41444
rect 26509 41440 26740 41442
rect 26509 41384 26514 41440
rect 26570 41384 26740 41440
rect 26509 41382 26740 41384
rect 26509 41379 26575 41382
rect 26734 41380 26740 41382
rect 26804 41380 26810 41444
rect 24301 41306 24367 41309
rect 23016 41304 24367 41306
rect 23016 41248 24306 41304
rect 24362 41248 24367 41304
rect 23016 41246 24367 41248
rect 0 41216 800 41246
rect 1577 41243 1643 41246
rect 24301 41243 24367 41246
rect 24761 41306 24827 41309
rect 24894 41306 24900 41308
rect 24761 41304 24900 41306
rect 24761 41248 24766 41304
rect 24822 41248 24900 41304
rect 24761 41246 24900 41248
rect 24761 41243 24827 41246
rect 24894 41244 24900 41246
rect 24964 41244 24970 41308
rect 26509 41306 26575 41309
rect 27294 41306 27354 41654
rect 27521 41651 27587 41654
rect 27662 41578 27722 41790
rect 28165 41716 28231 41717
rect 30741 41716 30807 41717
rect 28165 41712 28212 41716
rect 28276 41714 28282 41716
rect 30046 41714 30052 41716
rect 28165 41656 28170 41712
rect 28165 41652 28212 41656
rect 28276 41654 28322 41714
rect 29870 41654 30052 41714
rect 28276 41652 28282 41654
rect 28165 41651 28231 41652
rect 26509 41304 27354 41306
rect 26509 41248 26514 41304
rect 26570 41248 27354 41304
rect 26509 41246 27354 41248
rect 27478 41518 27722 41578
rect 26509 41243 26575 41246
rect 24209 41170 24275 41173
rect 25405 41172 25471 41173
rect 26969 41172 27035 41173
rect 24342 41170 24348 41172
rect 24209 41168 24348 41170
rect 24209 41112 24214 41168
rect 24270 41112 24348 41168
rect 24209 41110 24348 41112
rect 24209 41107 24275 41110
rect 24342 41108 24348 41110
rect 24412 41108 24418 41172
rect 25405 41168 25452 41172
rect 25516 41170 25522 41172
rect 25405 41112 25410 41168
rect 25405 41108 25452 41112
rect 25516 41110 25562 41170
rect 25516 41108 25522 41110
rect 26918 41108 26924 41172
rect 26988 41170 27035 41172
rect 26988 41168 27080 41170
rect 27030 41112 27080 41168
rect 26988 41110 27080 41112
rect 26988 41108 27035 41110
rect 25405 41107 25471 41108
rect 26969 41107 27035 41108
rect 27478 41037 27538 41518
rect 28073 41440 28139 41445
rect 28073 41384 28078 41440
rect 28134 41384 28139 41440
rect 28073 41379 28139 41384
rect 28257 41442 28323 41445
rect 28533 41442 28599 41445
rect 28257 41440 28599 41442
rect 28257 41384 28262 41440
rect 28318 41384 28538 41440
rect 28594 41384 28599 41440
rect 28257 41382 28599 41384
rect 28257 41379 28323 41382
rect 28533 41379 28599 41382
rect 28717 41442 28783 41445
rect 29729 41442 29795 41445
rect 28717 41440 29795 41442
rect 28717 41384 28722 41440
rect 28778 41384 29734 41440
rect 29790 41384 29795 41440
rect 28717 41382 29795 41384
rect 29870 41442 29930 41654
rect 30046 41652 30052 41654
rect 30116 41652 30122 41716
rect 30741 41714 30788 41716
rect 30696 41712 30788 41714
rect 30696 41656 30746 41712
rect 30696 41654 30788 41656
rect 30741 41652 30788 41654
rect 30852 41652 30858 41716
rect 30974 41714 31034 41790
rect 30974 41654 31218 41714
rect 30741 41651 30807 41652
rect 31158 41608 31218 41654
rect 30281 41576 30347 41581
rect 30833 41580 30899 41581
rect 30281 41520 30286 41576
rect 30342 41520 30347 41576
rect 30281 41515 30347 41520
rect 30782 41516 30788 41580
rect 30852 41578 30899 41580
rect 30852 41576 30944 41578
rect 30894 41520 30944 41576
rect 30852 41518 30944 41520
rect 31158 41518 32000 41608
rect 30852 41516 30899 41518
rect 30833 41515 30899 41516
rect 30005 41442 30071 41445
rect 29870 41440 30071 41442
rect 29870 41384 30010 41440
rect 30066 41384 30071 41440
rect 29870 41382 30071 41384
rect 28717 41379 28783 41382
rect 29729 41379 29795 41382
rect 30005 41379 30071 41382
rect 28076 41308 28136 41379
rect 28022 41244 28028 41308
rect 28092 41246 28136 41308
rect 30284 41306 30344 41515
rect 31200 41488 32000 41518
rect 28260 41246 30344 41306
rect 28092 41244 28098 41246
rect 27705 41170 27771 41173
rect 28260 41170 28320 41246
rect 27705 41168 28320 41170
rect 27705 41112 27710 41168
rect 27766 41112 28320 41168
rect 27705 41110 28320 41112
rect 28533 41170 28599 41173
rect 28901 41170 28967 41173
rect 29545 41170 29611 41173
rect 30598 41170 30604 41172
rect 28533 41168 29010 41170
rect 28533 41112 28538 41168
rect 28594 41112 28906 41168
rect 28962 41112 29010 41168
rect 28533 41110 29010 41112
rect 27705 41107 27771 41110
rect 28533 41107 28599 41110
rect 28901 41107 29010 41110
rect 29545 41168 30604 41170
rect 29545 41112 29550 41168
rect 29606 41112 30604 41168
rect 29545 41110 30604 41112
rect 29545 41107 29611 41110
rect 30598 41108 30604 41110
rect 30668 41108 30674 41172
rect 25957 41034 26023 41037
rect 25592 41032 26023 41034
rect 25592 40976 25962 41032
rect 26018 40976 26023 41032
rect 25592 40974 26023 40976
rect 27478 41032 27587 41037
rect 27705 41036 27771 41037
rect 27478 40976 27526 41032
rect 27582 40976 27587 41032
rect 27478 40974 27587 40976
rect 21265 40898 21331 40901
rect 23289 40898 23355 40901
rect 21265 40896 23355 40898
rect 21265 40840 21270 40896
rect 21326 40840 23294 40896
rect 23350 40840 23355 40896
rect 21265 40838 23355 40840
rect 21265 40835 21331 40838
rect 23289 40835 23355 40838
rect 25221 40898 25287 40901
rect 25446 40898 25452 40900
rect 25221 40896 25452 40898
rect 25221 40840 25226 40896
rect 25282 40840 25452 40896
rect 25221 40838 25452 40840
rect 25221 40835 25287 40838
rect 25446 40836 25452 40838
rect 25516 40836 25522 40900
rect 5909 40832 6229 40833
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6229 40832
rect 5909 40767 6229 40768
rect 15840 40832 16160 40833
rect 15840 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15840 40767 16160 40768
rect 24025 40762 24091 40765
rect 25221 40762 25287 40765
rect 25592 40762 25652 40974
rect 25957 40971 26023 40974
rect 27521 40971 27587 40974
rect 27654 40972 27660 41036
rect 27724 41034 27771 41036
rect 27724 41032 27816 41034
rect 27766 40976 27816 41032
rect 27724 40974 27816 40976
rect 27981 41032 28047 41037
rect 27981 40976 27986 41032
rect 28042 40976 28047 41032
rect 27724 40972 27771 40974
rect 27705 40971 27771 40972
rect 27981 40971 28047 40976
rect 28809 41032 28875 41037
rect 28809 40976 28814 41032
rect 28870 40976 28875 41032
rect 28809 40971 28875 40976
rect 27984 40901 28044 40971
rect 27286 40836 27292 40900
rect 27356 40898 27362 40900
rect 27654 40898 27660 40900
rect 27356 40838 27660 40898
rect 27356 40836 27362 40838
rect 27654 40836 27660 40838
rect 27724 40836 27730 40900
rect 27981 40896 28047 40901
rect 27981 40840 27986 40896
rect 28042 40840 28047 40896
rect 27981 40835 28047 40840
rect 28625 40898 28691 40901
rect 28812 40898 28872 40971
rect 28625 40896 28872 40898
rect 28625 40840 28630 40896
rect 28686 40840 28872 40896
rect 28625 40838 28872 40840
rect 28950 40901 29010 41107
rect 29126 40972 29132 41036
rect 29196 41034 29202 41036
rect 29545 41034 29611 41037
rect 29196 41032 29611 41034
rect 29196 40976 29550 41032
rect 29606 40976 29611 41032
rect 29196 40974 29611 40976
rect 29196 40972 29202 40974
rect 28950 40896 29059 40901
rect 28950 40840 28998 40896
rect 29054 40840 29059 40896
rect 28950 40838 29059 40840
rect 28625 40835 28691 40838
rect 28993 40835 29059 40838
rect 25770 40832 26090 40833
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26090 40832
rect 25770 40767 26090 40768
rect 29134 40762 29194 40972
rect 29545 40971 29611 40974
rect 29913 41034 29979 41037
rect 31200 41034 32000 41064
rect 29913 41032 32000 41034
rect 29913 40976 29918 41032
rect 29974 40976 32000 41032
rect 29913 40974 32000 40976
rect 29913 40971 29979 40974
rect 31200 40944 32000 40974
rect 24025 40760 25652 40762
rect 24025 40704 24030 40760
rect 24086 40704 25226 40760
rect 25282 40704 25652 40760
rect 24025 40702 25652 40704
rect 26374 40702 29194 40762
rect 30649 40762 30715 40765
rect 30782 40762 30788 40764
rect 30649 40760 30788 40762
rect 30649 40704 30654 40760
rect 30710 40704 30788 40760
rect 30649 40702 30788 40704
rect 24025 40699 24091 40702
rect 25221 40699 25287 40702
rect 0 40626 800 40656
rect 1577 40626 1643 40629
rect 0 40624 1643 40626
rect 0 40568 1582 40624
rect 1638 40568 1643 40624
rect 0 40566 1643 40568
rect 0 40536 800 40566
rect 1577 40563 1643 40566
rect 19885 40626 19951 40629
rect 26374 40626 26434 40702
rect 30649 40699 30715 40702
rect 30782 40700 30788 40702
rect 30852 40700 30858 40764
rect 31200 40626 32000 40656
rect 19885 40624 26434 40626
rect 19885 40568 19890 40624
rect 19946 40568 26434 40624
rect 19885 40566 26434 40568
rect 26512 40566 32000 40626
rect 19885 40563 19951 40566
rect 25129 40490 25195 40493
rect 25865 40490 25931 40493
rect 25129 40488 25931 40490
rect 25129 40432 25134 40488
rect 25190 40432 25870 40488
rect 25926 40432 25931 40488
rect 25129 40430 25931 40432
rect 25129 40427 25195 40430
rect 25865 40427 25931 40430
rect 26049 40490 26115 40493
rect 26325 40490 26391 40493
rect 26049 40488 26391 40490
rect 26049 40432 26054 40488
rect 26110 40432 26330 40488
rect 26386 40432 26391 40488
rect 26049 40430 26391 40432
rect 26049 40427 26115 40430
rect 26325 40427 26391 40430
rect 25630 40292 25636 40356
rect 25700 40354 25706 40356
rect 25773 40354 25839 40357
rect 25700 40352 25839 40354
rect 25700 40296 25778 40352
rect 25834 40296 25839 40352
rect 25700 40294 25839 40296
rect 25700 40292 25706 40294
rect 25773 40291 25839 40294
rect 10874 40288 11194 40289
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 40223 11194 40224
rect 20805 40288 21125 40289
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 40223 21125 40224
rect 22093 40218 22159 40221
rect 26512 40218 26572 40566
rect 31200 40536 32000 40566
rect 29637 40490 29703 40493
rect 30046 40490 30052 40492
rect 29637 40488 30052 40490
rect 29637 40432 29642 40488
rect 29698 40432 30052 40488
rect 29637 40430 30052 40432
rect 29637 40427 29703 40430
rect 30046 40428 30052 40430
rect 30116 40428 30122 40492
rect 22093 40216 26572 40218
rect 22093 40160 22098 40216
rect 22154 40160 26572 40216
rect 22093 40158 26572 40160
rect 27797 40218 27863 40221
rect 31200 40218 32000 40248
rect 27797 40216 32000 40218
rect 27797 40160 27802 40216
rect 27858 40160 32000 40216
rect 27797 40158 32000 40160
rect 22093 40155 22159 40158
rect 27797 40155 27863 40158
rect 31200 40128 32000 40158
rect 27470 40020 27476 40084
rect 27540 40082 27546 40084
rect 27797 40082 27863 40085
rect 27540 40080 27863 40082
rect 27540 40024 27802 40080
rect 27858 40024 27863 40080
rect 27540 40022 27863 40024
rect 27540 40020 27546 40022
rect 27797 40019 27863 40022
rect 0 39946 800 39976
rect 1577 39946 1643 39949
rect 0 39944 1643 39946
rect 0 39888 1582 39944
rect 1638 39888 1643 39944
rect 0 39886 1643 39888
rect 0 39856 800 39886
rect 1577 39883 1643 39886
rect 24158 39884 24164 39948
rect 24228 39946 24234 39948
rect 28165 39946 28231 39949
rect 24228 39944 28231 39946
rect 24228 39888 28170 39944
rect 28226 39888 28231 39944
rect 24228 39886 28231 39888
rect 24228 39884 24234 39886
rect 28165 39883 28231 39886
rect 30782 39884 30788 39948
rect 30852 39946 30858 39948
rect 31886 39946 31892 39948
rect 30852 39886 31892 39946
rect 30852 39884 30858 39886
rect 31886 39884 31892 39886
rect 31956 39884 31962 39948
rect 27102 39748 27108 39812
rect 27172 39810 27178 39812
rect 28533 39810 28599 39813
rect 27172 39808 28599 39810
rect 27172 39752 28538 39808
rect 28594 39752 28599 39808
rect 27172 39750 28599 39752
rect 27172 39748 27178 39750
rect 28533 39747 28599 39750
rect 5909 39744 6229 39745
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6229 39744
rect 5909 39679 6229 39680
rect 15840 39744 16160 39745
rect 15840 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15840 39679 16160 39680
rect 25770 39744 26090 39745
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26090 39744
rect 25770 39679 26090 39680
rect 27613 39674 27679 39677
rect 31200 39674 32000 39704
rect 27613 39672 32000 39674
rect 27613 39616 27618 39672
rect 27674 39616 32000 39672
rect 27613 39614 32000 39616
rect 27613 39611 27679 39614
rect 31200 39584 32000 39614
rect 26141 39540 26207 39541
rect 26141 39536 26188 39540
rect 26252 39538 26258 39540
rect 26141 39480 26146 39536
rect 26141 39476 26188 39480
rect 26252 39478 26298 39538
rect 26252 39476 26258 39478
rect 26141 39475 26207 39476
rect 25957 39402 26023 39405
rect 26366 39402 26372 39404
rect 25957 39400 26372 39402
rect 25957 39344 25962 39400
rect 26018 39344 26372 39400
rect 25957 39342 26372 39344
rect 25957 39339 26023 39342
rect 26366 39340 26372 39342
rect 26436 39340 26442 39404
rect 29126 39340 29132 39404
rect 29196 39402 29202 39404
rect 30414 39402 30420 39404
rect 29196 39342 30420 39402
rect 29196 39340 29202 39342
rect 30414 39340 30420 39342
rect 30484 39340 30490 39404
rect 0 39266 800 39296
rect 1577 39266 1643 39269
rect 26417 39268 26483 39269
rect 0 39264 1643 39266
rect 0 39208 1582 39264
rect 1638 39208 1643 39264
rect 0 39206 1643 39208
rect 0 39176 800 39206
rect 1577 39203 1643 39206
rect 26366 39204 26372 39268
rect 26436 39266 26483 39268
rect 28165 39266 28231 39269
rect 31200 39266 32000 39296
rect 26436 39264 26528 39266
rect 26478 39208 26528 39264
rect 26436 39206 26528 39208
rect 28165 39264 32000 39266
rect 28165 39208 28170 39264
rect 28226 39208 32000 39264
rect 28165 39206 32000 39208
rect 26436 39204 26483 39206
rect 26417 39203 26483 39204
rect 28165 39203 28231 39206
rect 10874 39200 11194 39201
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 39135 11194 39136
rect 20805 39200 21125 39201
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 31200 39176 32000 39206
rect 20805 39135 21125 39136
rect 26325 39128 26391 39133
rect 26325 39072 26330 39128
rect 26386 39072 26391 39128
rect 26325 39067 26391 39072
rect 23606 38932 23612 38996
rect 23676 38994 23682 38996
rect 23841 38994 23907 38997
rect 23676 38992 23907 38994
rect 23676 38936 23846 38992
rect 23902 38936 23907 38992
rect 23676 38934 23907 38936
rect 23676 38932 23682 38934
rect 23841 38931 23907 38934
rect 25865 38994 25931 38997
rect 26182 38994 26188 38996
rect 25865 38992 26188 38994
rect 25865 38936 25870 38992
rect 25926 38936 26188 38992
rect 25865 38934 26188 38936
rect 25865 38931 25931 38934
rect 26182 38932 26188 38934
rect 26252 38932 26258 38996
rect 24577 38858 24643 38861
rect 24534 38856 24643 38858
rect 24534 38800 24582 38856
rect 24638 38800 24643 38856
rect 24534 38795 24643 38800
rect 25630 38796 25636 38860
rect 25700 38858 25706 38860
rect 25865 38858 25931 38861
rect 25700 38856 25931 38858
rect 25700 38800 25870 38856
rect 25926 38800 25931 38856
rect 25700 38798 25931 38800
rect 25700 38796 25706 38798
rect 25865 38795 25931 38798
rect 12065 38722 12131 38725
rect 14089 38722 14155 38725
rect 12065 38720 14155 38722
rect 12065 38664 12070 38720
rect 12126 38664 14094 38720
rect 14150 38664 14155 38720
rect 12065 38662 14155 38664
rect 12065 38659 12131 38662
rect 14089 38659 14155 38662
rect 5909 38656 6229 38657
rect 0 38586 800 38616
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6229 38656
rect 5909 38591 6229 38592
rect 15840 38656 16160 38657
rect 15840 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15840 38591 16160 38592
rect 1577 38586 1643 38589
rect 0 38584 1643 38586
rect 0 38528 1582 38584
rect 1638 38528 1643 38584
rect 0 38526 1643 38528
rect 0 38496 800 38526
rect 1577 38523 1643 38526
rect 24534 38453 24594 38795
rect 26328 38725 26388 39067
rect 26509 38992 26575 38997
rect 26509 38936 26514 38992
rect 26570 38936 26575 38992
rect 26509 38931 26575 38936
rect 30414 38932 30420 38996
rect 30484 38994 30490 38996
rect 31702 38994 31708 38996
rect 30484 38934 31708 38994
rect 30484 38932 30490 38934
rect 31702 38932 31708 38934
rect 31772 38932 31778 38996
rect 26512 38861 26572 38931
rect 26509 38856 26575 38861
rect 26509 38800 26514 38856
rect 26570 38800 26575 38856
rect 26509 38795 26575 38800
rect 26325 38720 26391 38725
rect 24669 38670 24735 38673
rect 24669 38668 24778 38670
rect 24669 38612 24674 38668
rect 24730 38612 24778 38668
rect 24669 38607 24778 38612
rect 24853 38668 24919 38673
rect 24853 38612 24858 38668
rect 24914 38612 24919 38668
rect 26325 38664 26330 38720
rect 26386 38664 26391 38720
rect 26325 38659 26391 38664
rect 28901 38722 28967 38725
rect 31200 38722 32000 38752
rect 28901 38720 32000 38722
rect 28901 38664 28906 38720
rect 28962 38664 32000 38720
rect 28901 38662 32000 38664
rect 28901 38659 28967 38662
rect 24853 38607 24919 38612
rect 25770 38656 26090 38657
rect 23381 38450 23447 38453
rect 24534 38450 24643 38453
rect 23381 38448 24643 38450
rect 23381 38392 23386 38448
rect 23442 38392 24582 38448
rect 24638 38392 24643 38448
rect 23381 38390 24643 38392
rect 23381 38387 23447 38390
rect 24577 38387 24643 38390
rect 24718 38317 24778 38607
rect 24856 38452 24916 38607
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26090 38656
rect 31200 38632 32000 38662
rect 25770 38591 26090 38592
rect 25262 38524 25268 38588
rect 25332 38586 25338 38588
rect 25589 38586 25655 38589
rect 26417 38588 26483 38589
rect 26366 38586 26372 38588
rect 25332 38584 25655 38586
rect 25332 38528 25594 38584
rect 25650 38528 25655 38584
rect 25332 38526 25655 38528
rect 26326 38526 26372 38586
rect 26436 38584 26483 38588
rect 26478 38528 26483 38584
rect 25332 38524 25338 38526
rect 25589 38523 25655 38526
rect 26366 38524 26372 38526
rect 26436 38524 26483 38528
rect 26417 38523 26483 38524
rect 24856 38390 24900 38452
rect 24894 38388 24900 38390
rect 24964 38388 24970 38452
rect 25773 38450 25839 38453
rect 26049 38450 26115 38453
rect 27981 38452 28047 38453
rect 27981 38450 28028 38452
rect 25773 38448 26115 38450
rect 25773 38392 25778 38448
rect 25834 38392 26054 38448
rect 26110 38392 26115 38448
rect 25773 38390 26115 38392
rect 27936 38448 28028 38450
rect 27936 38392 27986 38448
rect 27936 38390 28028 38392
rect 25773 38387 25839 38390
rect 26049 38387 26115 38390
rect 27981 38388 28028 38390
rect 28092 38388 28098 38452
rect 27981 38387 28047 38388
rect 21725 38314 21791 38317
rect 24526 38314 24532 38316
rect 21725 38312 24532 38314
rect 21725 38256 21730 38312
rect 21786 38256 24532 38312
rect 21725 38254 24532 38256
rect 21725 38251 21791 38254
rect 24526 38252 24532 38254
rect 24596 38252 24602 38316
rect 24669 38312 24778 38317
rect 28165 38314 28231 38317
rect 24669 38256 24674 38312
rect 24730 38256 24778 38312
rect 24669 38254 24778 38256
rect 25776 38312 28231 38314
rect 25776 38256 28170 38312
rect 28226 38256 28231 38312
rect 25776 38254 28231 38256
rect 24669 38251 24735 38254
rect 22185 38178 22251 38181
rect 24853 38178 24919 38181
rect 25078 38178 25084 38180
rect 22185 38176 24778 38178
rect 22185 38120 22190 38176
rect 22246 38120 24778 38176
rect 22185 38118 24778 38120
rect 22185 38115 22251 38118
rect 10874 38112 11194 38113
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 38047 11194 38048
rect 20805 38112 21125 38113
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 38047 21125 38048
rect 23565 38044 23631 38045
rect 23565 38042 23612 38044
rect 23520 38040 23612 38042
rect 23520 37984 23570 38040
rect 23520 37982 23612 37984
rect 23565 37980 23612 37982
rect 23676 37980 23682 38044
rect 24718 38042 24778 38118
rect 24853 38176 25084 38178
rect 24853 38120 24858 38176
rect 24914 38120 25084 38176
rect 24853 38118 25084 38120
rect 24853 38115 24919 38118
rect 25078 38116 25084 38118
rect 25148 38116 25154 38180
rect 25446 38116 25452 38180
rect 25516 38178 25522 38180
rect 25589 38178 25655 38181
rect 25516 38176 25655 38178
rect 25516 38120 25594 38176
rect 25650 38120 25655 38176
rect 25516 38118 25655 38120
rect 25516 38116 25522 38118
rect 25589 38115 25655 38118
rect 25776 38042 25836 38254
rect 28165 38251 28231 38254
rect 28625 38314 28691 38317
rect 31200 38314 32000 38344
rect 28625 38312 32000 38314
rect 28625 38256 28630 38312
rect 28686 38256 32000 38312
rect 28625 38254 32000 38256
rect 28625 38251 28691 38254
rect 31200 38224 32000 38254
rect 26601 38178 26667 38181
rect 26918 38178 26924 38180
rect 26601 38176 26924 38178
rect 26601 38120 26606 38176
rect 26662 38120 26924 38176
rect 26601 38118 26924 38120
rect 26601 38115 26667 38118
rect 26918 38116 26924 38118
rect 26988 38116 26994 38180
rect 28022 38116 28028 38180
rect 28092 38178 28098 38180
rect 29453 38178 29519 38181
rect 28092 38176 29519 38178
rect 28092 38120 29458 38176
rect 29514 38120 29519 38176
rect 28092 38118 29519 38120
rect 28092 38116 28098 38118
rect 29453 38115 29519 38118
rect 24718 37982 25836 38042
rect 28625 38042 28691 38045
rect 31150 38042 31156 38044
rect 28625 38040 31156 38042
rect 28625 37984 28630 38040
rect 28686 37984 31156 38040
rect 28625 37982 31156 37984
rect 23565 37979 23631 37980
rect 28625 37979 28691 37982
rect 31150 37980 31156 37982
rect 31220 37980 31226 38044
rect 31334 37980 31340 38044
rect 31404 38042 31410 38044
rect 31845 38042 31911 38045
rect 31404 38040 31911 38042
rect 31404 37984 31850 38040
rect 31906 37984 31911 38040
rect 31404 37982 31911 37984
rect 31404 37980 31410 37982
rect 31845 37979 31911 37982
rect 0 37906 800 37936
rect 1577 37906 1643 37909
rect 0 37904 1643 37906
rect 0 37848 1582 37904
rect 1638 37848 1643 37904
rect 0 37846 1643 37848
rect 0 37816 800 37846
rect 1577 37843 1643 37846
rect 22921 37906 22987 37909
rect 24853 37906 24919 37909
rect 22921 37904 24919 37906
rect 22921 37848 22926 37904
rect 22982 37848 24858 37904
rect 24914 37848 24919 37904
rect 22921 37846 24919 37848
rect 22921 37843 22987 37846
rect 24853 37843 24919 37846
rect 25446 37844 25452 37908
rect 25516 37906 25522 37908
rect 26182 37906 26188 37908
rect 25516 37846 26188 37906
rect 25516 37844 25522 37846
rect 26182 37844 26188 37846
rect 26252 37844 26258 37908
rect 24025 37772 24091 37773
rect 23974 37708 23980 37772
rect 24044 37770 24091 37772
rect 24044 37768 24136 37770
rect 24086 37712 24136 37768
rect 24044 37710 24136 37712
rect 24044 37708 24091 37710
rect 27470 37708 27476 37772
rect 27540 37770 27546 37772
rect 28717 37770 28783 37773
rect 27540 37768 28783 37770
rect 27540 37712 28722 37768
rect 28778 37712 28783 37768
rect 27540 37710 28783 37712
rect 27540 37708 27546 37710
rect 24025 37707 24091 37708
rect 28717 37707 28783 37710
rect 30005 37770 30071 37773
rect 31200 37770 32000 37800
rect 30005 37768 32000 37770
rect 30005 37712 30010 37768
rect 30066 37712 32000 37768
rect 30005 37710 32000 37712
rect 30005 37707 30071 37710
rect 31200 37680 32000 37710
rect 24853 37636 24919 37637
rect 24853 37632 24900 37636
rect 24964 37634 24970 37636
rect 24853 37576 24858 37632
rect 24853 37572 24900 37576
rect 24964 37574 25010 37634
rect 24964 37572 24970 37574
rect 24853 37571 24919 37572
rect 5909 37568 6229 37569
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6229 37568
rect 5909 37503 6229 37504
rect 15840 37568 16160 37569
rect 15840 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15840 37503 16160 37504
rect 25770 37568 26090 37569
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26090 37568
rect 25770 37503 26090 37504
rect 18689 37498 18755 37501
rect 24710 37498 24716 37500
rect 18689 37496 24716 37498
rect 18689 37440 18694 37496
rect 18750 37440 24716 37496
rect 18689 37438 24716 37440
rect 18689 37435 18755 37438
rect 24710 37436 24716 37438
rect 24780 37498 24786 37500
rect 25221 37498 25287 37501
rect 26918 37498 26924 37500
rect 24780 37496 25287 37498
rect 24780 37440 25226 37496
rect 25282 37440 25287 37496
rect 24780 37438 25287 37440
rect 24780 37436 24786 37438
rect 25221 37435 25287 37438
rect 26190 37438 26924 37498
rect 0 37362 800 37392
rect 1393 37362 1459 37365
rect 0 37360 1459 37362
rect 0 37304 1398 37360
rect 1454 37304 1459 37360
rect 0 37302 1459 37304
rect 0 37272 800 37302
rect 1393 37299 1459 37302
rect 18229 37362 18295 37365
rect 18965 37362 19031 37365
rect 18229 37360 19031 37362
rect 18229 37304 18234 37360
rect 18290 37304 18970 37360
rect 19026 37304 19031 37360
rect 18229 37302 19031 37304
rect 18229 37299 18295 37302
rect 18965 37299 19031 37302
rect 19885 37362 19951 37365
rect 26190 37362 26250 37438
rect 26918 37436 26924 37438
rect 26988 37436 26994 37500
rect 19885 37360 26250 37362
rect 19885 37304 19890 37360
rect 19946 37304 26250 37360
rect 19885 37302 26250 37304
rect 19885 37299 19951 37302
rect 26366 37300 26372 37364
rect 26436 37362 26442 37364
rect 27981 37362 28047 37365
rect 26436 37360 28047 37362
rect 26436 37304 27986 37360
rect 28042 37304 28047 37360
rect 26436 37302 28047 37304
rect 26436 37300 26442 37302
rect 27981 37299 28047 37302
rect 29361 37362 29427 37365
rect 31200 37362 32000 37392
rect 29361 37360 32000 37362
rect 29361 37304 29366 37360
rect 29422 37304 32000 37360
rect 29361 37302 32000 37304
rect 29361 37299 29427 37302
rect 31200 37272 32000 37302
rect 25262 37164 25268 37228
rect 25332 37226 25338 37228
rect 25497 37226 25563 37229
rect 25332 37224 25563 37226
rect 25332 37168 25502 37224
rect 25558 37168 25563 37224
rect 25332 37166 25563 37168
rect 25332 37164 25338 37166
rect 25497 37163 25563 37166
rect 28257 37226 28323 37229
rect 30414 37226 30420 37228
rect 28257 37224 30420 37226
rect 28257 37168 28262 37224
rect 28318 37168 30420 37224
rect 28257 37166 30420 37168
rect 28257 37163 28323 37166
rect 30414 37164 30420 37166
rect 30484 37164 30490 37228
rect 26049 37090 26115 37093
rect 26734 37090 26740 37092
rect 26049 37088 26740 37090
rect 26049 37032 26054 37088
rect 26110 37032 26740 37088
rect 26049 37030 26740 37032
rect 26049 37027 26115 37030
rect 26734 37028 26740 37030
rect 26804 37028 26810 37092
rect 31150 37028 31156 37092
rect 31220 37090 31226 37092
rect 31385 37090 31451 37093
rect 31220 37088 31451 37090
rect 31220 37032 31390 37088
rect 31446 37032 31451 37088
rect 31220 37030 31451 37032
rect 31220 37028 31226 37030
rect 31385 37027 31451 37030
rect 10874 37024 11194 37025
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 36959 11194 36960
rect 20805 37024 21125 37025
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 20805 36959 21125 36960
rect 15377 36954 15443 36957
rect 15929 36954 15995 36957
rect 15377 36952 15995 36954
rect 15377 36896 15382 36952
rect 15438 36896 15934 36952
rect 15990 36896 15995 36952
rect 15377 36894 15995 36896
rect 15377 36891 15443 36894
rect 15929 36891 15995 36894
rect 22921 36954 22987 36957
rect 28257 36954 28323 36957
rect 22921 36952 28323 36954
rect 22921 36896 22926 36952
rect 22982 36896 28262 36952
rect 28318 36896 28323 36952
rect 22921 36894 28323 36896
rect 22921 36891 22987 36894
rect 28257 36891 28323 36894
rect 9489 36818 9555 36821
rect 29821 36818 29887 36821
rect 9489 36816 29887 36818
rect 9489 36760 9494 36816
rect 9550 36760 29826 36816
rect 29882 36760 29887 36816
rect 9489 36758 29887 36760
rect 9489 36755 9555 36758
rect 29821 36755 29887 36758
rect 30005 36818 30071 36821
rect 31200 36818 32000 36848
rect 30005 36816 32000 36818
rect 30005 36760 30010 36816
rect 30066 36760 32000 36816
rect 30005 36758 32000 36760
rect 30005 36755 30071 36758
rect 31200 36728 32000 36758
rect 0 36682 800 36712
rect 1577 36682 1643 36685
rect 0 36680 1643 36682
rect 0 36624 1582 36680
rect 1638 36624 1643 36680
rect 0 36622 1643 36624
rect 0 36592 800 36622
rect 1577 36619 1643 36622
rect 10409 36682 10475 36685
rect 15837 36682 15903 36685
rect 10409 36680 15903 36682
rect 10409 36624 10414 36680
rect 10470 36624 15842 36680
rect 15898 36624 15903 36680
rect 10409 36622 15903 36624
rect 10409 36619 10475 36622
rect 15837 36619 15903 36622
rect 24894 36620 24900 36684
rect 24964 36682 24970 36684
rect 25681 36682 25747 36685
rect 24964 36680 25747 36682
rect 24964 36624 25686 36680
rect 25742 36624 25747 36680
rect 24964 36622 25747 36624
rect 24964 36620 24970 36622
rect 25681 36619 25747 36622
rect 26417 36682 26483 36685
rect 26550 36682 26556 36684
rect 26417 36680 26556 36682
rect 26417 36624 26422 36680
rect 26478 36624 26556 36680
rect 26417 36622 26556 36624
rect 26417 36619 26483 36622
rect 26550 36620 26556 36622
rect 26620 36620 26626 36684
rect 26693 36682 26759 36685
rect 30005 36684 30071 36685
rect 26693 36680 26802 36682
rect 26693 36624 26698 36680
rect 26754 36624 26802 36680
rect 26693 36619 26802 36624
rect 30005 36680 30052 36684
rect 30116 36682 30122 36684
rect 30005 36624 30010 36680
rect 30005 36620 30052 36624
rect 30116 36622 30162 36682
rect 30116 36620 30122 36622
rect 30005 36619 30071 36620
rect 5909 36480 6229 36481
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6229 36480
rect 5909 36415 6229 36416
rect 15840 36480 16160 36481
rect 15840 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15840 36415 16160 36416
rect 25770 36480 26090 36481
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26090 36480
rect 25770 36415 26090 36416
rect 26601 36410 26667 36413
rect 26742 36410 26802 36619
rect 29913 36546 29979 36549
rect 29913 36544 30114 36546
rect 29913 36488 29918 36544
rect 29974 36488 30114 36544
rect 29913 36486 30114 36488
rect 29913 36483 29979 36486
rect 26601 36408 26802 36410
rect 26601 36352 26606 36408
rect 26662 36352 26802 36408
rect 26601 36350 26802 36352
rect 30054 36410 30114 36486
rect 31200 36410 32000 36440
rect 30054 36350 32000 36410
rect 26601 36347 26667 36350
rect 31200 36320 32000 36350
rect 26509 36274 26575 36277
rect 24902 36272 26575 36274
rect 24902 36216 26514 36272
rect 26570 36216 26575 36272
rect 24902 36214 26575 36216
rect 24761 36138 24827 36141
rect 24902 36138 24962 36214
rect 26509 36211 26575 36214
rect 29913 36274 29979 36277
rect 30966 36274 30972 36276
rect 29913 36272 30972 36274
rect 29913 36216 29918 36272
rect 29974 36216 30972 36272
rect 29913 36214 30972 36216
rect 29913 36211 29979 36214
rect 30966 36212 30972 36214
rect 31036 36212 31042 36276
rect 24761 36136 24962 36138
rect 24761 36080 24766 36136
rect 24822 36080 24962 36136
rect 24761 36078 24962 36080
rect 24761 36075 24827 36078
rect 25446 36076 25452 36140
rect 25516 36138 25522 36140
rect 25589 36138 25655 36141
rect 25516 36136 25655 36138
rect 25516 36080 25594 36136
rect 25650 36080 25655 36136
rect 25516 36078 25655 36080
rect 25516 36076 25522 36078
rect 25589 36075 25655 36078
rect 31293 36138 31359 36141
rect 31518 36138 31524 36140
rect 31293 36136 31524 36138
rect 31293 36080 31298 36136
rect 31354 36080 31524 36136
rect 31293 36078 31524 36080
rect 31293 36075 31359 36078
rect 31518 36076 31524 36078
rect 31588 36076 31594 36140
rect 0 36002 800 36032
rect 1577 36002 1643 36005
rect 0 36000 1643 36002
rect 0 35944 1582 36000
rect 1638 35944 1643 36000
rect 0 35942 1643 35944
rect 0 35912 800 35942
rect 1577 35939 1643 35942
rect 25446 35940 25452 36004
rect 25516 36002 25522 36004
rect 26049 36002 26115 36005
rect 25516 36000 26115 36002
rect 25516 35944 26054 36000
rect 26110 35944 26115 36000
rect 25516 35942 26115 35944
rect 25516 35940 25522 35942
rect 26049 35939 26115 35942
rect 10874 35936 11194 35937
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 35871 11194 35872
rect 20805 35936 21125 35937
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 20805 35871 21125 35872
rect 25078 35804 25084 35868
rect 25148 35866 25154 35868
rect 25865 35866 25931 35869
rect 25148 35864 25931 35866
rect 25148 35808 25870 35864
rect 25926 35808 25931 35864
rect 25148 35806 25931 35808
rect 25148 35804 25154 35806
rect 25865 35803 25931 35806
rect 30189 35866 30255 35869
rect 31200 35866 32000 35896
rect 30189 35864 32000 35866
rect 30189 35808 30194 35864
rect 30250 35808 32000 35864
rect 30189 35806 32000 35808
rect 30189 35803 30255 35806
rect 31200 35776 32000 35806
rect 25262 35668 25268 35732
rect 25332 35730 25338 35732
rect 25773 35730 25839 35733
rect 25332 35728 25839 35730
rect 25332 35672 25778 35728
rect 25834 35672 25839 35728
rect 25332 35670 25839 35672
rect 25332 35668 25338 35670
rect 25773 35667 25839 35670
rect 27521 35730 27587 35733
rect 28257 35730 28323 35733
rect 27521 35728 28323 35730
rect 27521 35672 27526 35728
rect 27582 35672 28262 35728
rect 28318 35672 28323 35728
rect 27521 35670 28323 35672
rect 27521 35667 27587 35670
rect 28257 35667 28323 35670
rect 27613 35458 27679 35461
rect 31200 35458 32000 35488
rect 27613 35456 32000 35458
rect 27613 35400 27618 35456
rect 27674 35400 32000 35456
rect 27613 35398 32000 35400
rect 27613 35395 27679 35398
rect 5909 35392 6229 35393
rect 0 35322 800 35352
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6229 35392
rect 5909 35327 6229 35328
rect 15840 35392 16160 35393
rect 15840 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15840 35327 16160 35328
rect 25770 35392 26090 35393
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26090 35392
rect 31200 35368 32000 35398
rect 25770 35327 26090 35328
rect 1577 35322 1643 35325
rect 24117 35324 24183 35325
rect 24117 35322 24164 35324
rect 0 35320 1643 35322
rect 0 35264 1582 35320
rect 1638 35264 1643 35320
rect 0 35262 1643 35264
rect 24072 35320 24164 35322
rect 24072 35264 24122 35320
rect 24072 35262 24164 35264
rect 0 35232 800 35262
rect 1577 35259 1643 35262
rect 24117 35260 24164 35262
rect 24228 35260 24234 35324
rect 24117 35259 24183 35260
rect 19701 35050 19767 35053
rect 19701 35048 19810 35050
rect 19701 34992 19706 35048
rect 19762 34992 19810 35048
rect 19701 34987 19810 34992
rect 10874 34848 11194 34849
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 34783 11194 34784
rect 0 34642 800 34672
rect 19750 34645 19810 34987
rect 28165 34914 28231 34917
rect 31200 34914 32000 34944
rect 28165 34912 32000 34914
rect 28165 34856 28170 34912
rect 28226 34856 32000 34912
rect 28165 34854 32000 34856
rect 28165 34851 28231 34854
rect 20805 34848 21125 34849
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 31200 34824 32000 34854
rect 20805 34783 21125 34784
rect 1577 34642 1643 34645
rect 0 34640 1643 34642
rect 0 34584 1582 34640
rect 1638 34584 1643 34640
rect 0 34582 1643 34584
rect 0 34552 800 34582
rect 1577 34579 1643 34582
rect 19701 34640 19810 34645
rect 19701 34584 19706 34640
rect 19762 34584 19810 34640
rect 19701 34582 19810 34584
rect 19701 34579 19767 34582
rect 28901 34506 28967 34509
rect 31200 34506 32000 34536
rect 28901 34504 32000 34506
rect 28901 34448 28906 34504
rect 28962 34448 32000 34504
rect 28901 34446 32000 34448
rect 28901 34443 28967 34446
rect 31200 34416 32000 34446
rect 5909 34304 6229 34305
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6229 34304
rect 5909 34239 6229 34240
rect 15840 34304 16160 34305
rect 15840 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15840 34239 16160 34240
rect 25770 34304 26090 34305
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26090 34304
rect 25770 34239 26090 34240
rect 30097 34234 30163 34237
rect 30230 34234 30236 34236
rect 30097 34232 30236 34234
rect 30097 34176 30102 34232
rect 30158 34176 30236 34232
rect 30097 34174 30236 34176
rect 30097 34171 30163 34174
rect 30230 34172 30236 34174
rect 30300 34172 30306 34236
rect 17350 34036 17356 34100
rect 17420 34098 17426 34100
rect 25773 34098 25839 34101
rect 17420 34096 25839 34098
rect 17420 34040 25778 34096
rect 25834 34040 25839 34096
rect 17420 34038 25839 34040
rect 17420 34036 17426 34038
rect 25773 34035 25839 34038
rect 30005 34098 30071 34101
rect 31200 34098 32000 34128
rect 30005 34096 32000 34098
rect 30005 34040 30010 34096
rect 30066 34040 32000 34096
rect 30005 34038 32000 34040
rect 30005 34035 30071 34038
rect 31200 34008 32000 34038
rect 0 33962 800 33992
rect 1393 33962 1459 33965
rect 0 33960 1459 33962
rect 0 33904 1398 33960
rect 1454 33904 1459 33960
rect 0 33902 1459 33904
rect 0 33872 800 33902
rect 1393 33899 1459 33902
rect 24209 33826 24275 33829
rect 24342 33826 24348 33828
rect 24209 33824 24348 33826
rect 24209 33768 24214 33824
rect 24270 33768 24348 33824
rect 24209 33766 24348 33768
rect 24209 33763 24275 33766
rect 24342 33764 24348 33766
rect 24412 33764 24418 33828
rect 10874 33760 11194 33761
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 33695 11194 33696
rect 20805 33760 21125 33761
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 33695 21125 33696
rect 27153 33556 27219 33557
rect 27102 33554 27108 33556
rect 27062 33494 27108 33554
rect 27172 33552 27219 33556
rect 27214 33496 27219 33552
rect 27102 33492 27108 33494
rect 27172 33492 27219 33496
rect 27153 33491 27219 33492
rect 28901 33554 28967 33557
rect 31200 33554 32000 33584
rect 28901 33552 32000 33554
rect 28901 33496 28906 33552
rect 28962 33496 32000 33552
rect 28901 33494 32000 33496
rect 28901 33491 28967 33494
rect 31200 33464 32000 33494
rect 0 33282 800 33312
rect 1577 33282 1643 33285
rect 0 33280 1643 33282
rect 0 33224 1582 33280
rect 1638 33224 1643 33280
rect 0 33222 1643 33224
rect 0 33192 800 33222
rect 1577 33219 1643 33222
rect 5909 33216 6229 33217
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6229 33216
rect 5909 33151 6229 33152
rect 15840 33216 16160 33217
rect 15840 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15840 33151 16160 33152
rect 25770 33216 26090 33217
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26090 33216
rect 25770 33151 26090 33152
rect 29269 33146 29335 33149
rect 31200 33146 32000 33176
rect 29269 33144 32000 33146
rect 29269 33088 29274 33144
rect 29330 33088 32000 33144
rect 29269 33086 32000 33088
rect 29269 33083 29335 33086
rect 31200 33056 32000 33086
rect 25630 32948 25636 33012
rect 25700 33010 25706 33012
rect 25773 33010 25839 33013
rect 25700 33008 25839 33010
rect 25700 32952 25778 33008
rect 25834 32952 25839 33008
rect 25700 32950 25839 32952
rect 25700 32948 25706 32950
rect 25773 32947 25839 32950
rect 21265 32874 21331 32877
rect 22921 32874 22987 32877
rect 21265 32872 22987 32874
rect 21265 32816 21270 32872
rect 21326 32816 22926 32872
rect 22982 32816 22987 32872
rect 21265 32814 22987 32816
rect 21265 32811 21331 32814
rect 22921 32811 22987 32814
rect 25405 32874 25471 32877
rect 25630 32874 25636 32876
rect 25405 32872 25636 32874
rect 25405 32816 25410 32872
rect 25466 32816 25636 32872
rect 25405 32814 25636 32816
rect 25405 32811 25471 32814
rect 25630 32812 25636 32814
rect 25700 32812 25706 32876
rect 29126 32874 29132 32876
rect 28720 32814 29132 32874
rect 0 32738 800 32768
rect 28720 32741 28780 32814
rect 29126 32812 29132 32814
rect 29196 32812 29202 32876
rect 1393 32738 1459 32741
rect 0 32736 1459 32738
rect 0 32680 1398 32736
rect 1454 32680 1459 32736
rect 0 32678 1459 32680
rect 0 32648 800 32678
rect 1393 32675 1459 32678
rect 28073 32738 28139 32741
rect 28073 32736 28274 32738
rect 28073 32680 28078 32736
rect 28134 32680 28274 32736
rect 28073 32678 28274 32680
rect 28073 32675 28139 32678
rect 10874 32672 11194 32673
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 32607 11194 32608
rect 20805 32672 21125 32673
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 20805 32607 21125 32608
rect 26182 32540 26188 32604
rect 26252 32602 26258 32604
rect 26918 32602 26924 32604
rect 26252 32542 26924 32602
rect 26252 32540 26258 32542
rect 26918 32540 26924 32542
rect 26988 32602 26994 32604
rect 28073 32602 28139 32605
rect 26988 32600 28139 32602
rect 26988 32544 28078 32600
rect 28134 32544 28139 32600
rect 26988 32542 28139 32544
rect 26988 32540 26994 32542
rect 28073 32539 28139 32542
rect 26918 32404 26924 32468
rect 26988 32466 26994 32468
rect 27613 32466 27679 32469
rect 28214 32466 28274 32678
rect 28717 32736 28783 32741
rect 28717 32680 28722 32736
rect 28778 32680 28783 32736
rect 28717 32675 28783 32680
rect 29126 32676 29132 32740
rect 29196 32738 29202 32740
rect 29913 32738 29979 32741
rect 29196 32736 29979 32738
rect 29196 32680 29918 32736
rect 29974 32680 29979 32736
rect 29196 32678 29979 32680
rect 29196 32676 29202 32678
rect 29913 32675 29979 32678
rect 28809 32600 28875 32605
rect 28809 32544 28814 32600
rect 28870 32544 28875 32600
rect 28809 32539 28875 32544
rect 28993 32600 29059 32605
rect 28993 32544 28998 32600
rect 29054 32544 29059 32600
rect 28993 32539 29059 32544
rect 30005 32602 30071 32605
rect 31200 32602 32000 32632
rect 30005 32600 32000 32602
rect 30005 32544 30010 32600
rect 30066 32544 32000 32600
rect 30005 32542 32000 32544
rect 30005 32539 30071 32542
rect 26988 32464 27679 32466
rect 26988 32408 27618 32464
rect 27674 32408 27679 32464
rect 26988 32406 27679 32408
rect 26988 32404 26994 32406
rect 27613 32403 27679 32406
rect 28076 32406 28274 32466
rect 28076 32333 28136 32406
rect 27286 32268 27292 32332
rect 27356 32330 27362 32332
rect 27705 32330 27771 32333
rect 27356 32328 27771 32330
rect 27356 32272 27710 32328
rect 27766 32272 27771 32328
rect 27356 32270 27771 32272
rect 27356 32268 27362 32270
rect 27705 32267 27771 32270
rect 28073 32328 28139 32333
rect 28812 32330 28872 32539
rect 28073 32272 28078 32328
rect 28134 32272 28139 32328
rect 28073 32267 28139 32272
rect 28214 32270 28872 32330
rect 28996 32330 29056 32539
rect 31200 32512 32000 32542
rect 29177 32330 29243 32333
rect 28996 32328 29243 32330
rect 28996 32272 29182 32328
rect 29238 32272 29243 32328
rect 28996 32270 29243 32272
rect 23197 32196 23263 32197
rect 23197 32194 23244 32196
rect 23152 32192 23244 32194
rect 23152 32136 23202 32192
rect 23152 32134 23244 32136
rect 23197 32132 23244 32134
rect 23308 32132 23314 32196
rect 26550 32132 26556 32196
rect 26620 32194 26626 32196
rect 26969 32194 27035 32197
rect 27654 32194 27660 32196
rect 26620 32192 27035 32194
rect 26620 32136 26974 32192
rect 27030 32136 27035 32192
rect 26620 32134 27035 32136
rect 26620 32132 26626 32134
rect 23197 32131 23263 32132
rect 26969 32131 27035 32134
rect 27478 32134 27660 32194
rect 5909 32128 6229 32129
rect 0 32058 800 32088
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6229 32128
rect 5909 32063 6229 32064
rect 15840 32128 16160 32129
rect 15840 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 15840 32063 16160 32064
rect 25770 32128 26090 32129
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26090 32128
rect 25770 32063 26090 32064
rect 1485 32058 1551 32061
rect 0 32056 1551 32058
rect 0 32000 1490 32056
rect 1546 32000 1551 32056
rect 0 31998 1551 32000
rect 0 31968 800 31998
rect 1485 31995 1551 31998
rect 24710 31996 24716 32060
rect 24780 32058 24786 32060
rect 25129 32058 25195 32061
rect 24780 32056 25195 32058
rect 24780 32000 25134 32056
rect 25190 32000 25195 32056
rect 24780 31998 25195 32000
rect 24780 31996 24786 31998
rect 25129 31995 25195 31998
rect 1853 31922 1919 31925
rect 26049 31922 26115 31925
rect 1853 31920 26115 31922
rect 1853 31864 1858 31920
rect 1914 31864 26054 31920
rect 26110 31864 26115 31920
rect 1853 31862 26115 31864
rect 1853 31859 1919 31862
rect 26049 31859 26115 31862
rect 23381 31770 23447 31773
rect 23246 31768 23447 31770
rect 23246 31712 23386 31768
rect 23442 31712 23447 31768
rect 25262 31724 25268 31788
rect 25332 31786 25338 31788
rect 25589 31786 25655 31789
rect 25332 31784 25655 31786
rect 25332 31728 25594 31784
rect 25650 31728 25655 31784
rect 25332 31726 25655 31728
rect 25332 31724 25338 31726
rect 25589 31723 25655 31726
rect 26969 31786 27035 31789
rect 27102 31786 27108 31788
rect 26969 31784 27108 31786
rect 26969 31728 26974 31784
rect 27030 31728 27108 31784
rect 26969 31726 27108 31728
rect 26969 31723 27035 31726
rect 27102 31724 27108 31726
rect 27172 31724 27178 31788
rect 27478 31786 27538 32134
rect 27654 32132 27660 32134
rect 27724 32132 27730 32196
rect 27705 32060 27771 32061
rect 27654 31996 27660 32060
rect 27724 32058 27771 32060
rect 28214 32058 28274 32270
rect 29177 32267 29243 32270
rect 29361 32330 29427 32333
rect 30966 32330 30972 32332
rect 29361 32328 30972 32330
rect 29361 32272 29366 32328
rect 29422 32272 30972 32328
rect 29361 32270 30972 32272
rect 29361 32267 29427 32270
rect 30966 32268 30972 32270
rect 31036 32268 31042 32332
rect 28901 32194 28967 32197
rect 31200 32194 32000 32224
rect 28901 32192 32000 32194
rect 28901 32136 28906 32192
rect 28962 32136 32000 32192
rect 28901 32134 32000 32136
rect 28901 32131 28967 32134
rect 31200 32104 32000 32134
rect 27724 32056 27816 32058
rect 27766 32000 27816 32056
rect 27724 31998 27816 32000
rect 28076 31998 28274 32058
rect 28625 32058 28691 32061
rect 28993 32058 29059 32061
rect 28625 32056 29059 32058
rect 28625 32000 28630 32056
rect 28686 32000 28998 32056
rect 29054 32000 29059 32056
rect 28625 31998 29059 32000
rect 27724 31996 27771 31998
rect 27705 31995 27771 31996
rect 28076 31789 28136 31998
rect 28625 31995 28691 31998
rect 28993 31995 29059 31998
rect 30833 32056 30899 32061
rect 30833 32000 30838 32056
rect 30894 32000 30899 32056
rect 30833 31995 30899 32000
rect 28206 31860 28212 31924
rect 28276 31922 28282 31924
rect 28993 31922 29059 31925
rect 28276 31920 29059 31922
rect 28276 31864 28998 31920
rect 29054 31864 29059 31920
rect 28276 31862 29059 31864
rect 28276 31860 28282 31862
rect 28993 31859 29059 31862
rect 30097 31922 30163 31925
rect 30414 31922 30420 31924
rect 30097 31920 30420 31922
rect 30097 31864 30102 31920
rect 30158 31864 30420 31920
rect 30097 31862 30420 31864
rect 30097 31859 30163 31862
rect 30414 31860 30420 31862
rect 30484 31860 30490 31924
rect 27613 31786 27679 31789
rect 27478 31784 27679 31786
rect 27478 31728 27618 31784
rect 27674 31728 27679 31784
rect 27478 31726 27679 31728
rect 27613 31723 27679 31726
rect 28073 31784 28139 31789
rect 28073 31728 28078 31784
rect 28134 31728 28139 31784
rect 28073 31723 28139 31728
rect 29729 31786 29795 31789
rect 30598 31786 30604 31788
rect 29729 31784 30604 31786
rect 29729 31728 29734 31784
rect 29790 31728 30604 31784
rect 29729 31726 30604 31728
rect 29729 31723 29795 31726
rect 30598 31724 30604 31726
rect 30668 31724 30674 31788
rect 23246 31710 23447 31712
rect 23246 31650 23306 31710
rect 23381 31707 23447 31710
rect 23062 31590 23306 31650
rect 26233 31650 26299 31653
rect 26366 31650 26372 31652
rect 26233 31648 26372 31650
rect 26233 31592 26238 31648
rect 26294 31592 26372 31648
rect 26233 31590 26372 31592
rect 10874 31584 11194 31585
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 31519 11194 31520
rect 20805 31584 21125 31585
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 20805 31519 21125 31520
rect 22921 31514 22987 31517
rect 23062 31514 23122 31590
rect 26233 31587 26299 31590
rect 26366 31588 26372 31590
rect 26436 31588 26442 31652
rect 30836 31650 30896 31995
rect 31150 31860 31156 31924
rect 31220 31922 31226 31924
rect 31753 31922 31819 31925
rect 31220 31920 31819 31922
rect 31220 31864 31758 31920
rect 31814 31864 31819 31920
rect 31220 31862 31819 31864
rect 31220 31860 31226 31862
rect 31753 31859 31819 31862
rect 31200 31650 32000 31680
rect 30836 31590 32000 31650
rect 31200 31560 32000 31590
rect 23289 31516 23355 31517
rect 23238 31514 23244 31516
rect 22921 31512 23122 31514
rect 22921 31456 22926 31512
rect 22982 31456 23122 31512
rect 22921 31454 23122 31456
rect 23198 31454 23244 31514
rect 23308 31512 23355 31516
rect 23350 31456 23355 31512
rect 22921 31451 22987 31454
rect 23238 31452 23244 31454
rect 23308 31452 23355 31456
rect 27654 31452 27660 31516
rect 27724 31514 27730 31516
rect 28441 31514 28507 31517
rect 27724 31512 28507 31514
rect 27724 31456 28446 31512
rect 28502 31456 28507 31512
rect 27724 31454 28507 31456
rect 27724 31452 27730 31454
rect 23289 31451 23355 31452
rect 28441 31451 28507 31454
rect 0 31378 800 31408
rect 1577 31378 1643 31381
rect 0 31376 1643 31378
rect 0 31320 1582 31376
rect 1638 31320 1643 31376
rect 0 31318 1643 31320
rect 0 31288 800 31318
rect 1577 31315 1643 31318
rect 24853 31378 24919 31381
rect 25078 31378 25084 31380
rect 24853 31376 25084 31378
rect 24853 31320 24858 31376
rect 24914 31320 25084 31376
rect 24853 31318 25084 31320
rect 24853 31315 24919 31318
rect 25078 31316 25084 31318
rect 25148 31316 25154 31380
rect 26141 31378 26207 31381
rect 26141 31376 26250 31378
rect 26141 31320 26146 31376
rect 26202 31320 26250 31376
rect 26141 31315 26250 31320
rect 27654 31316 27660 31380
rect 27724 31378 27730 31380
rect 28073 31378 28139 31381
rect 27724 31376 28139 31378
rect 27724 31320 28078 31376
rect 28134 31320 28139 31376
rect 27724 31318 28139 31320
rect 27724 31316 27730 31318
rect 28073 31315 28139 31318
rect 29545 31378 29611 31381
rect 30414 31378 30420 31380
rect 29545 31376 30420 31378
rect 29545 31320 29550 31376
rect 29606 31320 30420 31376
rect 29545 31318 30420 31320
rect 29545 31315 29611 31318
rect 30414 31316 30420 31318
rect 30484 31316 30490 31380
rect 25129 31242 25195 31245
rect 25446 31242 25452 31244
rect 25129 31240 25452 31242
rect 25129 31184 25134 31240
rect 25190 31184 25452 31240
rect 25129 31182 25452 31184
rect 25129 31179 25195 31182
rect 25446 31180 25452 31182
rect 25516 31180 25522 31244
rect 5909 31040 6229 31041
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6229 31040
rect 5909 30975 6229 30976
rect 15840 31040 16160 31041
rect 15840 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15840 30975 16160 30976
rect 25770 31040 26090 31041
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26090 31040
rect 25770 30975 26090 30976
rect 26049 30834 26115 30837
rect 26190 30834 26250 31315
rect 30557 31242 30623 31245
rect 31200 31242 32000 31272
rect 30557 31240 32000 31242
rect 30557 31184 30562 31240
rect 30618 31184 32000 31240
rect 30557 31182 32000 31184
rect 30557 31179 30623 31182
rect 31200 31152 32000 31182
rect 27470 31106 27476 31108
rect 26049 30832 26250 30834
rect 26049 30776 26054 30832
rect 26110 30776 26250 30832
rect 26049 30774 26250 30776
rect 27340 31046 27476 31106
rect 27340 30834 27400 31046
rect 27470 31044 27476 31046
rect 27540 31044 27546 31108
rect 30281 31106 30347 31109
rect 30598 31106 30604 31108
rect 30281 31104 30604 31106
rect 30281 31048 30286 31104
rect 30342 31048 30604 31104
rect 30281 31046 30604 31048
rect 30281 31043 30347 31046
rect 30598 31044 30604 31046
rect 30668 31044 30674 31108
rect 27521 30972 27587 30973
rect 27470 30908 27476 30972
rect 27540 30970 27587 30972
rect 27540 30968 27632 30970
rect 27582 30912 27632 30968
rect 27540 30910 27632 30912
rect 27540 30908 27587 30910
rect 28942 30908 28948 30972
rect 29012 30970 29018 30972
rect 30557 30970 30623 30973
rect 29012 30968 30623 30970
rect 29012 30912 30562 30968
rect 30618 30912 30623 30968
rect 29012 30910 30623 30912
rect 29012 30908 29018 30910
rect 27521 30907 27587 30908
rect 30557 30907 30623 30910
rect 31150 30908 31156 30972
rect 31220 30970 31226 30972
rect 31477 30970 31543 30973
rect 31220 30968 31543 30970
rect 31220 30912 31482 30968
rect 31538 30912 31543 30968
rect 31220 30910 31543 30912
rect 31220 30908 31226 30910
rect 31477 30907 31543 30910
rect 27521 30834 27587 30837
rect 27340 30832 27587 30834
rect 27340 30776 27526 30832
rect 27582 30776 27587 30832
rect 27340 30774 27587 30776
rect 26049 30771 26115 30774
rect 27521 30771 27587 30774
rect 28809 30834 28875 30837
rect 28942 30834 28948 30836
rect 28809 30832 28948 30834
rect 28809 30776 28814 30832
rect 28870 30776 28948 30832
rect 28809 30774 28948 30776
rect 28809 30771 28875 30774
rect 28942 30772 28948 30774
rect 29012 30772 29018 30836
rect 30373 30834 30439 30837
rect 29870 30832 30439 30834
rect 29870 30776 30378 30832
rect 30434 30776 30439 30832
rect 29870 30774 30439 30776
rect 0 30698 800 30728
rect 1577 30698 1643 30701
rect 0 30696 1643 30698
rect 0 30640 1582 30696
rect 1638 30640 1643 30696
rect 0 30638 1643 30640
rect 0 30608 800 30638
rect 1577 30635 1643 30638
rect 25037 30698 25103 30701
rect 25262 30698 25268 30700
rect 25037 30696 25268 30698
rect 25037 30640 25042 30696
rect 25098 30640 25268 30696
rect 25037 30638 25268 30640
rect 25037 30635 25103 30638
rect 25262 30636 25268 30638
rect 25332 30636 25338 30700
rect 29545 30562 29611 30565
rect 29870 30562 29930 30774
rect 30373 30771 30439 30774
rect 30097 30698 30163 30701
rect 31200 30698 32000 30728
rect 30097 30696 32000 30698
rect 30097 30640 30102 30696
rect 30158 30640 32000 30696
rect 30097 30638 32000 30640
rect 30097 30635 30163 30638
rect 31200 30608 32000 30638
rect 29545 30560 29930 30562
rect 29545 30504 29550 30560
rect 29606 30504 29930 30560
rect 29545 30502 29930 30504
rect 29545 30499 29611 30502
rect 10874 30496 11194 30497
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 10874 30431 11194 30432
rect 20805 30496 21125 30497
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 20805 30431 21125 30432
rect 26366 30364 26372 30428
rect 26436 30426 26442 30428
rect 26785 30426 26851 30429
rect 26436 30424 26851 30426
rect 26436 30368 26790 30424
rect 26846 30368 26851 30424
rect 26436 30366 26851 30368
rect 26436 30364 26442 30366
rect 26785 30363 26851 30366
rect 28901 30426 28967 30429
rect 30782 30426 30788 30428
rect 28901 30424 30788 30426
rect 28901 30368 28906 30424
rect 28962 30368 30788 30424
rect 28901 30366 30788 30368
rect 28901 30363 28967 30366
rect 30782 30364 30788 30366
rect 30852 30364 30858 30428
rect 24158 30228 24164 30292
rect 24228 30290 24234 30292
rect 30005 30290 30071 30293
rect 31200 30290 32000 30320
rect 24228 30230 28090 30290
rect 24228 30228 24234 30230
rect 25262 30092 25268 30156
rect 25332 30154 25338 30156
rect 25589 30154 25655 30157
rect 25332 30152 25655 30154
rect 25332 30096 25594 30152
rect 25650 30096 25655 30152
rect 25332 30094 25655 30096
rect 25332 30092 25338 30094
rect 25589 30091 25655 30094
rect 26182 30092 26188 30156
rect 26252 30154 26258 30156
rect 26252 30094 27630 30154
rect 26252 30092 26258 30094
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 27337 30018 27403 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 27294 30016 27403 30018
rect 27294 29960 27342 30016
rect 27398 29960 27403 30016
rect 27294 29955 27403 29960
rect 5909 29952 6229 29953
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6229 29952
rect 5909 29887 6229 29888
rect 15840 29952 16160 29953
rect 15840 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15840 29887 16160 29888
rect 25770 29952 26090 29953
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26090 29952
rect 25770 29887 26090 29888
rect 22093 29884 22159 29885
rect 27061 29884 27127 29885
rect 22093 29880 22140 29884
rect 22204 29882 22210 29884
rect 27061 29882 27108 29884
rect 22093 29824 22098 29880
rect 22093 29820 22140 29824
rect 22204 29822 22250 29882
rect 27016 29880 27108 29882
rect 27016 29824 27066 29880
rect 27016 29822 27108 29824
rect 22204 29820 22210 29822
rect 27061 29820 27108 29822
rect 27172 29820 27178 29884
rect 22093 29819 22159 29820
rect 27061 29819 27127 29820
rect 24894 29684 24900 29748
rect 24964 29746 24970 29748
rect 25773 29746 25839 29749
rect 26785 29748 26851 29749
rect 24964 29744 25839 29746
rect 24964 29688 25778 29744
rect 25834 29688 25839 29744
rect 24964 29686 25839 29688
rect 24964 29684 24970 29686
rect 25773 29683 25839 29686
rect 26734 29684 26740 29748
rect 26804 29746 26851 29748
rect 26804 29744 26896 29746
rect 26846 29688 26896 29744
rect 26804 29686 26896 29688
rect 26804 29684 26851 29686
rect 26785 29683 26851 29684
rect 26734 29548 26740 29612
rect 26804 29610 26810 29612
rect 27294 29610 27354 29955
rect 26804 29550 27354 29610
rect 27570 29610 27630 30094
rect 28030 29746 28090 30230
rect 30005 30288 32000 30290
rect 30005 30232 30010 30288
rect 30066 30232 32000 30288
rect 30005 30230 32000 30232
rect 30005 30227 30071 30230
rect 31200 30200 32000 30230
rect 28257 30018 28323 30021
rect 30598 30018 30604 30020
rect 28257 30016 30604 30018
rect 28257 29960 28262 30016
rect 28318 29960 30604 30016
rect 28257 29958 30604 29960
rect 28257 29955 28323 29958
rect 30598 29956 30604 29958
rect 30668 29956 30674 30020
rect 28206 29820 28212 29884
rect 28276 29882 28282 29884
rect 29545 29882 29611 29885
rect 28276 29880 29611 29882
rect 28276 29824 29550 29880
rect 29606 29824 29611 29880
rect 28276 29822 29611 29824
rect 28276 29820 28282 29822
rect 29545 29819 29611 29822
rect 28349 29746 28415 29749
rect 31200 29746 32000 29776
rect 28030 29686 28136 29746
rect 27889 29610 27955 29613
rect 27570 29608 27955 29610
rect 27570 29552 27894 29608
rect 27950 29552 27955 29608
rect 27570 29550 27955 29552
rect 26804 29548 26810 29550
rect 27889 29547 27955 29550
rect 28076 29477 28136 29686
rect 28349 29744 32000 29746
rect 28349 29688 28354 29744
rect 28410 29688 32000 29744
rect 28349 29686 32000 29688
rect 28349 29683 28415 29686
rect 31200 29656 32000 29686
rect 25957 29474 26023 29477
rect 25957 29472 27952 29474
rect 25957 29416 25962 29472
rect 26018 29416 27952 29472
rect 25957 29414 27952 29416
rect 25957 29411 26023 29414
rect 10874 29408 11194 29409
rect 0 29338 800 29368
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 29343 11194 29344
rect 20805 29408 21125 29409
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 29343 21125 29344
rect 1577 29338 1643 29341
rect 0 29336 1643 29338
rect 0 29280 1582 29336
rect 1638 29280 1643 29336
rect 0 29278 1643 29280
rect 0 29248 800 29278
rect 1577 29275 1643 29278
rect 26049 29338 26115 29341
rect 26182 29338 26188 29340
rect 26049 29336 26188 29338
rect 26049 29280 26054 29336
rect 26110 29280 26188 29336
rect 26049 29278 26188 29280
rect 26049 29275 26115 29278
rect 26182 29276 26188 29278
rect 26252 29276 26258 29340
rect 27521 29336 27587 29341
rect 27521 29280 27526 29336
rect 27582 29304 27587 29336
rect 27892 29338 27952 29414
rect 28073 29472 28139 29477
rect 28073 29416 28078 29472
rect 28134 29416 28139 29472
rect 28073 29411 28139 29416
rect 31200 29338 32000 29368
rect 27582 29280 27630 29304
rect 27521 29275 27630 29280
rect 27892 29278 32000 29338
rect 27524 29244 27630 29275
rect 31200 29248 32000 29278
rect 19609 29202 19675 29205
rect 26049 29202 26115 29205
rect 27286 29202 27292 29204
rect 19609 29200 27292 29202
rect 19609 29144 19614 29200
rect 19670 29144 26054 29200
rect 26110 29144 27292 29200
rect 19609 29142 27292 29144
rect 19609 29139 19675 29142
rect 26049 29139 26115 29142
rect 27286 29140 27292 29142
rect 27356 29140 27362 29204
rect 27570 29202 27630 29244
rect 28165 29202 28231 29205
rect 27570 29200 28231 29202
rect 27570 29144 28170 29200
rect 28226 29144 28231 29200
rect 27570 29142 28231 29144
rect 28165 29139 28231 29142
rect 12617 29066 12683 29069
rect 12801 29066 12867 29069
rect 19057 29066 19123 29069
rect 12617 29064 19123 29066
rect 12617 29008 12622 29064
rect 12678 29008 12806 29064
rect 12862 29008 19062 29064
rect 19118 29008 19123 29064
rect 12617 29006 19123 29008
rect 12617 29003 12683 29006
rect 12801 29003 12867 29006
rect 19057 29003 19123 29006
rect 27245 29066 27311 29069
rect 29453 29066 29519 29069
rect 27245 29064 29519 29066
rect 27245 29008 27250 29064
rect 27306 29008 29458 29064
rect 29514 29008 29519 29064
rect 27245 29006 29519 29008
rect 27245 29003 27311 29006
rect 29453 29003 29519 29006
rect 27889 28930 27955 28933
rect 28022 28930 28028 28932
rect 27889 28928 28028 28930
rect 27889 28872 27894 28928
rect 27950 28872 28028 28928
rect 27889 28870 28028 28872
rect 27889 28867 27955 28870
rect 28022 28868 28028 28870
rect 28092 28868 28098 28932
rect 5909 28864 6229 28865
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6229 28864
rect 5909 28799 6229 28800
rect 15840 28864 16160 28865
rect 15840 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15840 28799 16160 28800
rect 25770 28864 26090 28865
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26090 28864
rect 25770 28799 26090 28800
rect 13629 28794 13695 28797
rect 14733 28794 14799 28797
rect 13629 28792 14799 28794
rect 13629 28736 13634 28792
rect 13690 28736 14738 28792
rect 14794 28736 14799 28792
rect 13629 28734 14799 28736
rect 13629 28731 13695 28734
rect 14733 28731 14799 28734
rect 27521 28794 27587 28797
rect 30005 28794 30071 28797
rect 27521 28792 30071 28794
rect 27521 28736 27526 28792
rect 27582 28736 30010 28792
rect 30066 28736 30071 28792
rect 27521 28734 30071 28736
rect 27521 28731 27587 28734
rect 30005 28731 30071 28734
rect 30598 28732 30604 28796
rect 30668 28794 30674 28796
rect 31200 28794 32000 28824
rect 30668 28734 32000 28794
rect 30668 28732 30674 28734
rect 31200 28704 32000 28734
rect 0 28658 800 28688
rect 1577 28658 1643 28661
rect 0 28656 1643 28658
rect 0 28600 1582 28656
rect 1638 28600 1643 28656
rect 0 28598 1643 28600
rect 0 28568 800 28598
rect 1577 28595 1643 28598
rect 25037 28660 25103 28661
rect 25037 28656 25084 28660
rect 25148 28658 25154 28660
rect 25037 28600 25042 28656
rect 25037 28596 25084 28600
rect 25148 28598 25194 28658
rect 25148 28596 25154 28598
rect 25037 28595 25103 28596
rect 28901 28520 28967 28525
rect 28901 28464 28906 28520
rect 28962 28464 28967 28520
rect 28901 28459 28967 28464
rect 28904 28386 28964 28459
rect 31200 28386 32000 28416
rect 28904 28326 32000 28386
rect 10874 28320 11194 28321
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 28255 11194 28256
rect 20805 28320 21125 28321
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 31200 28296 32000 28326
rect 20805 28255 21125 28256
rect 14365 28250 14431 28253
rect 15510 28250 15516 28252
rect 14365 28248 15516 28250
rect 14365 28192 14370 28248
rect 14426 28192 15516 28248
rect 14365 28190 15516 28192
rect 14365 28187 14431 28190
rect 15510 28188 15516 28190
rect 15580 28250 15586 28252
rect 15837 28250 15903 28253
rect 15580 28248 15903 28250
rect 15580 28192 15842 28248
rect 15898 28192 15903 28248
rect 15580 28190 15903 28192
rect 15580 28188 15586 28190
rect 15837 28187 15903 28190
rect 0 28114 800 28144
rect 1577 28114 1643 28117
rect 15745 28114 15811 28117
rect 0 28112 1643 28114
rect 0 28056 1582 28112
rect 1638 28056 1643 28112
rect 0 28054 1643 28056
rect 0 28024 800 28054
rect 1577 28051 1643 28054
rect 15334 28112 15811 28114
rect 15334 28056 15750 28112
rect 15806 28056 15811 28112
rect 15334 28054 15811 28056
rect 5909 27776 6229 27777
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6229 27776
rect 5909 27711 6229 27712
rect 15334 27573 15394 28054
rect 15745 28051 15811 28054
rect 19190 28052 19196 28116
rect 19260 28114 19266 28116
rect 29361 28114 29427 28117
rect 19260 28112 29427 28114
rect 19260 28056 29366 28112
rect 29422 28056 29427 28112
rect 19260 28054 29427 28056
rect 19260 28052 19266 28054
rect 29361 28051 29427 28054
rect 25446 27916 25452 27980
rect 25516 27978 25522 27980
rect 25589 27978 25655 27981
rect 25516 27976 25655 27978
rect 25516 27920 25594 27976
rect 25650 27920 25655 27976
rect 25516 27918 25655 27920
rect 25516 27916 25522 27918
rect 25589 27915 25655 27918
rect 26366 27916 26372 27980
rect 26436 27978 26442 27980
rect 27245 27978 27311 27981
rect 26436 27976 27311 27978
rect 26436 27920 27250 27976
rect 27306 27920 27311 27976
rect 26436 27918 27311 27920
rect 26436 27916 26442 27918
rect 27245 27915 27311 27918
rect 27705 27978 27771 27981
rect 31200 27978 32000 28008
rect 27705 27976 32000 27978
rect 27705 27920 27710 27976
rect 27766 27920 32000 27976
rect 27705 27918 32000 27920
rect 27705 27915 27771 27918
rect 31200 27888 32000 27918
rect 15469 27844 15535 27845
rect 15469 27840 15516 27844
rect 15580 27842 15586 27844
rect 28993 27842 29059 27845
rect 29126 27842 29132 27844
rect 15469 27784 15474 27840
rect 15469 27780 15516 27784
rect 15580 27782 15626 27842
rect 28993 27840 29132 27842
rect 28993 27784 28998 27840
rect 29054 27784 29132 27840
rect 28993 27782 29132 27784
rect 15580 27780 15586 27782
rect 15469 27779 15535 27780
rect 28993 27779 29059 27782
rect 29126 27780 29132 27782
rect 29196 27780 29202 27844
rect 15840 27776 16160 27777
rect 15840 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15840 27711 16160 27712
rect 25770 27776 26090 27777
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26090 27776
rect 25770 27711 26090 27712
rect 15334 27568 15443 27573
rect 15334 27512 15382 27568
rect 15438 27512 15443 27568
rect 15334 27510 15443 27512
rect 15377 27507 15443 27510
rect 17534 27508 17540 27572
rect 17604 27570 17610 27572
rect 27705 27570 27771 27573
rect 17604 27568 27771 27570
rect 17604 27512 27710 27568
rect 27766 27512 27771 27568
rect 17604 27510 27771 27512
rect 17604 27508 17610 27510
rect 27705 27507 27771 27510
rect 0 27434 800 27464
rect 1577 27434 1643 27437
rect 0 27432 1643 27434
rect 0 27376 1582 27432
rect 1638 27376 1643 27432
rect 0 27374 1643 27376
rect 0 27344 800 27374
rect 1577 27371 1643 27374
rect 26918 27372 26924 27436
rect 26988 27434 26994 27436
rect 27705 27434 27771 27437
rect 26988 27432 27771 27434
rect 26988 27376 27710 27432
rect 27766 27376 27771 27432
rect 26988 27374 27771 27376
rect 26988 27372 26994 27374
rect 27705 27371 27771 27374
rect 28441 27432 28507 27437
rect 28441 27376 28446 27432
rect 28502 27376 28507 27432
rect 28441 27371 28507 27376
rect 28625 27434 28691 27437
rect 31200 27434 32000 27464
rect 28625 27432 32000 27434
rect 28625 27376 28630 27432
rect 28686 27376 32000 27432
rect 28625 27374 32000 27376
rect 28625 27371 28691 27374
rect 26366 27236 26372 27300
rect 26436 27298 26442 27300
rect 28444 27298 28504 27371
rect 31200 27344 32000 27374
rect 26436 27238 28504 27298
rect 26436 27236 26442 27238
rect 10874 27232 11194 27233
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 10874 27167 11194 27168
rect 20805 27232 21125 27233
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 27167 21125 27168
rect 25405 27164 25471 27165
rect 25405 27162 25452 27164
rect 25360 27160 25452 27162
rect 25360 27104 25410 27160
rect 25360 27102 25452 27104
rect 25405 27100 25452 27102
rect 25516 27100 25522 27164
rect 25405 27099 25471 27100
rect 16205 27026 16271 27029
rect 25681 27026 25747 27029
rect 16205 27024 16314 27026
rect 16205 26968 16210 27024
rect 16266 26968 16314 27024
rect 16205 26963 16314 26968
rect 0 26754 800 26784
rect 16254 26757 16314 26963
rect 25270 27024 25747 27026
rect 25270 26968 25686 27024
rect 25742 26968 25747 27024
rect 25270 26966 25747 26968
rect 25129 26890 25195 26893
rect 25270 26890 25330 26966
rect 25681 26963 25747 26966
rect 27153 27026 27219 27029
rect 27286 27026 27292 27028
rect 27153 27024 27292 27026
rect 27153 26968 27158 27024
rect 27214 26968 27292 27024
rect 27153 26966 27292 26968
rect 27153 26963 27219 26966
rect 27286 26964 27292 26966
rect 27356 26964 27362 27028
rect 30005 27026 30071 27029
rect 31200 27026 32000 27056
rect 30005 27024 32000 27026
rect 30005 26968 30010 27024
rect 30066 26968 32000 27024
rect 30005 26966 32000 26968
rect 30005 26963 30071 26966
rect 31200 26936 32000 26966
rect 25129 26888 25330 26890
rect 25129 26832 25134 26888
rect 25190 26832 25330 26888
rect 25129 26830 25330 26832
rect 25129 26827 25195 26830
rect 25630 26828 25636 26892
rect 25700 26890 25706 26892
rect 27245 26890 27311 26893
rect 25700 26888 27311 26890
rect 25700 26832 27250 26888
rect 27306 26832 27311 26888
rect 25700 26830 27311 26832
rect 25700 26828 25706 26830
rect 27245 26827 27311 26830
rect 1577 26754 1643 26757
rect 0 26752 1643 26754
rect 0 26696 1582 26752
rect 1638 26696 1643 26752
rect 0 26694 1643 26696
rect 16254 26752 16363 26757
rect 16254 26696 16302 26752
rect 16358 26696 16363 26752
rect 16254 26694 16363 26696
rect 0 26664 800 26694
rect 1577 26691 1643 26694
rect 16297 26691 16363 26694
rect 27429 26754 27495 26757
rect 28022 26754 28028 26756
rect 27429 26752 28028 26754
rect 27429 26696 27434 26752
rect 27490 26696 28028 26752
rect 27429 26694 28028 26696
rect 27429 26691 27495 26694
rect 28022 26692 28028 26694
rect 28092 26692 28098 26756
rect 5909 26688 6229 26689
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6229 26688
rect 5909 26623 6229 26624
rect 15840 26688 16160 26689
rect 15840 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15840 26623 16160 26624
rect 25770 26688 26090 26689
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26090 26688
rect 25770 26623 26090 26624
rect 27429 26618 27495 26621
rect 27654 26618 27660 26620
rect 27429 26616 27660 26618
rect 27429 26560 27434 26616
rect 27490 26560 27660 26616
rect 27429 26558 27660 26560
rect 27429 26555 27495 26558
rect 27654 26556 27660 26558
rect 27724 26556 27730 26620
rect 28901 26616 28967 26621
rect 28901 26560 28906 26616
rect 28962 26560 28967 26616
rect 28901 26555 28967 26560
rect 26049 26482 26115 26485
rect 26233 26482 26299 26485
rect 26049 26480 26299 26482
rect 26049 26424 26054 26480
rect 26110 26424 26238 26480
rect 26294 26424 26299 26480
rect 26049 26422 26299 26424
rect 28904 26482 28964 26555
rect 31200 26482 32000 26512
rect 28904 26422 32000 26482
rect 26049 26419 26115 26422
rect 26233 26419 26299 26422
rect 31200 26392 32000 26422
rect 10874 26144 11194 26145
rect 0 26074 800 26104
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 26079 11194 26080
rect 20805 26144 21125 26145
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 20805 26079 21125 26080
rect 1577 26074 1643 26077
rect 0 26072 1643 26074
rect 0 26016 1582 26072
rect 1638 26016 1643 26072
rect 0 26014 1643 26016
rect 0 25984 800 26014
rect 1577 26011 1643 26014
rect 28901 26074 28967 26077
rect 31200 26074 32000 26104
rect 28901 26072 32000 26074
rect 28901 26016 28906 26072
rect 28962 26016 32000 26072
rect 28901 26014 32000 26016
rect 28901 26011 28967 26014
rect 31200 25984 32000 26014
rect 28206 25876 28212 25940
rect 28276 25938 28282 25940
rect 28625 25938 28691 25941
rect 28901 25940 28967 25941
rect 28901 25938 28948 25940
rect 28276 25936 28691 25938
rect 28276 25880 28630 25936
rect 28686 25880 28691 25936
rect 28276 25878 28691 25880
rect 28856 25936 28948 25938
rect 28856 25880 28906 25936
rect 28856 25878 28948 25880
rect 28276 25876 28282 25878
rect 28625 25875 28691 25878
rect 28901 25876 28948 25878
rect 29012 25876 29018 25940
rect 28901 25875 28967 25876
rect 26550 25740 26556 25804
rect 26620 25802 26626 25804
rect 29085 25802 29151 25805
rect 26620 25800 29151 25802
rect 26620 25744 29090 25800
rect 29146 25744 29151 25800
rect 26620 25742 29151 25744
rect 26620 25740 26626 25742
rect 29085 25739 29151 25742
rect 5909 25600 6229 25601
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6229 25600
rect 5909 25535 6229 25536
rect 15840 25600 16160 25601
rect 15840 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15840 25535 16160 25536
rect 25770 25600 26090 25601
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26090 25600
rect 25770 25535 26090 25536
rect 30005 25530 30071 25533
rect 31200 25530 32000 25560
rect 30005 25528 32000 25530
rect 30005 25472 30010 25528
rect 30066 25472 32000 25528
rect 30005 25470 32000 25472
rect 30005 25467 30071 25470
rect 31200 25440 32000 25470
rect 0 25394 800 25424
rect 1577 25394 1643 25397
rect 0 25392 1643 25394
rect 0 25336 1582 25392
rect 1638 25336 1643 25392
rect 0 25334 1643 25336
rect 0 25304 800 25334
rect 1577 25331 1643 25334
rect 24853 25396 24919 25397
rect 24853 25392 24900 25396
rect 24964 25394 24970 25396
rect 24853 25336 24858 25392
rect 24853 25332 24900 25336
rect 24964 25334 25010 25394
rect 24964 25332 24970 25334
rect 24853 25331 24919 25332
rect 25313 25260 25379 25261
rect 25262 25258 25268 25260
rect 25222 25198 25268 25258
rect 25332 25256 25379 25260
rect 25374 25200 25379 25256
rect 25262 25196 25268 25198
rect 25332 25196 25379 25200
rect 25313 25195 25379 25196
rect 26785 25258 26851 25261
rect 26785 25256 26986 25258
rect 26785 25200 26790 25256
rect 26846 25200 26986 25256
rect 26785 25198 26986 25200
rect 26785 25195 26851 25198
rect 10874 25056 11194 25057
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 24991 11194 24992
rect 20805 25056 21125 25057
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 24991 21125 24992
rect 26926 24989 26986 25198
rect 27286 25196 27292 25260
rect 27356 25258 27362 25260
rect 27613 25258 27679 25261
rect 27356 25256 27679 25258
rect 27356 25200 27618 25256
rect 27674 25200 27679 25256
rect 27356 25198 27679 25200
rect 27356 25196 27362 25198
rect 27613 25195 27679 25198
rect 28349 25122 28415 25125
rect 31200 25122 32000 25152
rect 28349 25120 32000 25122
rect 28349 25064 28354 25120
rect 28410 25064 32000 25120
rect 28349 25062 32000 25064
rect 28349 25059 28415 25062
rect 31200 25032 32000 25062
rect 26877 24984 26986 24989
rect 26877 24928 26882 24984
rect 26938 24928 26986 24984
rect 26877 24926 26986 24928
rect 26877 24923 26943 24926
rect 21909 24850 21975 24853
rect 22134 24850 22140 24852
rect 21909 24848 22140 24850
rect 21909 24792 21914 24848
rect 21970 24792 22140 24848
rect 21909 24790 22140 24792
rect 21909 24787 21975 24790
rect 22134 24788 22140 24790
rect 22204 24850 22210 24852
rect 22921 24850 22987 24853
rect 24577 24850 24643 24853
rect 22204 24848 22987 24850
rect 22204 24792 22926 24848
rect 22982 24792 22987 24848
rect 22204 24790 22987 24792
rect 22204 24788 22210 24790
rect 22921 24787 22987 24790
rect 24350 24848 24643 24850
rect 24350 24792 24582 24848
rect 24638 24792 24643 24848
rect 24350 24790 24643 24792
rect 0 24714 800 24744
rect 24350 24717 24410 24790
rect 24577 24787 24643 24790
rect 30097 24850 30163 24853
rect 30230 24850 30236 24852
rect 30097 24848 30236 24850
rect 30097 24792 30102 24848
rect 30158 24792 30236 24848
rect 30097 24790 30236 24792
rect 30097 24787 30163 24790
rect 30230 24788 30236 24790
rect 30300 24788 30306 24852
rect 1577 24714 1643 24717
rect 0 24712 1643 24714
rect 0 24656 1582 24712
rect 1638 24656 1643 24712
rect 0 24654 1643 24656
rect 0 24624 800 24654
rect 1577 24651 1643 24654
rect 24301 24712 24410 24717
rect 26233 24716 26299 24717
rect 24301 24656 24306 24712
rect 24362 24656 24410 24712
rect 24301 24654 24410 24656
rect 24301 24651 24367 24654
rect 26182 24652 26188 24716
rect 26252 24714 26299 24716
rect 26252 24712 26344 24714
rect 26294 24656 26344 24712
rect 26252 24654 26344 24656
rect 26252 24652 26299 24654
rect 26233 24651 26299 24652
rect 28993 24578 29059 24581
rect 31200 24578 32000 24608
rect 28993 24576 32000 24578
rect 28993 24520 28998 24576
rect 29054 24520 32000 24576
rect 28993 24518 32000 24520
rect 28993 24515 29059 24518
rect 5909 24512 6229 24513
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6229 24512
rect 5909 24447 6229 24448
rect 15840 24512 16160 24513
rect 15840 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15840 24447 16160 24448
rect 25770 24512 26090 24513
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26090 24512
rect 31200 24488 32000 24518
rect 25770 24447 26090 24448
rect 24945 24170 25011 24173
rect 25262 24170 25268 24172
rect 24945 24168 25268 24170
rect 24945 24112 24950 24168
rect 25006 24112 25268 24168
rect 24945 24110 25268 24112
rect 24945 24107 25011 24110
rect 25262 24108 25268 24110
rect 25332 24108 25338 24172
rect 28901 24170 28967 24173
rect 31200 24170 32000 24200
rect 28901 24168 32000 24170
rect 28901 24112 28906 24168
rect 28962 24112 32000 24168
rect 28901 24110 32000 24112
rect 28901 24107 28967 24110
rect 31200 24080 32000 24110
rect 0 24034 800 24064
rect 1577 24034 1643 24037
rect 0 24032 1643 24034
rect 0 23976 1582 24032
rect 1638 23976 1643 24032
rect 0 23974 1643 23976
rect 0 23944 800 23974
rect 1577 23971 1643 23974
rect 26734 23972 26740 24036
rect 26804 24034 26810 24036
rect 27797 24034 27863 24037
rect 26804 24032 27863 24034
rect 26804 23976 27802 24032
rect 27858 23976 27863 24032
rect 26804 23974 27863 23976
rect 26804 23972 26810 23974
rect 27797 23971 27863 23974
rect 10874 23968 11194 23969
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 23903 11194 23904
rect 20805 23968 21125 23969
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 20805 23903 21125 23904
rect 27470 23836 27476 23900
rect 27540 23898 27546 23900
rect 28717 23898 28783 23901
rect 27540 23896 28783 23898
rect 27540 23840 28722 23896
rect 28778 23840 28783 23896
rect 27540 23838 28783 23840
rect 27540 23836 27546 23838
rect 28717 23835 28783 23838
rect 27797 23762 27863 23765
rect 28022 23762 28028 23764
rect 27797 23760 28028 23762
rect 27797 23704 27802 23760
rect 27858 23704 28028 23760
rect 27797 23702 28028 23704
rect 27797 23699 27863 23702
rect 28022 23700 28028 23702
rect 28092 23700 28098 23764
rect 28625 23626 28691 23629
rect 31200 23626 32000 23656
rect 28625 23624 32000 23626
rect 28625 23568 28630 23624
rect 28686 23568 32000 23624
rect 28625 23566 32000 23568
rect 28625 23563 28691 23566
rect 31200 23536 32000 23566
rect 0 23490 800 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 800 23430
rect 1577 23427 1643 23430
rect 5909 23424 6229 23425
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6229 23424
rect 5909 23359 6229 23360
rect 15840 23424 16160 23425
rect 15840 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15840 23359 16160 23360
rect 25770 23424 26090 23425
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26090 23424
rect 25770 23359 26090 23360
rect 22369 23218 22435 23221
rect 29177 23218 29243 23221
rect 31200 23218 32000 23248
rect 22369 23216 22570 23218
rect 22369 23160 22374 23216
rect 22430 23160 22570 23216
rect 22369 23158 22570 23160
rect 22369 23155 22435 23158
rect 10874 22880 11194 22881
rect 0 22810 800 22840
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 10874 22815 11194 22816
rect 20805 22880 21125 22881
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 20805 22815 21125 22816
rect 1577 22810 1643 22813
rect 0 22808 1643 22810
rect 0 22752 1582 22808
rect 1638 22752 1643 22808
rect 0 22750 1643 22752
rect 0 22720 800 22750
rect 1577 22747 1643 22750
rect 22510 22674 22570 23158
rect 29177 23216 32000 23218
rect 29177 23160 29182 23216
rect 29238 23160 32000 23216
rect 29177 23158 32000 23160
rect 29177 23155 29243 23158
rect 31200 23128 32000 23158
rect 24894 23020 24900 23084
rect 24964 23082 24970 23084
rect 25405 23082 25471 23085
rect 24964 23080 25471 23082
rect 24964 23024 25410 23080
rect 25466 23024 25471 23080
rect 24964 23022 25471 23024
rect 24964 23020 24970 23022
rect 25405 23019 25471 23022
rect 24710 22748 24716 22812
rect 24780 22810 24786 22812
rect 26182 22810 26188 22812
rect 24780 22750 26188 22810
rect 24780 22748 24786 22750
rect 26182 22748 26188 22750
rect 26252 22810 26258 22812
rect 26693 22810 26759 22813
rect 26252 22808 26759 22810
rect 26252 22752 26698 22808
rect 26754 22752 26759 22808
rect 26252 22750 26759 22752
rect 26252 22748 26258 22750
rect 26693 22747 26759 22750
rect 29913 22810 29979 22813
rect 31200 22810 32000 22840
rect 29913 22808 32000 22810
rect 29913 22752 29918 22808
rect 29974 22752 32000 22808
rect 29913 22750 32000 22752
rect 29913 22747 29979 22750
rect 31200 22720 32000 22750
rect 22645 22674 22711 22677
rect 22510 22672 22711 22674
rect 22510 22616 22650 22672
rect 22706 22616 22711 22672
rect 22510 22614 22711 22616
rect 22645 22611 22711 22614
rect 25589 22538 25655 22541
rect 30281 22538 30347 22541
rect 30414 22538 30420 22540
rect 25589 22536 26296 22538
rect 25589 22480 25594 22536
rect 25650 22480 26296 22536
rect 25589 22478 26296 22480
rect 25589 22475 25655 22478
rect 25037 22402 25103 22405
rect 25630 22402 25636 22404
rect 25037 22400 25636 22402
rect 25037 22344 25042 22400
rect 25098 22344 25636 22400
rect 25037 22342 25636 22344
rect 25037 22339 25103 22342
rect 25630 22340 25636 22342
rect 25700 22340 25706 22404
rect 5909 22336 6229 22337
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6229 22336
rect 5909 22271 6229 22272
rect 15840 22336 16160 22337
rect 15840 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15840 22271 16160 22272
rect 25770 22336 26090 22337
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26090 22336
rect 25770 22271 26090 22272
rect 0 22130 800 22160
rect 26236 22133 26296 22478
rect 30281 22536 30420 22538
rect 30281 22480 30286 22536
rect 30342 22480 30420 22536
rect 30281 22478 30420 22480
rect 30281 22475 30347 22478
rect 30414 22476 30420 22478
rect 30484 22476 30490 22540
rect 28901 22402 28967 22405
rect 28901 22400 30666 22402
rect 28901 22344 28906 22400
rect 28962 22344 30666 22400
rect 28901 22342 30666 22344
rect 28901 22339 28967 22342
rect 27429 22266 27495 22269
rect 30606 22266 30666 22342
rect 31200 22266 32000 22296
rect 27429 22264 28504 22266
rect 27429 22208 27434 22264
rect 27490 22208 28504 22264
rect 27429 22206 28504 22208
rect 30606 22206 32000 22266
rect 27429 22203 27495 22206
rect 28444 22133 28504 22206
rect 31200 22176 32000 22206
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 800 22070
rect 1577 22067 1643 22070
rect 24945 22130 25011 22133
rect 25446 22130 25452 22132
rect 24945 22128 25452 22130
rect 24945 22072 24950 22128
rect 25006 22072 25452 22128
rect 24945 22070 25452 22072
rect 24945 22067 25011 22070
rect 25446 22068 25452 22070
rect 25516 22068 25522 22132
rect 26233 22128 26299 22133
rect 26785 22132 26851 22133
rect 26233 22072 26238 22128
rect 26294 22072 26299 22128
rect 26233 22067 26299 22072
rect 26734 22068 26740 22132
rect 26804 22130 26851 22132
rect 26804 22128 26896 22130
rect 26846 22072 26896 22128
rect 26804 22070 26896 22072
rect 26804 22068 26851 22070
rect 27102 22068 27108 22132
rect 27172 22130 27178 22132
rect 27521 22130 27587 22133
rect 27172 22128 27587 22130
rect 27172 22072 27526 22128
rect 27582 22072 27587 22128
rect 27172 22070 27587 22072
rect 27172 22068 27178 22070
rect 26785 22067 26851 22068
rect 27521 22067 27587 22070
rect 28441 22128 28507 22133
rect 28441 22072 28446 22128
rect 28502 22072 28507 22128
rect 28441 22067 28507 22072
rect 29637 22130 29703 22133
rect 30097 22130 30163 22133
rect 30230 22130 30236 22132
rect 29637 22128 29930 22130
rect 29637 22072 29642 22128
rect 29698 22072 29930 22128
rect 29637 22070 29930 22072
rect 29637 22067 29703 22070
rect 25037 21994 25103 21997
rect 26877 21994 26943 21997
rect 27797 21996 27863 21997
rect 27797 21994 27844 21996
rect 25037 21992 25330 21994
rect 25037 21936 25042 21992
rect 25098 21936 25330 21992
rect 25037 21934 25330 21936
rect 25037 21931 25103 21934
rect 25270 21861 25330 21934
rect 26877 21992 27170 21994
rect 26877 21936 26882 21992
rect 26938 21936 27170 21992
rect 26877 21934 27170 21936
rect 27752 21992 27844 21994
rect 27752 21936 27802 21992
rect 27752 21934 27844 21936
rect 26877 21931 26943 21934
rect 25270 21856 25379 21861
rect 25270 21800 25318 21856
rect 25374 21800 25379 21856
rect 25270 21798 25379 21800
rect 27110 21858 27170 21934
rect 27797 21932 27844 21934
rect 27908 21932 27914 21996
rect 29126 21932 29132 21996
rect 29196 21994 29202 21996
rect 29870 21994 29930 22070
rect 30097 22128 30236 22130
rect 30097 22072 30102 22128
rect 30158 22072 30236 22128
rect 30097 22070 30236 22072
rect 30097 22067 30163 22070
rect 30230 22068 30236 22070
rect 30300 22068 30306 22132
rect 29196 21934 29930 21994
rect 29196 21932 29202 21934
rect 27797 21931 27863 21932
rect 27245 21858 27311 21861
rect 27110 21856 27311 21858
rect 27110 21800 27250 21856
rect 27306 21800 27311 21856
rect 27110 21798 27311 21800
rect 25313 21795 25379 21798
rect 27245 21795 27311 21798
rect 28073 21858 28139 21861
rect 28441 21858 28507 21861
rect 28073 21856 28507 21858
rect 28073 21800 28078 21856
rect 28134 21800 28446 21856
rect 28502 21800 28507 21856
rect 28073 21798 28507 21800
rect 28073 21795 28139 21798
rect 28441 21795 28507 21798
rect 28901 21858 28967 21861
rect 31200 21858 32000 21888
rect 28901 21856 32000 21858
rect 28901 21800 28906 21856
rect 28962 21800 32000 21856
rect 28901 21798 32000 21800
rect 28901 21795 28967 21798
rect 10874 21792 11194 21793
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 10874 21727 11194 21728
rect 20805 21792 21125 21793
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 31200 21768 32000 21798
rect 20805 21727 21125 21728
rect 24945 21724 25011 21725
rect 24894 21722 24900 21724
rect 24854 21662 24900 21722
rect 24964 21720 25011 21724
rect 25006 21664 25011 21720
rect 24894 21660 24900 21662
rect 24964 21660 25011 21664
rect 24945 21659 25011 21660
rect 0 21450 800 21480
rect 1577 21450 1643 21453
rect 25129 21452 25195 21453
rect 25078 21450 25084 21452
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 25038 21390 25084 21450
rect 25148 21448 25195 21452
rect 25190 21392 25195 21448
rect 0 21360 800 21390
rect 1577 21387 1643 21390
rect 25078 21388 25084 21390
rect 25148 21388 25195 21392
rect 25129 21387 25195 21388
rect 27613 21314 27679 21317
rect 31200 21314 32000 21344
rect 27613 21312 32000 21314
rect 27613 21256 27618 21312
rect 27674 21256 32000 21312
rect 27613 21254 32000 21256
rect 27613 21251 27679 21254
rect 5909 21248 6229 21249
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6229 21248
rect 5909 21183 6229 21184
rect 15840 21248 16160 21249
rect 15840 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15840 21183 16160 21184
rect 25770 21248 26090 21249
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26090 21248
rect 31200 21224 32000 21254
rect 25770 21183 26090 21184
rect 25630 20980 25636 21044
rect 25700 21042 25706 21044
rect 25773 21042 25839 21045
rect 25700 21040 25839 21042
rect 25700 20984 25778 21040
rect 25834 20984 25839 21040
rect 25700 20982 25839 20984
rect 25700 20980 25706 20982
rect 25773 20979 25839 20982
rect 28257 20906 28323 20909
rect 31200 20906 32000 20936
rect 28257 20904 32000 20906
rect 28257 20848 28262 20904
rect 28318 20848 32000 20904
rect 28257 20846 32000 20848
rect 28257 20843 28323 20846
rect 31200 20816 32000 20846
rect 0 20770 800 20800
rect 1577 20770 1643 20773
rect 26417 20772 26483 20773
rect 26366 20770 26372 20772
rect 0 20768 1643 20770
rect 0 20712 1582 20768
rect 1638 20712 1643 20768
rect 0 20710 1643 20712
rect 26326 20710 26372 20770
rect 26436 20768 26483 20772
rect 26478 20712 26483 20768
rect 0 20680 800 20710
rect 1577 20707 1643 20710
rect 26366 20708 26372 20710
rect 26436 20708 26483 20712
rect 26417 20707 26483 20708
rect 10874 20704 11194 20705
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 20639 11194 20640
rect 20805 20704 21125 20705
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 20805 20639 21125 20640
rect 28901 20362 28967 20365
rect 31200 20362 32000 20392
rect 28901 20360 32000 20362
rect 28901 20304 28906 20360
rect 28962 20304 32000 20360
rect 28901 20302 32000 20304
rect 28901 20299 28967 20302
rect 31200 20272 32000 20302
rect 5909 20160 6229 20161
rect 0 20090 800 20120
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6229 20160
rect 5909 20095 6229 20096
rect 15840 20160 16160 20161
rect 15840 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 15840 20095 16160 20096
rect 25770 20160 26090 20161
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26090 20160
rect 25770 20095 26090 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 29269 19954 29335 19957
rect 31200 19954 32000 19984
rect 29269 19952 32000 19954
rect 29269 19896 29274 19952
rect 29330 19896 32000 19952
rect 29269 19894 32000 19896
rect 29269 19891 29335 19894
rect 31200 19864 32000 19894
rect 26509 19818 26575 19821
rect 27061 19818 27127 19821
rect 26509 19816 27127 19818
rect 26509 19760 26514 19816
rect 26570 19760 27066 19816
rect 27122 19760 27127 19816
rect 26509 19758 27127 19760
rect 26509 19755 26575 19758
rect 27061 19755 27127 19758
rect 28717 19818 28783 19821
rect 30414 19818 30420 19820
rect 28717 19816 30420 19818
rect 28717 19760 28722 19816
rect 28778 19760 30420 19816
rect 28717 19758 30420 19760
rect 28717 19755 28783 19758
rect 30414 19756 30420 19758
rect 30484 19756 30490 19820
rect 25262 19620 25268 19684
rect 25332 19682 25338 19684
rect 26509 19682 26575 19685
rect 25332 19680 26575 19682
rect 25332 19624 26514 19680
rect 26570 19624 26575 19680
rect 25332 19622 26575 19624
rect 25332 19620 25338 19622
rect 26509 19619 26575 19622
rect 10874 19616 11194 19617
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 19551 11194 19552
rect 20805 19616 21125 19617
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 19551 21125 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 28809 19410 28875 19413
rect 31200 19410 32000 19440
rect 28809 19408 32000 19410
rect 28809 19352 28814 19408
rect 28870 19352 32000 19408
rect 28809 19350 32000 19352
rect 28809 19347 28875 19350
rect 31200 19320 32000 19350
rect 5909 19072 6229 19073
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6229 19072
rect 5909 19007 6229 19008
rect 15840 19072 16160 19073
rect 15840 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15840 19007 16160 19008
rect 25770 19072 26090 19073
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26090 19072
rect 25770 19007 26090 19008
rect 30005 19002 30071 19005
rect 31200 19002 32000 19032
rect 30005 19000 32000 19002
rect 30005 18944 30010 19000
rect 30066 18944 32000 19000
rect 30005 18942 32000 18944
rect 30005 18939 30071 18942
rect 31200 18912 32000 18942
rect 0 18866 800 18896
rect 1577 18866 1643 18869
rect 0 18864 1643 18866
rect 0 18808 1582 18864
rect 1638 18808 1643 18864
rect 0 18806 1643 18808
rect 0 18776 800 18806
rect 1577 18803 1643 18806
rect 25957 18730 26023 18733
rect 26182 18730 26188 18732
rect 25957 18728 26188 18730
rect 25957 18672 25962 18728
rect 26018 18672 26188 18728
rect 25957 18670 26188 18672
rect 25957 18667 26023 18670
rect 26182 18668 26188 18670
rect 26252 18668 26258 18732
rect 27521 18730 27587 18733
rect 28574 18730 28580 18732
rect 27521 18728 28580 18730
rect 27521 18672 27526 18728
rect 27582 18672 28580 18728
rect 27521 18670 28580 18672
rect 27521 18667 27587 18670
rect 28574 18668 28580 18670
rect 28644 18668 28650 18732
rect 10874 18528 11194 18529
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 18463 11194 18464
rect 20805 18528 21125 18529
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 18463 21125 18464
rect 25313 18458 25379 18461
rect 24902 18456 25379 18458
rect 24902 18400 25318 18456
rect 25374 18400 25379 18456
rect 24902 18398 25379 18400
rect 0 18186 800 18216
rect 24902 18189 24962 18398
rect 25313 18395 25379 18398
rect 29821 18458 29887 18461
rect 31200 18458 32000 18488
rect 29821 18456 32000 18458
rect 29821 18400 29826 18456
rect 29882 18400 32000 18456
rect 29821 18398 32000 18400
rect 29821 18395 29887 18398
rect 31200 18368 32000 18398
rect 27337 18322 27403 18325
rect 26742 18320 27403 18322
rect 26742 18264 27342 18320
rect 27398 18264 27403 18320
rect 26742 18262 27403 18264
rect 1577 18186 1643 18189
rect 0 18184 1643 18186
rect 0 18128 1582 18184
rect 1638 18128 1643 18184
rect 0 18126 1643 18128
rect 0 18096 800 18126
rect 1577 18123 1643 18126
rect 24853 18184 24962 18189
rect 24853 18128 24858 18184
rect 24914 18128 24962 18184
rect 24853 18126 24962 18128
rect 24853 18123 24919 18126
rect 25630 18124 25636 18188
rect 25700 18186 25706 18188
rect 25773 18186 25839 18189
rect 25700 18184 25839 18186
rect 25700 18128 25778 18184
rect 25834 18128 25839 18184
rect 25700 18126 25839 18128
rect 25700 18124 25706 18126
rect 25773 18123 25839 18126
rect 5909 17984 6229 17985
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6229 17984
rect 5909 17919 6229 17920
rect 15840 17984 16160 17985
rect 15840 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15840 17919 16160 17920
rect 25770 17984 26090 17985
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26090 17984
rect 25770 17919 26090 17920
rect 26049 17642 26115 17645
rect 26182 17642 26188 17644
rect 26049 17640 26188 17642
rect 26049 17584 26054 17640
rect 26110 17584 26188 17640
rect 26049 17582 26188 17584
rect 26049 17579 26115 17582
rect 26182 17580 26188 17582
rect 26252 17580 26258 17644
rect 26601 17642 26667 17645
rect 26742 17642 26802 18262
rect 27337 18259 27403 18262
rect 28993 18186 29059 18189
rect 29126 18186 29132 18188
rect 28993 18184 29132 18186
rect 28993 18128 28998 18184
rect 29054 18128 29132 18184
rect 28993 18126 29132 18128
rect 28993 18123 29059 18126
rect 29126 18124 29132 18126
rect 29196 18124 29202 18188
rect 29913 18050 29979 18053
rect 31200 18050 32000 18080
rect 29913 18048 32000 18050
rect 29913 17992 29918 18048
rect 29974 17992 32000 18048
rect 29913 17990 32000 17992
rect 29913 17987 29979 17990
rect 31200 17960 32000 17990
rect 26601 17640 26802 17642
rect 26601 17584 26606 17640
rect 26662 17584 26802 17640
rect 26601 17582 26802 17584
rect 26601 17579 26667 17582
rect 0 17506 800 17536
rect 1577 17506 1643 17509
rect 0 17504 1643 17506
rect 0 17448 1582 17504
rect 1638 17448 1643 17504
rect 0 17446 1643 17448
rect 0 17416 800 17446
rect 1577 17443 1643 17446
rect 28349 17506 28415 17509
rect 31200 17506 32000 17536
rect 28349 17504 32000 17506
rect 28349 17448 28354 17504
rect 28410 17448 32000 17504
rect 28349 17446 32000 17448
rect 28349 17443 28415 17446
rect 10874 17440 11194 17441
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10874 17375 11194 17376
rect 20805 17440 21125 17441
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 31200 17416 32000 17446
rect 20805 17375 21125 17376
rect 28809 17098 28875 17101
rect 31200 17098 32000 17128
rect 28809 17096 32000 17098
rect 28809 17040 28814 17096
rect 28870 17040 32000 17096
rect 28809 17038 32000 17040
rect 28809 17035 28875 17038
rect 31200 17008 32000 17038
rect 5909 16896 6229 16897
rect 0 16826 800 16856
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6229 16896
rect 5909 16831 6229 16832
rect 15840 16896 16160 16897
rect 15840 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15840 16831 16160 16832
rect 25770 16896 26090 16897
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26090 16896
rect 25770 16831 26090 16832
rect 1577 16826 1643 16829
rect 0 16824 1643 16826
rect 0 16768 1582 16824
rect 1638 16768 1643 16824
rect 0 16766 1643 16768
rect 0 16736 800 16766
rect 1577 16763 1643 16766
rect 16849 16826 16915 16829
rect 19241 16826 19307 16829
rect 16849 16824 19307 16826
rect 16849 16768 16854 16824
rect 16910 16768 19246 16824
rect 19302 16768 19307 16824
rect 16849 16766 19307 16768
rect 16849 16763 16915 16766
rect 19241 16763 19307 16766
rect 18873 16690 18939 16693
rect 19885 16690 19951 16693
rect 18873 16688 19951 16690
rect 18873 16632 18878 16688
rect 18934 16632 19890 16688
rect 19946 16632 19951 16688
rect 18873 16630 19951 16632
rect 18873 16627 18939 16630
rect 19885 16627 19951 16630
rect 28901 16690 28967 16693
rect 31200 16690 32000 16720
rect 28901 16688 32000 16690
rect 28901 16632 28906 16688
rect 28962 16632 32000 16688
rect 28901 16630 32000 16632
rect 28901 16627 28967 16630
rect 31200 16600 32000 16630
rect 18873 16554 18939 16557
rect 19517 16554 19583 16557
rect 18873 16552 19583 16554
rect 18873 16496 18878 16552
rect 18934 16496 19522 16552
rect 19578 16496 19583 16552
rect 18873 16494 19583 16496
rect 18873 16491 18939 16494
rect 19517 16491 19583 16494
rect 18689 16418 18755 16421
rect 19885 16418 19951 16421
rect 18689 16416 19951 16418
rect 18689 16360 18694 16416
rect 18750 16360 19890 16416
rect 19946 16360 19951 16416
rect 18689 16358 19951 16360
rect 18689 16355 18755 16358
rect 19885 16355 19951 16358
rect 10874 16352 11194 16353
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 16287 11194 16288
rect 20805 16352 21125 16353
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 20805 16287 21125 16288
rect 27613 16282 27679 16285
rect 27889 16282 27955 16285
rect 27613 16280 27955 16282
rect 27613 16224 27618 16280
rect 27674 16224 27894 16280
rect 27950 16224 27955 16280
rect 27613 16222 27955 16224
rect 27613 16219 27679 16222
rect 27889 16219 27955 16222
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 17718 16084 17724 16148
rect 17788 16146 17794 16148
rect 25037 16146 25103 16149
rect 17788 16144 25103 16146
rect 17788 16088 25042 16144
rect 25098 16088 25103 16144
rect 17788 16086 25103 16088
rect 17788 16084 17794 16086
rect 25037 16083 25103 16086
rect 30097 16146 30163 16149
rect 31200 16146 32000 16176
rect 30097 16144 32000 16146
rect 30097 16088 30102 16144
rect 30158 16088 32000 16144
rect 30097 16086 32000 16088
rect 30097 16083 30163 16086
rect 31200 16056 32000 16086
rect 18137 15874 18203 15877
rect 21173 15874 21239 15877
rect 18137 15872 21239 15874
rect 18137 15816 18142 15872
rect 18198 15816 21178 15872
rect 21234 15816 21239 15872
rect 18137 15814 21239 15816
rect 18137 15811 18203 15814
rect 21173 15811 21239 15814
rect 5909 15808 6229 15809
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6229 15808
rect 5909 15743 6229 15744
rect 15840 15808 16160 15809
rect 15840 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15840 15743 16160 15744
rect 25770 15808 26090 15809
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26090 15808
rect 25770 15743 26090 15744
rect 29913 15738 29979 15741
rect 31200 15738 32000 15768
rect 29913 15736 32000 15738
rect 29913 15680 29918 15736
rect 29974 15680 32000 15736
rect 29913 15678 32000 15680
rect 29913 15675 29979 15678
rect 31200 15648 32000 15678
rect 0 15466 800 15496
rect 1577 15466 1643 15469
rect 0 15464 1643 15466
rect 0 15408 1582 15464
rect 1638 15408 1643 15464
rect 0 15406 1643 15408
rect 0 15376 800 15406
rect 1577 15403 1643 15406
rect 27613 15466 27679 15469
rect 29494 15466 29500 15468
rect 27613 15464 29500 15466
rect 27613 15408 27618 15464
rect 27674 15408 29500 15464
rect 27613 15406 29500 15408
rect 27613 15403 27679 15406
rect 29494 15404 29500 15406
rect 29564 15404 29570 15468
rect 25589 15332 25655 15333
rect 25589 15328 25636 15332
rect 25700 15330 25706 15332
rect 25589 15272 25594 15328
rect 25589 15268 25636 15272
rect 25700 15270 25746 15330
rect 25700 15268 25706 15270
rect 25589 15267 25655 15268
rect 10874 15264 11194 15265
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 15199 11194 15200
rect 20805 15264 21125 15265
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 15199 21125 15200
rect 28257 15194 28323 15197
rect 28390 15194 28396 15196
rect 28257 15192 28396 15194
rect 28257 15136 28262 15192
rect 28318 15136 28396 15192
rect 28257 15134 28396 15136
rect 28257 15131 28323 15134
rect 28390 15132 28396 15134
rect 28460 15132 28466 15196
rect 29913 15194 29979 15197
rect 31200 15194 32000 15224
rect 29913 15192 32000 15194
rect 29913 15136 29918 15192
rect 29974 15136 32000 15192
rect 29913 15134 32000 15136
rect 29913 15131 29979 15134
rect 31200 15104 32000 15134
rect 0 14786 800 14816
rect 1577 14786 1643 14789
rect 0 14784 1643 14786
rect 0 14728 1582 14784
rect 1638 14728 1643 14784
rect 0 14726 1643 14728
rect 0 14696 800 14726
rect 1577 14723 1643 14726
rect 29821 14786 29887 14789
rect 31200 14786 32000 14816
rect 29821 14784 32000 14786
rect 29821 14728 29826 14784
rect 29882 14728 32000 14784
rect 29821 14726 32000 14728
rect 29821 14723 29887 14726
rect 5909 14720 6229 14721
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6229 14720
rect 5909 14655 6229 14656
rect 15840 14720 16160 14721
rect 15840 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15840 14655 16160 14656
rect 25770 14720 26090 14721
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26090 14720
rect 31200 14696 32000 14726
rect 25770 14655 26090 14656
rect 19517 14514 19583 14517
rect 27981 14514 28047 14517
rect 19517 14512 28047 14514
rect 19517 14456 19522 14512
rect 19578 14456 27986 14512
rect 28042 14456 28047 14512
rect 19517 14454 28047 14456
rect 19517 14451 19583 14454
rect 27981 14451 28047 14454
rect 0 14242 800 14272
rect 1577 14242 1643 14245
rect 0 14240 1643 14242
rect 0 14184 1582 14240
rect 1638 14184 1643 14240
rect 0 14182 1643 14184
rect 0 14152 800 14182
rect 1577 14179 1643 14182
rect 28901 14242 28967 14245
rect 31200 14242 32000 14272
rect 28901 14240 32000 14242
rect 28901 14184 28906 14240
rect 28962 14184 32000 14240
rect 28901 14182 32000 14184
rect 28901 14179 28967 14182
rect 10874 14176 11194 14177
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 14111 11194 14112
rect 20805 14176 21125 14177
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 31200 14152 32000 14182
rect 20805 14111 21125 14112
rect 25773 14106 25839 14109
rect 26785 14106 26851 14109
rect 25773 14104 26851 14106
rect 25773 14048 25778 14104
rect 25834 14048 26790 14104
rect 26846 14048 26851 14104
rect 25773 14046 26851 14048
rect 25773 14043 25839 14046
rect 26785 14043 26851 14046
rect 28533 14106 28599 14109
rect 29310 14106 29316 14108
rect 28533 14104 29316 14106
rect 28533 14048 28538 14104
rect 28594 14048 29316 14104
rect 28533 14046 29316 14048
rect 28533 14043 28599 14046
rect 29310 14044 29316 14046
rect 29380 14044 29386 14108
rect 27613 13834 27679 13837
rect 31200 13834 32000 13864
rect 27613 13832 32000 13834
rect 27613 13776 27618 13832
rect 27674 13776 32000 13832
rect 27613 13774 32000 13776
rect 27613 13771 27679 13774
rect 31200 13744 32000 13774
rect 5909 13632 6229 13633
rect 0 13562 800 13592
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6229 13632
rect 5909 13567 6229 13568
rect 15840 13632 16160 13633
rect 15840 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15840 13567 16160 13568
rect 25770 13632 26090 13633
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26090 13632
rect 25770 13567 26090 13568
rect 1577 13562 1643 13565
rect 0 13560 1643 13562
rect 0 13504 1582 13560
rect 1638 13504 1643 13560
rect 0 13502 1643 13504
rect 0 13472 800 13502
rect 1577 13499 1643 13502
rect 28993 13290 29059 13293
rect 31200 13290 32000 13320
rect 28993 13288 32000 13290
rect 28993 13232 28998 13288
rect 29054 13232 32000 13288
rect 28993 13230 32000 13232
rect 28993 13227 29059 13230
rect 31200 13200 32000 13230
rect 10874 13088 11194 13089
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10874 13023 11194 13024
rect 20805 13088 21125 13089
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 20805 13023 21125 13024
rect 0 12882 800 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 800 12822
rect 1577 12819 1643 12822
rect 28809 12882 28875 12885
rect 31200 12882 32000 12912
rect 28809 12880 32000 12882
rect 28809 12824 28814 12880
rect 28870 12824 32000 12880
rect 28809 12822 32000 12824
rect 28809 12819 28875 12822
rect 31200 12792 32000 12822
rect 5909 12544 6229 12545
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6229 12544
rect 5909 12479 6229 12480
rect 15840 12544 16160 12545
rect 15840 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15840 12479 16160 12480
rect 25770 12544 26090 12545
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26090 12544
rect 25770 12479 26090 12480
rect 28901 12338 28967 12341
rect 31200 12338 32000 12368
rect 28901 12336 32000 12338
rect 28901 12280 28906 12336
rect 28962 12280 32000 12336
rect 28901 12278 32000 12280
rect 28901 12275 28967 12278
rect 31200 12248 32000 12278
rect 0 12202 800 12232
rect 1577 12202 1643 12205
rect 0 12200 1643 12202
rect 0 12144 1582 12200
rect 1638 12144 1643 12200
rect 0 12142 1643 12144
rect 0 12112 800 12142
rect 1577 12139 1643 12142
rect 26141 12068 26207 12069
rect 26141 12064 26188 12068
rect 26252 12066 26258 12068
rect 26141 12008 26146 12064
rect 26141 12004 26188 12008
rect 26252 12006 26298 12066
rect 26252 12004 26258 12006
rect 26141 12003 26207 12004
rect 10874 12000 11194 12001
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 10874 11935 11194 11936
rect 20805 12000 21125 12001
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 20805 11935 21125 11936
rect 28165 11930 28231 11933
rect 31200 11930 32000 11960
rect 28165 11928 32000 11930
rect 28165 11872 28170 11928
rect 28226 11872 32000 11928
rect 28165 11870 32000 11872
rect 28165 11867 28231 11870
rect 31200 11840 32000 11870
rect 0 11522 800 11552
rect 1577 11522 1643 11525
rect 0 11520 1643 11522
rect 0 11464 1582 11520
rect 1638 11464 1643 11520
rect 0 11462 1643 11464
rect 0 11432 800 11462
rect 1577 11459 1643 11462
rect 29361 11522 29427 11525
rect 31200 11522 32000 11552
rect 29361 11520 32000 11522
rect 29361 11464 29366 11520
rect 29422 11464 32000 11520
rect 29361 11462 32000 11464
rect 29361 11459 29427 11462
rect 5909 11456 6229 11457
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6229 11456
rect 5909 11391 6229 11392
rect 15840 11456 16160 11457
rect 15840 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15840 11391 16160 11392
rect 25770 11456 26090 11457
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26090 11456
rect 31200 11432 32000 11462
rect 25770 11391 26090 11392
rect 19609 11250 19675 11253
rect 21357 11250 21423 11253
rect 19609 11248 21423 11250
rect 19609 11192 19614 11248
rect 19670 11192 21362 11248
rect 21418 11192 21423 11248
rect 19609 11190 21423 11192
rect 19609 11187 19675 11190
rect 21357 11187 21423 11190
rect 29269 10978 29335 10981
rect 31200 10978 32000 11008
rect 29269 10976 32000 10978
rect 29269 10920 29274 10976
rect 29330 10920 32000 10976
rect 29269 10918 32000 10920
rect 29269 10915 29335 10918
rect 10874 10912 11194 10913
rect 0 10842 800 10872
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 10847 11194 10848
rect 20805 10912 21125 10913
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 31200 10888 32000 10918
rect 20805 10847 21125 10848
rect 1577 10842 1643 10845
rect 0 10840 1643 10842
rect 0 10784 1582 10840
rect 1638 10784 1643 10840
rect 0 10782 1643 10784
rect 0 10752 800 10782
rect 1577 10779 1643 10782
rect 26509 10842 26575 10845
rect 26785 10842 26851 10845
rect 26509 10840 26851 10842
rect 26509 10784 26514 10840
rect 26570 10784 26790 10840
rect 26846 10784 26851 10840
rect 26509 10782 26851 10784
rect 26509 10779 26575 10782
rect 26785 10779 26851 10782
rect 29913 10570 29979 10573
rect 31200 10570 32000 10600
rect 29913 10568 32000 10570
rect 29913 10512 29918 10568
rect 29974 10512 32000 10568
rect 29913 10510 32000 10512
rect 29913 10507 29979 10510
rect 31200 10480 32000 10510
rect 5909 10368 6229 10369
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6229 10368
rect 5909 10303 6229 10304
rect 15840 10368 16160 10369
rect 15840 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15840 10303 16160 10304
rect 25770 10368 26090 10369
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26090 10368
rect 25770 10303 26090 10304
rect 0 10162 800 10192
rect 1577 10162 1643 10165
rect 0 10160 1643 10162
rect 0 10104 1582 10160
rect 1638 10104 1643 10160
rect 0 10102 1643 10104
rect 0 10072 800 10102
rect 1577 10099 1643 10102
rect 29729 10026 29795 10029
rect 31200 10026 32000 10056
rect 29729 10024 32000 10026
rect 29729 9968 29734 10024
rect 29790 9968 32000 10024
rect 29729 9966 32000 9968
rect 29729 9963 29795 9966
rect 31200 9936 32000 9966
rect 10874 9824 11194 9825
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 9759 11194 9760
rect 20805 9824 21125 9825
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 20805 9759 21125 9760
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 28717 9618 28783 9621
rect 31200 9618 32000 9648
rect 28717 9616 32000 9618
rect 28717 9560 28722 9616
rect 28778 9560 32000 9616
rect 28717 9558 32000 9560
rect 28717 9555 28783 9558
rect 31200 9528 32000 9558
rect 5909 9280 6229 9281
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6229 9280
rect 5909 9215 6229 9216
rect 15840 9280 16160 9281
rect 15840 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15840 9215 16160 9216
rect 25770 9280 26090 9281
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26090 9280
rect 25770 9215 26090 9216
rect 28901 9074 28967 9077
rect 31200 9074 32000 9104
rect 28901 9072 32000 9074
rect 28901 9016 28906 9072
rect 28962 9016 32000 9072
rect 28901 9014 32000 9016
rect 28901 9011 28967 9014
rect 31200 8984 32000 9014
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 10874 8736 11194 8737
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 8671 11194 8672
rect 20805 8736 21125 8737
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 8671 21125 8672
rect 28901 8666 28967 8669
rect 31200 8666 32000 8696
rect 28901 8664 32000 8666
rect 28901 8608 28906 8664
rect 28962 8608 32000 8664
rect 28901 8606 32000 8608
rect 28901 8603 28967 8606
rect 31200 8576 32000 8606
rect 0 8258 800 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 800 8198
rect 1577 8195 1643 8198
rect 5909 8192 6229 8193
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6229 8192
rect 5909 8127 6229 8128
rect 15840 8192 16160 8193
rect 15840 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15840 8127 16160 8128
rect 25770 8192 26090 8193
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26090 8192
rect 25770 8127 26090 8128
rect 29821 8122 29887 8125
rect 31200 8122 32000 8152
rect 29821 8120 32000 8122
rect 29821 8064 29826 8120
rect 29882 8064 32000 8120
rect 29821 8062 32000 8064
rect 29821 8059 29887 8062
rect 31200 8032 32000 8062
rect 27705 7714 27771 7717
rect 31200 7714 32000 7744
rect 27705 7712 32000 7714
rect 27705 7656 27710 7712
rect 27766 7656 32000 7712
rect 27705 7654 32000 7656
rect 27705 7651 27771 7654
rect 10874 7648 11194 7649
rect 0 7578 800 7608
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 7583 11194 7584
rect 20805 7648 21125 7649
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 31200 7624 32000 7654
rect 20805 7583 21125 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 27613 7170 27679 7173
rect 31200 7170 32000 7200
rect 27613 7168 32000 7170
rect 27613 7112 27618 7168
rect 27674 7112 32000 7168
rect 27613 7110 32000 7112
rect 27613 7107 27679 7110
rect 5909 7104 6229 7105
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6229 7104
rect 5909 7039 6229 7040
rect 15840 7104 16160 7105
rect 15840 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15840 7039 16160 7040
rect 25770 7104 26090 7105
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26090 7104
rect 31200 7080 32000 7110
rect 25770 7039 26090 7040
rect 0 6898 800 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 800 6838
rect 1577 6835 1643 6838
rect 28809 6762 28875 6765
rect 31200 6762 32000 6792
rect 28809 6760 32000 6762
rect 28809 6704 28814 6760
rect 28870 6704 32000 6760
rect 28809 6702 32000 6704
rect 28809 6699 28875 6702
rect 31200 6672 32000 6702
rect 10874 6560 11194 6561
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 6495 11194 6496
rect 20805 6560 21125 6561
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 6495 21125 6496
rect 29821 6490 29887 6493
rect 30046 6490 30052 6492
rect 29821 6488 30052 6490
rect 29821 6432 29826 6488
rect 29882 6432 30052 6488
rect 29821 6430 30052 6432
rect 29821 6427 29887 6430
rect 30046 6428 30052 6430
rect 30116 6428 30122 6492
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 30097 6218 30163 6221
rect 31200 6218 32000 6248
rect 30097 6216 32000 6218
rect 30097 6160 30102 6216
rect 30158 6160 32000 6216
rect 30097 6158 32000 6160
rect 30097 6155 30163 6158
rect 31200 6128 32000 6158
rect 5909 6016 6229 6017
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6229 6016
rect 5909 5951 6229 5952
rect 15840 6016 16160 6017
rect 15840 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15840 5951 16160 5952
rect 25770 6016 26090 6017
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26090 6016
rect 25770 5951 26090 5952
rect 31200 5720 32000 5840
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 10874 5472 11194 5473
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 5407 11194 5408
rect 20805 5472 21125 5473
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 20805 5407 21125 5408
rect 29678 5340 29684 5404
rect 29748 5402 29754 5404
rect 29821 5402 29887 5405
rect 29748 5400 29887 5402
rect 29748 5344 29826 5400
rect 29882 5344 29887 5400
rect 29748 5342 29887 5344
rect 29748 5340 29754 5342
rect 29821 5339 29887 5342
rect 31200 5312 32000 5432
rect 0 4994 800 5024
rect 1577 4994 1643 4997
rect 0 4992 1643 4994
rect 0 4936 1582 4992
rect 1638 4936 1643 4992
rect 0 4934 1643 4936
rect 0 4904 800 4934
rect 1577 4931 1643 4934
rect 5909 4928 6229 4929
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6229 4928
rect 5909 4863 6229 4864
rect 15840 4928 16160 4929
rect 15840 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15840 4863 16160 4864
rect 25770 4928 26090 4929
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26090 4928
rect 25770 4863 26090 4864
rect 28165 4858 28231 4861
rect 31200 4858 32000 4888
rect 28165 4856 32000 4858
rect 28165 4800 28170 4856
rect 28226 4800 32000 4856
rect 28165 4798 32000 4800
rect 28165 4795 28231 4798
rect 31200 4768 32000 4798
rect 28717 4724 28783 4725
rect 28717 4722 28764 4724
rect 28672 4720 28764 4722
rect 28672 4664 28722 4720
rect 28672 4662 28764 4664
rect 28717 4660 28764 4662
rect 28828 4660 28834 4724
rect 28717 4659 28783 4660
rect 27797 4450 27863 4453
rect 31200 4450 32000 4480
rect 27797 4448 32000 4450
rect 27797 4392 27802 4448
rect 27858 4392 32000 4448
rect 27797 4390 32000 4392
rect 27797 4387 27863 4390
rect 10874 4384 11194 4385
rect 0 4314 800 4344
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 10874 4319 11194 4320
rect 20805 4384 21125 4385
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 31200 4360 32000 4390
rect 20805 4319 21125 4320
rect 1577 4314 1643 4317
rect 0 4312 1643 4314
rect 0 4256 1582 4312
rect 1638 4256 1643 4312
rect 0 4254 1643 4256
rect 0 4224 800 4254
rect 1577 4251 1643 4254
rect 29821 4044 29887 4045
rect 29821 4042 29868 4044
rect 29776 4040 29868 4042
rect 29776 3984 29826 4040
rect 29776 3982 29868 3984
rect 29821 3980 29868 3982
rect 29932 3980 29938 4044
rect 29821 3979 29887 3980
rect 28165 3906 28231 3909
rect 31200 3906 32000 3936
rect 28165 3904 32000 3906
rect 28165 3848 28170 3904
rect 28226 3848 32000 3904
rect 28165 3846 32000 3848
rect 28165 3843 28231 3846
rect 5909 3840 6229 3841
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6229 3840
rect 5909 3775 6229 3776
rect 15840 3840 16160 3841
rect 15840 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15840 3775 16160 3776
rect 25770 3840 26090 3841
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26090 3840
rect 31200 3816 32000 3846
rect 25770 3775 26090 3776
rect 0 3634 800 3664
rect 1577 3634 1643 3637
rect 0 3632 1643 3634
rect 0 3576 1582 3632
rect 1638 3576 1643 3632
rect 0 3574 1643 3576
rect 0 3544 800 3574
rect 1577 3571 1643 3574
rect 28257 3498 28323 3501
rect 31200 3498 32000 3528
rect 28257 3496 32000 3498
rect 28257 3440 28262 3496
rect 28318 3440 32000 3496
rect 28257 3438 32000 3440
rect 28257 3435 28323 3438
rect 31200 3408 32000 3438
rect 10874 3296 11194 3297
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 3231 11194 3232
rect 20805 3296 21125 3297
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 3231 21125 3232
rect 0 2954 800 2984
rect 1577 2954 1643 2957
rect 0 2952 1643 2954
rect 0 2896 1582 2952
rect 1638 2896 1643 2952
rect 0 2894 1643 2896
rect 0 2864 800 2894
rect 1577 2891 1643 2894
rect 28901 2954 28967 2957
rect 31200 2954 32000 2984
rect 28901 2952 32000 2954
rect 28901 2896 28906 2952
rect 28962 2896 32000 2952
rect 28901 2894 32000 2896
rect 28901 2891 28967 2894
rect 31200 2864 32000 2894
rect 5909 2752 6229 2753
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6229 2752
rect 5909 2687 6229 2688
rect 15840 2752 16160 2753
rect 15840 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15840 2687 16160 2688
rect 25770 2752 26090 2753
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26090 2752
rect 25770 2687 26090 2688
rect 29729 2546 29795 2549
rect 31200 2546 32000 2576
rect 29729 2544 32000 2546
rect 29729 2488 29734 2544
rect 29790 2488 32000 2544
rect 29729 2486 32000 2488
rect 29729 2483 29795 2486
rect 31200 2456 32000 2486
rect 0 2274 800 2304
rect 2313 2274 2379 2277
rect 0 2272 2379 2274
rect 0 2216 2318 2272
rect 2374 2216 2379 2272
rect 0 2214 2379 2216
rect 0 2184 800 2214
rect 2313 2211 2379 2214
rect 10874 2208 11194 2209
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2143 11194 2144
rect 20805 2208 21125 2209
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 20805 2143 21125 2144
rect 28717 2002 28783 2005
rect 31200 2002 32000 2032
rect 28717 2000 32000 2002
rect 28717 1944 28722 2000
rect 28778 1944 32000 2000
rect 28717 1942 32000 1944
rect 28717 1939 28783 1942
rect 31200 1912 32000 1942
rect 0 1594 800 1624
rect 1393 1594 1459 1597
rect 0 1592 1459 1594
rect 0 1536 1398 1592
rect 1454 1536 1459 1592
rect 0 1534 1459 1536
rect 0 1504 800 1534
rect 1393 1531 1459 1534
rect 28809 1594 28875 1597
rect 31200 1594 32000 1624
rect 28809 1592 32000 1594
rect 28809 1536 28814 1592
rect 28870 1536 32000 1592
rect 28809 1534 32000 1536
rect 28809 1531 28875 1534
rect 31200 1504 32000 1534
rect 29637 1050 29703 1053
rect 31200 1050 32000 1080
rect 29637 1048 32000 1050
rect 29637 992 29642 1048
rect 29698 992 32000 1048
rect 29637 990 32000 992
rect 29637 987 29703 990
rect 31200 960 32000 990
rect 0 914 800 944
rect 1577 914 1643 917
rect 0 912 1643 914
rect 0 856 1582 912
rect 1638 856 1643 912
rect 0 854 1643 856
rect 0 824 800 854
rect 1577 851 1643 854
rect 28717 642 28783 645
rect 31200 642 32000 672
rect 28717 640 32000 642
rect 28717 584 28722 640
rect 28778 584 32000 640
rect 28717 582 32000 584
rect 28717 579 28783 582
rect 31200 552 32000 582
rect 0 370 800 400
rect 2865 370 2931 373
rect 0 368 2931 370
rect 0 312 2870 368
rect 2926 312 2931 368
rect 0 310 2931 312
rect 0 280 800 310
rect 2865 307 2931 310
rect 28257 234 28323 237
rect 31200 234 32000 264
rect 28257 232 32000 234
rect 28257 176 28262 232
rect 28318 176 32000 232
rect 28257 174 32000 176
rect 28257 171 28323 174
rect 31200 144 32000 174
<< via3 >>
rect 5917 77820 5981 77824
rect 5917 77764 5921 77820
rect 5921 77764 5977 77820
rect 5977 77764 5981 77820
rect 5917 77760 5981 77764
rect 5997 77820 6061 77824
rect 5997 77764 6001 77820
rect 6001 77764 6057 77820
rect 6057 77764 6061 77820
rect 5997 77760 6061 77764
rect 6077 77820 6141 77824
rect 6077 77764 6081 77820
rect 6081 77764 6137 77820
rect 6137 77764 6141 77820
rect 6077 77760 6141 77764
rect 6157 77820 6221 77824
rect 6157 77764 6161 77820
rect 6161 77764 6217 77820
rect 6217 77764 6221 77820
rect 6157 77760 6221 77764
rect 15848 77820 15912 77824
rect 15848 77764 15852 77820
rect 15852 77764 15908 77820
rect 15908 77764 15912 77820
rect 15848 77760 15912 77764
rect 15928 77820 15992 77824
rect 15928 77764 15932 77820
rect 15932 77764 15988 77820
rect 15988 77764 15992 77820
rect 15928 77760 15992 77764
rect 16008 77820 16072 77824
rect 16008 77764 16012 77820
rect 16012 77764 16068 77820
rect 16068 77764 16072 77820
rect 16008 77760 16072 77764
rect 16088 77820 16152 77824
rect 16088 77764 16092 77820
rect 16092 77764 16148 77820
rect 16148 77764 16152 77820
rect 16088 77760 16152 77764
rect 25778 77820 25842 77824
rect 25778 77764 25782 77820
rect 25782 77764 25838 77820
rect 25838 77764 25842 77820
rect 25778 77760 25842 77764
rect 25858 77820 25922 77824
rect 25858 77764 25862 77820
rect 25862 77764 25918 77820
rect 25918 77764 25922 77820
rect 25858 77760 25922 77764
rect 25938 77820 26002 77824
rect 25938 77764 25942 77820
rect 25942 77764 25998 77820
rect 25998 77764 26002 77820
rect 25938 77760 26002 77764
rect 26018 77820 26082 77824
rect 26018 77764 26022 77820
rect 26022 77764 26078 77820
rect 26078 77764 26082 77820
rect 26018 77760 26082 77764
rect 10882 77276 10946 77280
rect 10882 77220 10886 77276
rect 10886 77220 10942 77276
rect 10942 77220 10946 77276
rect 10882 77216 10946 77220
rect 10962 77276 11026 77280
rect 10962 77220 10966 77276
rect 10966 77220 11022 77276
rect 11022 77220 11026 77276
rect 10962 77216 11026 77220
rect 11042 77276 11106 77280
rect 11042 77220 11046 77276
rect 11046 77220 11102 77276
rect 11102 77220 11106 77276
rect 11042 77216 11106 77220
rect 11122 77276 11186 77280
rect 11122 77220 11126 77276
rect 11126 77220 11182 77276
rect 11182 77220 11186 77276
rect 11122 77216 11186 77220
rect 20813 77276 20877 77280
rect 20813 77220 20817 77276
rect 20817 77220 20873 77276
rect 20873 77220 20877 77276
rect 20813 77216 20877 77220
rect 20893 77276 20957 77280
rect 20893 77220 20897 77276
rect 20897 77220 20953 77276
rect 20953 77220 20957 77276
rect 20893 77216 20957 77220
rect 20973 77276 21037 77280
rect 20973 77220 20977 77276
rect 20977 77220 21033 77276
rect 21033 77220 21037 77276
rect 20973 77216 21037 77220
rect 21053 77276 21117 77280
rect 21053 77220 21057 77276
rect 21057 77220 21113 77276
rect 21113 77220 21117 77276
rect 21053 77216 21117 77220
rect 5917 76732 5981 76736
rect 5917 76676 5921 76732
rect 5921 76676 5977 76732
rect 5977 76676 5981 76732
rect 5917 76672 5981 76676
rect 5997 76732 6061 76736
rect 5997 76676 6001 76732
rect 6001 76676 6057 76732
rect 6057 76676 6061 76732
rect 5997 76672 6061 76676
rect 6077 76732 6141 76736
rect 6077 76676 6081 76732
rect 6081 76676 6137 76732
rect 6137 76676 6141 76732
rect 6077 76672 6141 76676
rect 6157 76732 6221 76736
rect 6157 76676 6161 76732
rect 6161 76676 6217 76732
rect 6217 76676 6221 76732
rect 6157 76672 6221 76676
rect 15848 76732 15912 76736
rect 15848 76676 15852 76732
rect 15852 76676 15908 76732
rect 15908 76676 15912 76732
rect 15848 76672 15912 76676
rect 15928 76732 15992 76736
rect 15928 76676 15932 76732
rect 15932 76676 15988 76732
rect 15988 76676 15992 76732
rect 15928 76672 15992 76676
rect 16008 76732 16072 76736
rect 16008 76676 16012 76732
rect 16012 76676 16068 76732
rect 16068 76676 16072 76732
rect 16008 76672 16072 76676
rect 16088 76732 16152 76736
rect 16088 76676 16092 76732
rect 16092 76676 16148 76732
rect 16148 76676 16152 76732
rect 16088 76672 16152 76676
rect 25778 76732 25842 76736
rect 25778 76676 25782 76732
rect 25782 76676 25838 76732
rect 25838 76676 25842 76732
rect 25778 76672 25842 76676
rect 25858 76732 25922 76736
rect 25858 76676 25862 76732
rect 25862 76676 25918 76732
rect 25918 76676 25922 76732
rect 25858 76672 25922 76676
rect 25938 76732 26002 76736
rect 25938 76676 25942 76732
rect 25942 76676 25998 76732
rect 25998 76676 26002 76732
rect 25938 76672 26002 76676
rect 26018 76732 26082 76736
rect 26018 76676 26022 76732
rect 26022 76676 26078 76732
rect 26078 76676 26082 76732
rect 26018 76672 26082 76676
rect 10882 76188 10946 76192
rect 10882 76132 10886 76188
rect 10886 76132 10942 76188
rect 10942 76132 10946 76188
rect 10882 76128 10946 76132
rect 10962 76188 11026 76192
rect 10962 76132 10966 76188
rect 10966 76132 11022 76188
rect 11022 76132 11026 76188
rect 10962 76128 11026 76132
rect 11042 76188 11106 76192
rect 11042 76132 11046 76188
rect 11046 76132 11102 76188
rect 11102 76132 11106 76188
rect 11042 76128 11106 76132
rect 11122 76188 11186 76192
rect 11122 76132 11126 76188
rect 11126 76132 11182 76188
rect 11182 76132 11186 76188
rect 11122 76128 11186 76132
rect 20813 76188 20877 76192
rect 20813 76132 20817 76188
rect 20817 76132 20873 76188
rect 20873 76132 20877 76188
rect 20813 76128 20877 76132
rect 20893 76188 20957 76192
rect 20893 76132 20897 76188
rect 20897 76132 20953 76188
rect 20953 76132 20957 76188
rect 20893 76128 20957 76132
rect 20973 76188 21037 76192
rect 20973 76132 20977 76188
rect 20977 76132 21033 76188
rect 21033 76132 21037 76188
rect 20973 76128 21037 76132
rect 21053 76188 21117 76192
rect 21053 76132 21057 76188
rect 21057 76132 21113 76188
rect 21113 76132 21117 76188
rect 21053 76128 21117 76132
rect 5917 75644 5981 75648
rect 5917 75588 5921 75644
rect 5921 75588 5977 75644
rect 5977 75588 5981 75644
rect 5917 75584 5981 75588
rect 5997 75644 6061 75648
rect 5997 75588 6001 75644
rect 6001 75588 6057 75644
rect 6057 75588 6061 75644
rect 5997 75584 6061 75588
rect 6077 75644 6141 75648
rect 6077 75588 6081 75644
rect 6081 75588 6137 75644
rect 6137 75588 6141 75644
rect 6077 75584 6141 75588
rect 6157 75644 6221 75648
rect 6157 75588 6161 75644
rect 6161 75588 6217 75644
rect 6217 75588 6221 75644
rect 6157 75584 6221 75588
rect 15848 75644 15912 75648
rect 15848 75588 15852 75644
rect 15852 75588 15908 75644
rect 15908 75588 15912 75644
rect 15848 75584 15912 75588
rect 15928 75644 15992 75648
rect 15928 75588 15932 75644
rect 15932 75588 15988 75644
rect 15988 75588 15992 75644
rect 15928 75584 15992 75588
rect 16008 75644 16072 75648
rect 16008 75588 16012 75644
rect 16012 75588 16068 75644
rect 16068 75588 16072 75644
rect 16008 75584 16072 75588
rect 16088 75644 16152 75648
rect 16088 75588 16092 75644
rect 16092 75588 16148 75644
rect 16148 75588 16152 75644
rect 16088 75584 16152 75588
rect 25778 75644 25842 75648
rect 25778 75588 25782 75644
rect 25782 75588 25838 75644
rect 25838 75588 25842 75644
rect 25778 75584 25842 75588
rect 25858 75644 25922 75648
rect 25858 75588 25862 75644
rect 25862 75588 25918 75644
rect 25918 75588 25922 75644
rect 25858 75584 25922 75588
rect 25938 75644 26002 75648
rect 25938 75588 25942 75644
rect 25942 75588 25998 75644
rect 25998 75588 26002 75644
rect 25938 75584 26002 75588
rect 26018 75644 26082 75648
rect 26018 75588 26022 75644
rect 26022 75588 26078 75644
rect 26078 75588 26082 75644
rect 26018 75584 26082 75588
rect 10882 75100 10946 75104
rect 10882 75044 10886 75100
rect 10886 75044 10942 75100
rect 10942 75044 10946 75100
rect 10882 75040 10946 75044
rect 10962 75100 11026 75104
rect 10962 75044 10966 75100
rect 10966 75044 11022 75100
rect 11022 75044 11026 75100
rect 10962 75040 11026 75044
rect 11042 75100 11106 75104
rect 11042 75044 11046 75100
rect 11046 75044 11102 75100
rect 11102 75044 11106 75100
rect 11042 75040 11106 75044
rect 11122 75100 11186 75104
rect 11122 75044 11126 75100
rect 11126 75044 11182 75100
rect 11182 75044 11186 75100
rect 11122 75040 11186 75044
rect 20813 75100 20877 75104
rect 20813 75044 20817 75100
rect 20817 75044 20873 75100
rect 20873 75044 20877 75100
rect 20813 75040 20877 75044
rect 20893 75100 20957 75104
rect 20893 75044 20897 75100
rect 20897 75044 20953 75100
rect 20953 75044 20957 75100
rect 20893 75040 20957 75044
rect 20973 75100 21037 75104
rect 20973 75044 20977 75100
rect 20977 75044 21033 75100
rect 21033 75044 21037 75100
rect 20973 75040 21037 75044
rect 21053 75100 21117 75104
rect 21053 75044 21057 75100
rect 21057 75044 21113 75100
rect 21113 75044 21117 75100
rect 21053 75040 21117 75044
rect 5917 74556 5981 74560
rect 5917 74500 5921 74556
rect 5921 74500 5977 74556
rect 5977 74500 5981 74556
rect 5917 74496 5981 74500
rect 5997 74556 6061 74560
rect 5997 74500 6001 74556
rect 6001 74500 6057 74556
rect 6057 74500 6061 74556
rect 5997 74496 6061 74500
rect 6077 74556 6141 74560
rect 6077 74500 6081 74556
rect 6081 74500 6137 74556
rect 6137 74500 6141 74556
rect 6077 74496 6141 74500
rect 6157 74556 6221 74560
rect 6157 74500 6161 74556
rect 6161 74500 6217 74556
rect 6217 74500 6221 74556
rect 6157 74496 6221 74500
rect 15848 74556 15912 74560
rect 15848 74500 15852 74556
rect 15852 74500 15908 74556
rect 15908 74500 15912 74556
rect 15848 74496 15912 74500
rect 15928 74556 15992 74560
rect 15928 74500 15932 74556
rect 15932 74500 15988 74556
rect 15988 74500 15992 74556
rect 15928 74496 15992 74500
rect 16008 74556 16072 74560
rect 16008 74500 16012 74556
rect 16012 74500 16068 74556
rect 16068 74500 16072 74556
rect 16008 74496 16072 74500
rect 16088 74556 16152 74560
rect 16088 74500 16092 74556
rect 16092 74500 16148 74556
rect 16148 74500 16152 74556
rect 16088 74496 16152 74500
rect 25778 74556 25842 74560
rect 25778 74500 25782 74556
rect 25782 74500 25838 74556
rect 25838 74500 25842 74556
rect 25778 74496 25842 74500
rect 25858 74556 25922 74560
rect 25858 74500 25862 74556
rect 25862 74500 25918 74556
rect 25918 74500 25922 74556
rect 25858 74496 25922 74500
rect 25938 74556 26002 74560
rect 25938 74500 25942 74556
rect 25942 74500 25998 74556
rect 25998 74500 26002 74556
rect 25938 74496 26002 74500
rect 26018 74556 26082 74560
rect 26018 74500 26022 74556
rect 26022 74500 26078 74556
rect 26078 74500 26082 74556
rect 26018 74496 26082 74500
rect 10882 74012 10946 74016
rect 10882 73956 10886 74012
rect 10886 73956 10942 74012
rect 10942 73956 10946 74012
rect 10882 73952 10946 73956
rect 10962 74012 11026 74016
rect 10962 73956 10966 74012
rect 10966 73956 11022 74012
rect 11022 73956 11026 74012
rect 10962 73952 11026 73956
rect 11042 74012 11106 74016
rect 11042 73956 11046 74012
rect 11046 73956 11102 74012
rect 11102 73956 11106 74012
rect 11042 73952 11106 73956
rect 11122 74012 11186 74016
rect 11122 73956 11126 74012
rect 11126 73956 11182 74012
rect 11182 73956 11186 74012
rect 11122 73952 11186 73956
rect 20813 74012 20877 74016
rect 20813 73956 20817 74012
rect 20817 73956 20873 74012
rect 20873 73956 20877 74012
rect 20813 73952 20877 73956
rect 20893 74012 20957 74016
rect 20893 73956 20897 74012
rect 20897 73956 20953 74012
rect 20953 73956 20957 74012
rect 20893 73952 20957 73956
rect 20973 74012 21037 74016
rect 20973 73956 20977 74012
rect 20977 73956 21033 74012
rect 21033 73956 21037 74012
rect 20973 73952 21037 73956
rect 21053 74012 21117 74016
rect 21053 73956 21057 74012
rect 21057 73956 21113 74012
rect 21113 73956 21117 74012
rect 21053 73952 21117 73956
rect 5917 73468 5981 73472
rect 5917 73412 5921 73468
rect 5921 73412 5977 73468
rect 5977 73412 5981 73468
rect 5917 73408 5981 73412
rect 5997 73468 6061 73472
rect 5997 73412 6001 73468
rect 6001 73412 6057 73468
rect 6057 73412 6061 73468
rect 5997 73408 6061 73412
rect 6077 73468 6141 73472
rect 6077 73412 6081 73468
rect 6081 73412 6137 73468
rect 6137 73412 6141 73468
rect 6077 73408 6141 73412
rect 6157 73468 6221 73472
rect 6157 73412 6161 73468
rect 6161 73412 6217 73468
rect 6217 73412 6221 73468
rect 6157 73408 6221 73412
rect 15848 73468 15912 73472
rect 15848 73412 15852 73468
rect 15852 73412 15908 73468
rect 15908 73412 15912 73468
rect 15848 73408 15912 73412
rect 15928 73468 15992 73472
rect 15928 73412 15932 73468
rect 15932 73412 15988 73468
rect 15988 73412 15992 73468
rect 15928 73408 15992 73412
rect 16008 73468 16072 73472
rect 16008 73412 16012 73468
rect 16012 73412 16068 73468
rect 16068 73412 16072 73468
rect 16008 73408 16072 73412
rect 16088 73468 16152 73472
rect 16088 73412 16092 73468
rect 16092 73412 16148 73468
rect 16148 73412 16152 73468
rect 16088 73408 16152 73412
rect 25778 73468 25842 73472
rect 25778 73412 25782 73468
rect 25782 73412 25838 73468
rect 25838 73412 25842 73468
rect 25778 73408 25842 73412
rect 25858 73468 25922 73472
rect 25858 73412 25862 73468
rect 25862 73412 25918 73468
rect 25918 73412 25922 73468
rect 25858 73408 25922 73412
rect 25938 73468 26002 73472
rect 25938 73412 25942 73468
rect 25942 73412 25998 73468
rect 25998 73412 26002 73468
rect 25938 73408 26002 73412
rect 26018 73468 26082 73472
rect 26018 73412 26022 73468
rect 26022 73412 26078 73468
rect 26078 73412 26082 73468
rect 26018 73408 26082 73412
rect 10882 72924 10946 72928
rect 10882 72868 10886 72924
rect 10886 72868 10942 72924
rect 10942 72868 10946 72924
rect 10882 72864 10946 72868
rect 10962 72924 11026 72928
rect 10962 72868 10966 72924
rect 10966 72868 11022 72924
rect 11022 72868 11026 72924
rect 10962 72864 11026 72868
rect 11042 72924 11106 72928
rect 11042 72868 11046 72924
rect 11046 72868 11102 72924
rect 11102 72868 11106 72924
rect 11042 72864 11106 72868
rect 11122 72924 11186 72928
rect 11122 72868 11126 72924
rect 11126 72868 11182 72924
rect 11182 72868 11186 72924
rect 11122 72864 11186 72868
rect 20813 72924 20877 72928
rect 20813 72868 20817 72924
rect 20817 72868 20873 72924
rect 20873 72868 20877 72924
rect 20813 72864 20877 72868
rect 20893 72924 20957 72928
rect 20893 72868 20897 72924
rect 20897 72868 20953 72924
rect 20953 72868 20957 72924
rect 20893 72864 20957 72868
rect 20973 72924 21037 72928
rect 20973 72868 20977 72924
rect 20977 72868 21033 72924
rect 21033 72868 21037 72924
rect 20973 72864 21037 72868
rect 21053 72924 21117 72928
rect 21053 72868 21057 72924
rect 21057 72868 21113 72924
rect 21113 72868 21117 72924
rect 21053 72864 21117 72868
rect 5917 72380 5981 72384
rect 5917 72324 5921 72380
rect 5921 72324 5977 72380
rect 5977 72324 5981 72380
rect 5917 72320 5981 72324
rect 5997 72380 6061 72384
rect 5997 72324 6001 72380
rect 6001 72324 6057 72380
rect 6057 72324 6061 72380
rect 5997 72320 6061 72324
rect 6077 72380 6141 72384
rect 6077 72324 6081 72380
rect 6081 72324 6137 72380
rect 6137 72324 6141 72380
rect 6077 72320 6141 72324
rect 6157 72380 6221 72384
rect 6157 72324 6161 72380
rect 6161 72324 6217 72380
rect 6217 72324 6221 72380
rect 6157 72320 6221 72324
rect 15848 72380 15912 72384
rect 15848 72324 15852 72380
rect 15852 72324 15908 72380
rect 15908 72324 15912 72380
rect 15848 72320 15912 72324
rect 15928 72380 15992 72384
rect 15928 72324 15932 72380
rect 15932 72324 15988 72380
rect 15988 72324 15992 72380
rect 15928 72320 15992 72324
rect 16008 72380 16072 72384
rect 16008 72324 16012 72380
rect 16012 72324 16068 72380
rect 16068 72324 16072 72380
rect 16008 72320 16072 72324
rect 16088 72380 16152 72384
rect 16088 72324 16092 72380
rect 16092 72324 16148 72380
rect 16148 72324 16152 72380
rect 16088 72320 16152 72324
rect 25778 72380 25842 72384
rect 25778 72324 25782 72380
rect 25782 72324 25838 72380
rect 25838 72324 25842 72380
rect 25778 72320 25842 72324
rect 25858 72380 25922 72384
rect 25858 72324 25862 72380
rect 25862 72324 25918 72380
rect 25918 72324 25922 72380
rect 25858 72320 25922 72324
rect 25938 72380 26002 72384
rect 25938 72324 25942 72380
rect 25942 72324 25998 72380
rect 25998 72324 26002 72380
rect 25938 72320 26002 72324
rect 26018 72380 26082 72384
rect 26018 72324 26022 72380
rect 26022 72324 26078 72380
rect 26078 72324 26082 72380
rect 26018 72320 26082 72324
rect 10882 71836 10946 71840
rect 10882 71780 10886 71836
rect 10886 71780 10942 71836
rect 10942 71780 10946 71836
rect 10882 71776 10946 71780
rect 10962 71836 11026 71840
rect 10962 71780 10966 71836
rect 10966 71780 11022 71836
rect 11022 71780 11026 71836
rect 10962 71776 11026 71780
rect 11042 71836 11106 71840
rect 11042 71780 11046 71836
rect 11046 71780 11102 71836
rect 11102 71780 11106 71836
rect 11042 71776 11106 71780
rect 11122 71836 11186 71840
rect 11122 71780 11126 71836
rect 11126 71780 11182 71836
rect 11182 71780 11186 71836
rect 11122 71776 11186 71780
rect 20813 71836 20877 71840
rect 20813 71780 20817 71836
rect 20817 71780 20873 71836
rect 20873 71780 20877 71836
rect 20813 71776 20877 71780
rect 20893 71836 20957 71840
rect 20893 71780 20897 71836
rect 20897 71780 20953 71836
rect 20953 71780 20957 71836
rect 20893 71776 20957 71780
rect 20973 71836 21037 71840
rect 20973 71780 20977 71836
rect 20977 71780 21033 71836
rect 21033 71780 21037 71836
rect 20973 71776 21037 71780
rect 21053 71836 21117 71840
rect 21053 71780 21057 71836
rect 21057 71780 21113 71836
rect 21113 71780 21117 71836
rect 21053 71776 21117 71780
rect 5917 71292 5981 71296
rect 5917 71236 5921 71292
rect 5921 71236 5977 71292
rect 5977 71236 5981 71292
rect 5917 71232 5981 71236
rect 5997 71292 6061 71296
rect 5997 71236 6001 71292
rect 6001 71236 6057 71292
rect 6057 71236 6061 71292
rect 5997 71232 6061 71236
rect 6077 71292 6141 71296
rect 6077 71236 6081 71292
rect 6081 71236 6137 71292
rect 6137 71236 6141 71292
rect 6077 71232 6141 71236
rect 6157 71292 6221 71296
rect 6157 71236 6161 71292
rect 6161 71236 6217 71292
rect 6217 71236 6221 71292
rect 6157 71232 6221 71236
rect 15848 71292 15912 71296
rect 15848 71236 15852 71292
rect 15852 71236 15908 71292
rect 15908 71236 15912 71292
rect 15848 71232 15912 71236
rect 15928 71292 15992 71296
rect 15928 71236 15932 71292
rect 15932 71236 15988 71292
rect 15988 71236 15992 71292
rect 15928 71232 15992 71236
rect 16008 71292 16072 71296
rect 16008 71236 16012 71292
rect 16012 71236 16068 71292
rect 16068 71236 16072 71292
rect 16008 71232 16072 71236
rect 16088 71292 16152 71296
rect 16088 71236 16092 71292
rect 16092 71236 16148 71292
rect 16148 71236 16152 71292
rect 16088 71232 16152 71236
rect 25778 71292 25842 71296
rect 25778 71236 25782 71292
rect 25782 71236 25838 71292
rect 25838 71236 25842 71292
rect 25778 71232 25842 71236
rect 25858 71292 25922 71296
rect 25858 71236 25862 71292
rect 25862 71236 25918 71292
rect 25918 71236 25922 71292
rect 25858 71232 25922 71236
rect 25938 71292 26002 71296
rect 25938 71236 25942 71292
rect 25942 71236 25998 71292
rect 25998 71236 26002 71292
rect 25938 71232 26002 71236
rect 26018 71292 26082 71296
rect 26018 71236 26022 71292
rect 26022 71236 26078 71292
rect 26078 71236 26082 71292
rect 26018 71232 26082 71236
rect 10882 70748 10946 70752
rect 10882 70692 10886 70748
rect 10886 70692 10942 70748
rect 10942 70692 10946 70748
rect 10882 70688 10946 70692
rect 10962 70748 11026 70752
rect 10962 70692 10966 70748
rect 10966 70692 11022 70748
rect 11022 70692 11026 70748
rect 10962 70688 11026 70692
rect 11042 70748 11106 70752
rect 11042 70692 11046 70748
rect 11046 70692 11102 70748
rect 11102 70692 11106 70748
rect 11042 70688 11106 70692
rect 11122 70748 11186 70752
rect 11122 70692 11126 70748
rect 11126 70692 11182 70748
rect 11182 70692 11186 70748
rect 11122 70688 11186 70692
rect 20813 70748 20877 70752
rect 20813 70692 20817 70748
rect 20817 70692 20873 70748
rect 20873 70692 20877 70748
rect 20813 70688 20877 70692
rect 20893 70748 20957 70752
rect 20893 70692 20897 70748
rect 20897 70692 20953 70748
rect 20953 70692 20957 70748
rect 20893 70688 20957 70692
rect 20973 70748 21037 70752
rect 20973 70692 20977 70748
rect 20977 70692 21033 70748
rect 21033 70692 21037 70748
rect 20973 70688 21037 70692
rect 21053 70748 21117 70752
rect 21053 70692 21057 70748
rect 21057 70692 21113 70748
rect 21113 70692 21117 70748
rect 21053 70688 21117 70692
rect 5917 70204 5981 70208
rect 5917 70148 5921 70204
rect 5921 70148 5977 70204
rect 5977 70148 5981 70204
rect 5917 70144 5981 70148
rect 5997 70204 6061 70208
rect 5997 70148 6001 70204
rect 6001 70148 6057 70204
rect 6057 70148 6061 70204
rect 5997 70144 6061 70148
rect 6077 70204 6141 70208
rect 6077 70148 6081 70204
rect 6081 70148 6137 70204
rect 6137 70148 6141 70204
rect 6077 70144 6141 70148
rect 6157 70204 6221 70208
rect 6157 70148 6161 70204
rect 6161 70148 6217 70204
rect 6217 70148 6221 70204
rect 6157 70144 6221 70148
rect 15848 70204 15912 70208
rect 15848 70148 15852 70204
rect 15852 70148 15908 70204
rect 15908 70148 15912 70204
rect 15848 70144 15912 70148
rect 15928 70204 15992 70208
rect 15928 70148 15932 70204
rect 15932 70148 15988 70204
rect 15988 70148 15992 70204
rect 15928 70144 15992 70148
rect 16008 70204 16072 70208
rect 16008 70148 16012 70204
rect 16012 70148 16068 70204
rect 16068 70148 16072 70204
rect 16008 70144 16072 70148
rect 16088 70204 16152 70208
rect 16088 70148 16092 70204
rect 16092 70148 16148 70204
rect 16148 70148 16152 70204
rect 16088 70144 16152 70148
rect 25778 70204 25842 70208
rect 25778 70148 25782 70204
rect 25782 70148 25838 70204
rect 25838 70148 25842 70204
rect 25778 70144 25842 70148
rect 25858 70204 25922 70208
rect 25858 70148 25862 70204
rect 25862 70148 25918 70204
rect 25918 70148 25922 70204
rect 25858 70144 25922 70148
rect 25938 70204 26002 70208
rect 25938 70148 25942 70204
rect 25942 70148 25998 70204
rect 25998 70148 26002 70204
rect 25938 70144 26002 70148
rect 26018 70204 26082 70208
rect 26018 70148 26022 70204
rect 26022 70148 26078 70204
rect 26078 70148 26082 70204
rect 26018 70144 26082 70148
rect 29132 70000 29196 70004
rect 29132 69944 29182 70000
rect 29182 69944 29196 70000
rect 29132 69940 29196 69944
rect 10882 69660 10946 69664
rect 10882 69604 10886 69660
rect 10886 69604 10942 69660
rect 10942 69604 10946 69660
rect 10882 69600 10946 69604
rect 10962 69660 11026 69664
rect 10962 69604 10966 69660
rect 10966 69604 11022 69660
rect 11022 69604 11026 69660
rect 10962 69600 11026 69604
rect 11042 69660 11106 69664
rect 11042 69604 11046 69660
rect 11046 69604 11102 69660
rect 11102 69604 11106 69660
rect 11042 69600 11106 69604
rect 11122 69660 11186 69664
rect 11122 69604 11126 69660
rect 11126 69604 11182 69660
rect 11182 69604 11186 69660
rect 11122 69600 11186 69604
rect 20813 69660 20877 69664
rect 20813 69604 20817 69660
rect 20817 69604 20873 69660
rect 20873 69604 20877 69660
rect 20813 69600 20877 69604
rect 20893 69660 20957 69664
rect 20893 69604 20897 69660
rect 20897 69604 20953 69660
rect 20953 69604 20957 69660
rect 20893 69600 20957 69604
rect 20973 69660 21037 69664
rect 20973 69604 20977 69660
rect 20977 69604 21033 69660
rect 21033 69604 21037 69660
rect 20973 69600 21037 69604
rect 21053 69660 21117 69664
rect 21053 69604 21057 69660
rect 21057 69604 21113 69660
rect 21113 69604 21117 69660
rect 21053 69600 21117 69604
rect 5917 69116 5981 69120
rect 5917 69060 5921 69116
rect 5921 69060 5977 69116
rect 5977 69060 5981 69116
rect 5917 69056 5981 69060
rect 5997 69116 6061 69120
rect 5997 69060 6001 69116
rect 6001 69060 6057 69116
rect 6057 69060 6061 69116
rect 5997 69056 6061 69060
rect 6077 69116 6141 69120
rect 6077 69060 6081 69116
rect 6081 69060 6137 69116
rect 6137 69060 6141 69116
rect 6077 69056 6141 69060
rect 6157 69116 6221 69120
rect 6157 69060 6161 69116
rect 6161 69060 6217 69116
rect 6217 69060 6221 69116
rect 6157 69056 6221 69060
rect 15848 69116 15912 69120
rect 15848 69060 15852 69116
rect 15852 69060 15908 69116
rect 15908 69060 15912 69116
rect 15848 69056 15912 69060
rect 15928 69116 15992 69120
rect 15928 69060 15932 69116
rect 15932 69060 15988 69116
rect 15988 69060 15992 69116
rect 15928 69056 15992 69060
rect 16008 69116 16072 69120
rect 16008 69060 16012 69116
rect 16012 69060 16068 69116
rect 16068 69060 16072 69116
rect 16008 69056 16072 69060
rect 16088 69116 16152 69120
rect 16088 69060 16092 69116
rect 16092 69060 16148 69116
rect 16148 69060 16152 69116
rect 16088 69056 16152 69060
rect 25778 69116 25842 69120
rect 25778 69060 25782 69116
rect 25782 69060 25838 69116
rect 25838 69060 25842 69116
rect 25778 69056 25842 69060
rect 25858 69116 25922 69120
rect 25858 69060 25862 69116
rect 25862 69060 25918 69116
rect 25918 69060 25922 69116
rect 25858 69056 25922 69060
rect 25938 69116 26002 69120
rect 25938 69060 25942 69116
rect 25942 69060 25998 69116
rect 25998 69060 26002 69116
rect 25938 69056 26002 69060
rect 26018 69116 26082 69120
rect 26018 69060 26022 69116
rect 26022 69060 26078 69116
rect 26078 69060 26082 69116
rect 26018 69056 26082 69060
rect 10882 68572 10946 68576
rect 10882 68516 10886 68572
rect 10886 68516 10942 68572
rect 10942 68516 10946 68572
rect 10882 68512 10946 68516
rect 10962 68572 11026 68576
rect 10962 68516 10966 68572
rect 10966 68516 11022 68572
rect 11022 68516 11026 68572
rect 10962 68512 11026 68516
rect 11042 68572 11106 68576
rect 11042 68516 11046 68572
rect 11046 68516 11102 68572
rect 11102 68516 11106 68572
rect 11042 68512 11106 68516
rect 11122 68572 11186 68576
rect 11122 68516 11126 68572
rect 11126 68516 11182 68572
rect 11182 68516 11186 68572
rect 11122 68512 11186 68516
rect 20813 68572 20877 68576
rect 20813 68516 20817 68572
rect 20817 68516 20873 68572
rect 20873 68516 20877 68572
rect 20813 68512 20877 68516
rect 20893 68572 20957 68576
rect 20893 68516 20897 68572
rect 20897 68516 20953 68572
rect 20953 68516 20957 68572
rect 20893 68512 20957 68516
rect 20973 68572 21037 68576
rect 20973 68516 20977 68572
rect 20977 68516 21033 68572
rect 21033 68516 21037 68572
rect 20973 68512 21037 68516
rect 21053 68572 21117 68576
rect 21053 68516 21057 68572
rect 21057 68516 21113 68572
rect 21113 68516 21117 68572
rect 21053 68512 21117 68516
rect 5917 68028 5981 68032
rect 5917 67972 5921 68028
rect 5921 67972 5977 68028
rect 5977 67972 5981 68028
rect 5917 67968 5981 67972
rect 5997 68028 6061 68032
rect 5997 67972 6001 68028
rect 6001 67972 6057 68028
rect 6057 67972 6061 68028
rect 5997 67968 6061 67972
rect 6077 68028 6141 68032
rect 6077 67972 6081 68028
rect 6081 67972 6137 68028
rect 6137 67972 6141 68028
rect 6077 67968 6141 67972
rect 6157 68028 6221 68032
rect 6157 67972 6161 68028
rect 6161 67972 6217 68028
rect 6217 67972 6221 68028
rect 6157 67968 6221 67972
rect 15848 68028 15912 68032
rect 15848 67972 15852 68028
rect 15852 67972 15908 68028
rect 15908 67972 15912 68028
rect 15848 67968 15912 67972
rect 15928 68028 15992 68032
rect 15928 67972 15932 68028
rect 15932 67972 15988 68028
rect 15988 67972 15992 68028
rect 15928 67968 15992 67972
rect 16008 68028 16072 68032
rect 16008 67972 16012 68028
rect 16012 67972 16068 68028
rect 16068 67972 16072 68028
rect 16008 67968 16072 67972
rect 16088 68028 16152 68032
rect 16088 67972 16092 68028
rect 16092 67972 16148 68028
rect 16148 67972 16152 68028
rect 16088 67968 16152 67972
rect 25778 68028 25842 68032
rect 25778 67972 25782 68028
rect 25782 67972 25838 68028
rect 25838 67972 25842 68028
rect 25778 67968 25842 67972
rect 25858 68028 25922 68032
rect 25858 67972 25862 68028
rect 25862 67972 25918 68028
rect 25918 67972 25922 68028
rect 25858 67968 25922 67972
rect 25938 68028 26002 68032
rect 25938 67972 25942 68028
rect 25942 67972 25998 68028
rect 25998 67972 26002 68028
rect 25938 67968 26002 67972
rect 26018 68028 26082 68032
rect 26018 67972 26022 68028
rect 26022 67972 26078 68028
rect 26078 67972 26082 68028
rect 26018 67968 26082 67972
rect 27108 67492 27172 67556
rect 10882 67484 10946 67488
rect 10882 67428 10886 67484
rect 10886 67428 10942 67484
rect 10942 67428 10946 67484
rect 10882 67424 10946 67428
rect 10962 67484 11026 67488
rect 10962 67428 10966 67484
rect 10966 67428 11022 67484
rect 11022 67428 11026 67484
rect 10962 67424 11026 67428
rect 11042 67484 11106 67488
rect 11042 67428 11046 67484
rect 11046 67428 11102 67484
rect 11102 67428 11106 67484
rect 11042 67424 11106 67428
rect 11122 67484 11186 67488
rect 11122 67428 11126 67484
rect 11126 67428 11182 67484
rect 11182 67428 11186 67484
rect 11122 67424 11186 67428
rect 20813 67484 20877 67488
rect 20813 67428 20817 67484
rect 20817 67428 20873 67484
rect 20873 67428 20877 67484
rect 20813 67424 20877 67428
rect 20893 67484 20957 67488
rect 20893 67428 20897 67484
rect 20897 67428 20953 67484
rect 20953 67428 20957 67484
rect 20893 67424 20957 67428
rect 20973 67484 21037 67488
rect 20973 67428 20977 67484
rect 20977 67428 21033 67484
rect 21033 67428 21037 67484
rect 20973 67424 21037 67428
rect 21053 67484 21117 67488
rect 21053 67428 21057 67484
rect 21057 67428 21113 67484
rect 21113 67428 21117 67484
rect 21053 67424 21117 67428
rect 5917 66940 5981 66944
rect 5917 66884 5921 66940
rect 5921 66884 5977 66940
rect 5977 66884 5981 66940
rect 5917 66880 5981 66884
rect 5997 66940 6061 66944
rect 5997 66884 6001 66940
rect 6001 66884 6057 66940
rect 6057 66884 6061 66940
rect 5997 66880 6061 66884
rect 6077 66940 6141 66944
rect 6077 66884 6081 66940
rect 6081 66884 6137 66940
rect 6137 66884 6141 66940
rect 6077 66880 6141 66884
rect 6157 66940 6221 66944
rect 6157 66884 6161 66940
rect 6161 66884 6217 66940
rect 6217 66884 6221 66940
rect 6157 66880 6221 66884
rect 15848 66940 15912 66944
rect 15848 66884 15852 66940
rect 15852 66884 15908 66940
rect 15908 66884 15912 66940
rect 15848 66880 15912 66884
rect 15928 66940 15992 66944
rect 15928 66884 15932 66940
rect 15932 66884 15988 66940
rect 15988 66884 15992 66940
rect 15928 66880 15992 66884
rect 16008 66940 16072 66944
rect 16008 66884 16012 66940
rect 16012 66884 16068 66940
rect 16068 66884 16072 66940
rect 16008 66880 16072 66884
rect 16088 66940 16152 66944
rect 16088 66884 16092 66940
rect 16092 66884 16148 66940
rect 16148 66884 16152 66940
rect 16088 66880 16152 66884
rect 25778 66940 25842 66944
rect 25778 66884 25782 66940
rect 25782 66884 25838 66940
rect 25838 66884 25842 66940
rect 25778 66880 25842 66884
rect 25858 66940 25922 66944
rect 25858 66884 25862 66940
rect 25862 66884 25918 66940
rect 25918 66884 25922 66940
rect 25858 66880 25922 66884
rect 25938 66940 26002 66944
rect 25938 66884 25942 66940
rect 25942 66884 25998 66940
rect 25998 66884 26002 66940
rect 25938 66880 26002 66884
rect 26018 66940 26082 66944
rect 26018 66884 26022 66940
rect 26022 66884 26078 66940
rect 26078 66884 26082 66940
rect 26018 66880 26082 66884
rect 26372 66812 26436 66876
rect 10882 66396 10946 66400
rect 10882 66340 10886 66396
rect 10886 66340 10942 66396
rect 10942 66340 10946 66396
rect 10882 66336 10946 66340
rect 10962 66396 11026 66400
rect 10962 66340 10966 66396
rect 10966 66340 11022 66396
rect 11022 66340 11026 66396
rect 10962 66336 11026 66340
rect 11042 66396 11106 66400
rect 11042 66340 11046 66396
rect 11046 66340 11102 66396
rect 11102 66340 11106 66396
rect 11042 66336 11106 66340
rect 11122 66396 11186 66400
rect 11122 66340 11126 66396
rect 11126 66340 11182 66396
rect 11182 66340 11186 66396
rect 11122 66336 11186 66340
rect 20813 66396 20877 66400
rect 20813 66340 20817 66396
rect 20817 66340 20873 66396
rect 20873 66340 20877 66396
rect 20813 66336 20877 66340
rect 20893 66396 20957 66400
rect 20893 66340 20897 66396
rect 20897 66340 20953 66396
rect 20953 66340 20957 66396
rect 20893 66336 20957 66340
rect 20973 66396 21037 66400
rect 20973 66340 20977 66396
rect 20977 66340 21033 66396
rect 21033 66340 21037 66396
rect 20973 66336 21037 66340
rect 21053 66396 21117 66400
rect 21053 66340 21057 66396
rect 21057 66340 21113 66396
rect 21113 66340 21117 66396
rect 21053 66336 21117 66340
rect 25084 65996 25148 66060
rect 5917 65852 5981 65856
rect 5917 65796 5921 65852
rect 5921 65796 5977 65852
rect 5977 65796 5981 65852
rect 5917 65792 5981 65796
rect 5997 65852 6061 65856
rect 5997 65796 6001 65852
rect 6001 65796 6057 65852
rect 6057 65796 6061 65852
rect 5997 65792 6061 65796
rect 6077 65852 6141 65856
rect 6077 65796 6081 65852
rect 6081 65796 6137 65852
rect 6137 65796 6141 65852
rect 6077 65792 6141 65796
rect 6157 65852 6221 65856
rect 6157 65796 6161 65852
rect 6161 65796 6217 65852
rect 6217 65796 6221 65852
rect 6157 65792 6221 65796
rect 15848 65852 15912 65856
rect 15848 65796 15852 65852
rect 15852 65796 15908 65852
rect 15908 65796 15912 65852
rect 15848 65792 15912 65796
rect 15928 65852 15992 65856
rect 15928 65796 15932 65852
rect 15932 65796 15988 65852
rect 15988 65796 15992 65852
rect 15928 65792 15992 65796
rect 16008 65852 16072 65856
rect 16008 65796 16012 65852
rect 16012 65796 16068 65852
rect 16068 65796 16072 65852
rect 16008 65792 16072 65796
rect 16088 65852 16152 65856
rect 16088 65796 16092 65852
rect 16092 65796 16148 65852
rect 16148 65796 16152 65852
rect 16088 65792 16152 65796
rect 25778 65852 25842 65856
rect 25778 65796 25782 65852
rect 25782 65796 25838 65852
rect 25838 65796 25842 65852
rect 25778 65792 25842 65796
rect 25858 65852 25922 65856
rect 25858 65796 25862 65852
rect 25862 65796 25918 65852
rect 25918 65796 25922 65852
rect 25858 65792 25922 65796
rect 25938 65852 26002 65856
rect 25938 65796 25942 65852
rect 25942 65796 25998 65852
rect 25998 65796 26002 65852
rect 25938 65792 26002 65796
rect 26018 65852 26082 65856
rect 26018 65796 26022 65852
rect 26022 65796 26078 65852
rect 26078 65796 26082 65852
rect 26018 65792 26082 65796
rect 27660 65588 27724 65652
rect 28396 65648 28460 65652
rect 28396 65592 28446 65648
rect 28446 65592 28460 65648
rect 28396 65588 28460 65592
rect 10882 65308 10946 65312
rect 10882 65252 10886 65308
rect 10886 65252 10942 65308
rect 10942 65252 10946 65308
rect 10882 65248 10946 65252
rect 10962 65308 11026 65312
rect 10962 65252 10966 65308
rect 10966 65252 11022 65308
rect 11022 65252 11026 65308
rect 10962 65248 11026 65252
rect 11042 65308 11106 65312
rect 11042 65252 11046 65308
rect 11046 65252 11102 65308
rect 11102 65252 11106 65308
rect 11042 65248 11106 65252
rect 11122 65308 11186 65312
rect 11122 65252 11126 65308
rect 11126 65252 11182 65308
rect 11182 65252 11186 65308
rect 11122 65248 11186 65252
rect 20813 65308 20877 65312
rect 20813 65252 20817 65308
rect 20817 65252 20873 65308
rect 20873 65252 20877 65308
rect 20813 65248 20877 65252
rect 20893 65308 20957 65312
rect 20893 65252 20897 65308
rect 20897 65252 20953 65308
rect 20953 65252 20957 65308
rect 20893 65248 20957 65252
rect 20973 65308 21037 65312
rect 20973 65252 20977 65308
rect 20977 65252 21033 65308
rect 21033 65252 21037 65308
rect 20973 65248 21037 65252
rect 21053 65308 21117 65312
rect 21053 65252 21057 65308
rect 21057 65252 21113 65308
rect 21113 65252 21117 65308
rect 21053 65248 21117 65252
rect 28764 64908 28828 64972
rect 5917 64764 5981 64768
rect 5917 64708 5921 64764
rect 5921 64708 5977 64764
rect 5977 64708 5981 64764
rect 5917 64704 5981 64708
rect 5997 64764 6061 64768
rect 5997 64708 6001 64764
rect 6001 64708 6057 64764
rect 6057 64708 6061 64764
rect 5997 64704 6061 64708
rect 6077 64764 6141 64768
rect 6077 64708 6081 64764
rect 6081 64708 6137 64764
rect 6137 64708 6141 64764
rect 6077 64704 6141 64708
rect 6157 64764 6221 64768
rect 6157 64708 6161 64764
rect 6161 64708 6217 64764
rect 6217 64708 6221 64764
rect 6157 64704 6221 64708
rect 15848 64764 15912 64768
rect 15848 64708 15852 64764
rect 15852 64708 15908 64764
rect 15908 64708 15912 64764
rect 15848 64704 15912 64708
rect 15928 64764 15992 64768
rect 15928 64708 15932 64764
rect 15932 64708 15988 64764
rect 15988 64708 15992 64764
rect 15928 64704 15992 64708
rect 16008 64764 16072 64768
rect 16008 64708 16012 64764
rect 16012 64708 16068 64764
rect 16068 64708 16072 64764
rect 16008 64704 16072 64708
rect 16088 64764 16152 64768
rect 16088 64708 16092 64764
rect 16092 64708 16148 64764
rect 16148 64708 16152 64764
rect 16088 64704 16152 64708
rect 25778 64764 25842 64768
rect 25778 64708 25782 64764
rect 25782 64708 25838 64764
rect 25838 64708 25842 64764
rect 25778 64704 25842 64708
rect 25858 64764 25922 64768
rect 25858 64708 25862 64764
rect 25862 64708 25918 64764
rect 25918 64708 25922 64764
rect 25858 64704 25922 64708
rect 25938 64764 26002 64768
rect 25938 64708 25942 64764
rect 25942 64708 25998 64764
rect 25998 64708 26002 64764
rect 25938 64704 26002 64708
rect 26018 64764 26082 64768
rect 26018 64708 26022 64764
rect 26022 64708 26078 64764
rect 26078 64708 26082 64764
rect 26018 64704 26082 64708
rect 10882 64220 10946 64224
rect 10882 64164 10886 64220
rect 10886 64164 10942 64220
rect 10942 64164 10946 64220
rect 10882 64160 10946 64164
rect 10962 64220 11026 64224
rect 10962 64164 10966 64220
rect 10966 64164 11022 64220
rect 11022 64164 11026 64220
rect 10962 64160 11026 64164
rect 11042 64220 11106 64224
rect 11042 64164 11046 64220
rect 11046 64164 11102 64220
rect 11102 64164 11106 64220
rect 11042 64160 11106 64164
rect 11122 64220 11186 64224
rect 11122 64164 11126 64220
rect 11126 64164 11182 64220
rect 11182 64164 11186 64220
rect 11122 64160 11186 64164
rect 20813 64220 20877 64224
rect 20813 64164 20817 64220
rect 20817 64164 20873 64220
rect 20873 64164 20877 64220
rect 20813 64160 20877 64164
rect 20893 64220 20957 64224
rect 20893 64164 20897 64220
rect 20897 64164 20953 64220
rect 20953 64164 20957 64220
rect 20893 64160 20957 64164
rect 20973 64220 21037 64224
rect 20973 64164 20977 64220
rect 20977 64164 21033 64220
rect 21033 64164 21037 64220
rect 20973 64160 21037 64164
rect 21053 64220 21117 64224
rect 21053 64164 21057 64220
rect 21057 64164 21113 64220
rect 21113 64164 21117 64220
rect 21053 64160 21117 64164
rect 27844 64092 27908 64156
rect 28212 64016 28276 64020
rect 28212 63960 28262 64016
rect 28262 63960 28276 64016
rect 28212 63956 28276 63960
rect 26556 63684 26620 63748
rect 5917 63676 5981 63680
rect 5917 63620 5921 63676
rect 5921 63620 5977 63676
rect 5977 63620 5981 63676
rect 5917 63616 5981 63620
rect 5997 63676 6061 63680
rect 5997 63620 6001 63676
rect 6001 63620 6057 63676
rect 6057 63620 6061 63676
rect 5997 63616 6061 63620
rect 6077 63676 6141 63680
rect 6077 63620 6081 63676
rect 6081 63620 6137 63676
rect 6137 63620 6141 63676
rect 6077 63616 6141 63620
rect 6157 63676 6221 63680
rect 6157 63620 6161 63676
rect 6161 63620 6217 63676
rect 6217 63620 6221 63676
rect 6157 63616 6221 63620
rect 15848 63676 15912 63680
rect 15848 63620 15852 63676
rect 15852 63620 15908 63676
rect 15908 63620 15912 63676
rect 15848 63616 15912 63620
rect 15928 63676 15992 63680
rect 15928 63620 15932 63676
rect 15932 63620 15988 63676
rect 15988 63620 15992 63676
rect 15928 63616 15992 63620
rect 16008 63676 16072 63680
rect 16008 63620 16012 63676
rect 16012 63620 16068 63676
rect 16068 63620 16072 63676
rect 16008 63616 16072 63620
rect 16088 63676 16152 63680
rect 16088 63620 16092 63676
rect 16092 63620 16148 63676
rect 16148 63620 16152 63676
rect 16088 63616 16152 63620
rect 25778 63676 25842 63680
rect 25778 63620 25782 63676
rect 25782 63620 25838 63676
rect 25838 63620 25842 63676
rect 25778 63616 25842 63620
rect 25858 63676 25922 63680
rect 25858 63620 25862 63676
rect 25862 63620 25918 63676
rect 25918 63620 25922 63676
rect 25858 63616 25922 63620
rect 25938 63676 26002 63680
rect 25938 63620 25942 63676
rect 25942 63620 25998 63676
rect 25998 63620 26002 63676
rect 25938 63616 26002 63620
rect 26018 63676 26082 63680
rect 26018 63620 26022 63676
rect 26022 63620 26078 63676
rect 26078 63620 26082 63676
rect 26018 63616 26082 63620
rect 28948 63412 29012 63476
rect 10882 63132 10946 63136
rect 10882 63076 10886 63132
rect 10886 63076 10942 63132
rect 10942 63076 10946 63132
rect 10882 63072 10946 63076
rect 10962 63132 11026 63136
rect 10962 63076 10966 63132
rect 10966 63076 11022 63132
rect 11022 63076 11026 63132
rect 10962 63072 11026 63076
rect 11042 63132 11106 63136
rect 11042 63076 11046 63132
rect 11046 63076 11102 63132
rect 11102 63076 11106 63132
rect 11042 63072 11106 63076
rect 11122 63132 11186 63136
rect 11122 63076 11126 63132
rect 11126 63076 11182 63132
rect 11182 63076 11186 63132
rect 11122 63072 11186 63076
rect 20813 63132 20877 63136
rect 20813 63076 20817 63132
rect 20817 63076 20873 63132
rect 20873 63076 20877 63132
rect 20813 63072 20877 63076
rect 20893 63132 20957 63136
rect 20893 63076 20897 63132
rect 20897 63076 20953 63132
rect 20953 63076 20957 63132
rect 20893 63072 20957 63076
rect 20973 63132 21037 63136
rect 20973 63076 20977 63132
rect 20977 63076 21033 63132
rect 21033 63076 21037 63132
rect 20973 63072 21037 63076
rect 21053 63132 21117 63136
rect 21053 63076 21057 63132
rect 21057 63076 21113 63132
rect 21113 63076 21117 63132
rect 21053 63072 21117 63076
rect 28396 63064 28460 63068
rect 28396 63008 28410 63064
rect 28410 63008 28460 63064
rect 27476 62928 27540 62932
rect 27476 62872 27526 62928
rect 27526 62872 27540 62928
rect 27476 62868 27540 62872
rect 28396 63004 28460 63008
rect 28580 63064 28644 63068
rect 28580 63008 28594 63064
rect 28594 63008 28644 63064
rect 28580 63004 28644 63008
rect 5917 62588 5981 62592
rect 5917 62532 5921 62588
rect 5921 62532 5977 62588
rect 5977 62532 5981 62588
rect 5917 62528 5981 62532
rect 5997 62588 6061 62592
rect 5997 62532 6001 62588
rect 6001 62532 6057 62588
rect 6057 62532 6061 62588
rect 5997 62528 6061 62532
rect 6077 62588 6141 62592
rect 6077 62532 6081 62588
rect 6081 62532 6137 62588
rect 6137 62532 6141 62588
rect 6077 62528 6141 62532
rect 6157 62588 6221 62592
rect 6157 62532 6161 62588
rect 6161 62532 6217 62588
rect 6217 62532 6221 62588
rect 6157 62528 6221 62532
rect 15848 62588 15912 62592
rect 15848 62532 15852 62588
rect 15852 62532 15908 62588
rect 15908 62532 15912 62588
rect 15848 62528 15912 62532
rect 15928 62588 15992 62592
rect 15928 62532 15932 62588
rect 15932 62532 15988 62588
rect 15988 62532 15992 62588
rect 15928 62528 15992 62532
rect 16008 62588 16072 62592
rect 16008 62532 16012 62588
rect 16012 62532 16068 62588
rect 16068 62532 16072 62588
rect 16008 62528 16072 62532
rect 16088 62588 16152 62592
rect 16088 62532 16092 62588
rect 16092 62532 16148 62588
rect 16148 62532 16152 62588
rect 16088 62528 16152 62532
rect 25778 62588 25842 62592
rect 25778 62532 25782 62588
rect 25782 62532 25838 62588
rect 25838 62532 25842 62588
rect 25778 62528 25842 62532
rect 25858 62588 25922 62592
rect 25858 62532 25862 62588
rect 25862 62532 25918 62588
rect 25918 62532 25922 62588
rect 25858 62528 25922 62532
rect 25938 62588 26002 62592
rect 25938 62532 25942 62588
rect 25942 62532 25998 62588
rect 25998 62532 26002 62588
rect 25938 62528 26002 62532
rect 26018 62588 26082 62592
rect 26018 62532 26022 62588
rect 26022 62532 26078 62588
rect 26078 62532 26082 62588
rect 26018 62528 26082 62532
rect 25268 62384 25332 62388
rect 25268 62328 25282 62384
rect 25282 62328 25332 62384
rect 25268 62324 25332 62328
rect 26188 62324 26252 62388
rect 28396 62052 28460 62116
rect 10882 62044 10946 62048
rect 10882 61988 10886 62044
rect 10886 61988 10942 62044
rect 10942 61988 10946 62044
rect 10882 61984 10946 61988
rect 10962 62044 11026 62048
rect 10962 61988 10966 62044
rect 10966 61988 11022 62044
rect 11022 61988 11026 62044
rect 10962 61984 11026 61988
rect 11042 62044 11106 62048
rect 11042 61988 11046 62044
rect 11046 61988 11102 62044
rect 11102 61988 11106 62044
rect 11042 61984 11106 61988
rect 11122 62044 11186 62048
rect 11122 61988 11126 62044
rect 11126 61988 11182 62044
rect 11182 61988 11186 62044
rect 11122 61984 11186 61988
rect 20813 62044 20877 62048
rect 20813 61988 20817 62044
rect 20817 61988 20873 62044
rect 20873 61988 20877 62044
rect 20813 61984 20877 61988
rect 20893 62044 20957 62048
rect 20893 61988 20897 62044
rect 20897 61988 20953 62044
rect 20953 61988 20957 62044
rect 20893 61984 20957 61988
rect 20973 62044 21037 62048
rect 20973 61988 20977 62044
rect 20977 61988 21033 62044
rect 21033 61988 21037 62044
rect 20973 61984 21037 61988
rect 21053 62044 21117 62048
rect 21053 61988 21057 62044
rect 21057 61988 21113 62044
rect 21113 61988 21117 62044
rect 21053 61984 21117 61988
rect 28580 61704 28644 61708
rect 28580 61648 28630 61704
rect 28630 61648 28644 61704
rect 28580 61644 28644 61648
rect 28764 61568 28828 61572
rect 28764 61512 28778 61568
rect 28778 61512 28828 61568
rect 28764 61508 28828 61512
rect 5917 61500 5981 61504
rect 5917 61444 5921 61500
rect 5921 61444 5977 61500
rect 5977 61444 5981 61500
rect 5917 61440 5981 61444
rect 5997 61500 6061 61504
rect 5997 61444 6001 61500
rect 6001 61444 6057 61500
rect 6057 61444 6061 61500
rect 5997 61440 6061 61444
rect 6077 61500 6141 61504
rect 6077 61444 6081 61500
rect 6081 61444 6137 61500
rect 6137 61444 6141 61500
rect 6077 61440 6141 61444
rect 6157 61500 6221 61504
rect 6157 61444 6161 61500
rect 6161 61444 6217 61500
rect 6217 61444 6221 61500
rect 6157 61440 6221 61444
rect 15848 61500 15912 61504
rect 15848 61444 15852 61500
rect 15852 61444 15908 61500
rect 15908 61444 15912 61500
rect 15848 61440 15912 61444
rect 15928 61500 15992 61504
rect 15928 61444 15932 61500
rect 15932 61444 15988 61500
rect 15988 61444 15992 61500
rect 15928 61440 15992 61444
rect 16008 61500 16072 61504
rect 16008 61444 16012 61500
rect 16012 61444 16068 61500
rect 16068 61444 16072 61500
rect 16008 61440 16072 61444
rect 16088 61500 16152 61504
rect 16088 61444 16092 61500
rect 16092 61444 16148 61500
rect 16148 61444 16152 61500
rect 16088 61440 16152 61444
rect 25778 61500 25842 61504
rect 25778 61444 25782 61500
rect 25782 61444 25838 61500
rect 25838 61444 25842 61500
rect 25778 61440 25842 61444
rect 25858 61500 25922 61504
rect 25858 61444 25862 61500
rect 25862 61444 25918 61500
rect 25918 61444 25922 61500
rect 25858 61440 25922 61444
rect 25938 61500 26002 61504
rect 25938 61444 25942 61500
rect 25942 61444 25998 61500
rect 25998 61444 26002 61500
rect 25938 61440 26002 61444
rect 26018 61500 26082 61504
rect 26018 61444 26022 61500
rect 26022 61444 26078 61500
rect 26078 61444 26082 61500
rect 26018 61440 26082 61444
rect 26924 61372 26988 61436
rect 29316 61372 29380 61436
rect 26740 61236 26804 61300
rect 28580 61236 28644 61300
rect 29132 61236 29196 61300
rect 28212 61100 28276 61164
rect 29500 61100 29564 61164
rect 26556 60964 26620 61028
rect 28212 60964 28276 61028
rect 10882 60956 10946 60960
rect 10882 60900 10886 60956
rect 10886 60900 10942 60956
rect 10942 60900 10946 60956
rect 10882 60896 10946 60900
rect 10962 60956 11026 60960
rect 10962 60900 10966 60956
rect 10966 60900 11022 60956
rect 11022 60900 11026 60956
rect 10962 60896 11026 60900
rect 11042 60956 11106 60960
rect 11042 60900 11046 60956
rect 11046 60900 11102 60956
rect 11102 60900 11106 60956
rect 11042 60896 11106 60900
rect 11122 60956 11186 60960
rect 11122 60900 11126 60956
rect 11126 60900 11182 60956
rect 11182 60900 11186 60956
rect 11122 60896 11186 60900
rect 20813 60956 20877 60960
rect 20813 60900 20817 60956
rect 20817 60900 20873 60956
rect 20873 60900 20877 60956
rect 20813 60896 20877 60900
rect 20893 60956 20957 60960
rect 20893 60900 20897 60956
rect 20897 60900 20953 60956
rect 20953 60900 20957 60956
rect 20893 60896 20957 60900
rect 20973 60956 21037 60960
rect 20973 60900 20977 60956
rect 20977 60900 21033 60956
rect 21033 60900 21037 60956
rect 20973 60896 21037 60900
rect 21053 60956 21117 60960
rect 21053 60900 21057 60956
rect 21057 60900 21113 60956
rect 21113 60900 21117 60956
rect 21053 60896 21117 60900
rect 25268 60888 25332 60892
rect 25268 60832 25318 60888
rect 25318 60832 25332 60888
rect 25268 60828 25332 60832
rect 26372 60828 26436 60892
rect 5917 60412 5981 60416
rect 5917 60356 5921 60412
rect 5921 60356 5977 60412
rect 5977 60356 5981 60412
rect 5917 60352 5981 60356
rect 5997 60412 6061 60416
rect 5997 60356 6001 60412
rect 6001 60356 6057 60412
rect 6057 60356 6061 60412
rect 5997 60352 6061 60356
rect 6077 60412 6141 60416
rect 6077 60356 6081 60412
rect 6081 60356 6137 60412
rect 6137 60356 6141 60412
rect 6077 60352 6141 60356
rect 6157 60412 6221 60416
rect 6157 60356 6161 60412
rect 6161 60356 6217 60412
rect 6217 60356 6221 60412
rect 6157 60352 6221 60356
rect 15848 60412 15912 60416
rect 15848 60356 15852 60412
rect 15852 60356 15908 60412
rect 15908 60356 15912 60412
rect 15848 60352 15912 60356
rect 15928 60412 15992 60416
rect 15928 60356 15932 60412
rect 15932 60356 15988 60412
rect 15988 60356 15992 60412
rect 15928 60352 15992 60356
rect 16008 60412 16072 60416
rect 16008 60356 16012 60412
rect 16012 60356 16068 60412
rect 16068 60356 16072 60412
rect 16008 60352 16072 60356
rect 16088 60412 16152 60416
rect 16088 60356 16092 60412
rect 16092 60356 16148 60412
rect 16148 60356 16152 60412
rect 16088 60352 16152 60356
rect 27292 60556 27356 60620
rect 26740 60420 26804 60484
rect 25778 60412 25842 60416
rect 25778 60356 25782 60412
rect 25782 60356 25838 60412
rect 25838 60356 25842 60412
rect 25778 60352 25842 60356
rect 25858 60412 25922 60416
rect 25858 60356 25862 60412
rect 25862 60356 25918 60412
rect 25918 60356 25922 60412
rect 25858 60352 25922 60356
rect 25938 60412 26002 60416
rect 25938 60356 25942 60412
rect 25942 60356 25998 60412
rect 25998 60356 26002 60412
rect 25938 60352 26002 60356
rect 26018 60412 26082 60416
rect 26018 60356 26022 60412
rect 26022 60356 26078 60412
rect 26078 60356 26082 60412
rect 26018 60352 26082 60356
rect 26924 60284 26988 60348
rect 29316 60480 29380 60484
rect 29316 60424 29366 60480
rect 29366 60424 29380 60480
rect 29316 60420 29380 60424
rect 28028 60284 28092 60348
rect 26188 60208 26252 60212
rect 26188 60152 26202 60208
rect 26202 60152 26252 60208
rect 26188 60148 26252 60152
rect 27844 60148 27908 60212
rect 28580 60148 28644 60212
rect 28212 60012 28276 60076
rect 28948 60012 29012 60076
rect 25268 59876 25332 59940
rect 10882 59868 10946 59872
rect 10882 59812 10886 59868
rect 10886 59812 10942 59868
rect 10942 59812 10946 59868
rect 10882 59808 10946 59812
rect 10962 59868 11026 59872
rect 10962 59812 10966 59868
rect 10966 59812 11022 59868
rect 11022 59812 11026 59868
rect 10962 59808 11026 59812
rect 11042 59868 11106 59872
rect 11042 59812 11046 59868
rect 11046 59812 11102 59868
rect 11102 59812 11106 59868
rect 11042 59808 11106 59812
rect 11122 59868 11186 59872
rect 11122 59812 11126 59868
rect 11126 59812 11182 59868
rect 11182 59812 11186 59868
rect 11122 59808 11186 59812
rect 20813 59868 20877 59872
rect 20813 59812 20817 59868
rect 20817 59812 20873 59868
rect 20873 59812 20877 59868
rect 20813 59808 20877 59812
rect 20893 59868 20957 59872
rect 20893 59812 20897 59868
rect 20897 59812 20953 59868
rect 20953 59812 20957 59868
rect 20893 59808 20957 59812
rect 20973 59868 21037 59872
rect 20973 59812 20977 59868
rect 20977 59812 21033 59868
rect 21033 59812 21037 59868
rect 20973 59808 21037 59812
rect 21053 59868 21117 59872
rect 21053 59812 21057 59868
rect 21057 59812 21113 59868
rect 21113 59812 21117 59868
rect 21053 59808 21117 59812
rect 27660 59740 27724 59804
rect 29684 59740 29748 59804
rect 25636 59604 25700 59668
rect 26556 59468 26620 59532
rect 28396 59468 28460 59532
rect 5917 59324 5981 59328
rect 5917 59268 5921 59324
rect 5921 59268 5977 59324
rect 5977 59268 5981 59324
rect 5917 59264 5981 59268
rect 5997 59324 6061 59328
rect 5997 59268 6001 59324
rect 6001 59268 6057 59324
rect 6057 59268 6061 59324
rect 5997 59264 6061 59268
rect 6077 59324 6141 59328
rect 6077 59268 6081 59324
rect 6081 59268 6137 59324
rect 6137 59268 6141 59324
rect 6077 59264 6141 59268
rect 6157 59324 6221 59328
rect 6157 59268 6161 59324
rect 6161 59268 6217 59324
rect 6217 59268 6221 59324
rect 6157 59264 6221 59268
rect 15848 59324 15912 59328
rect 15848 59268 15852 59324
rect 15852 59268 15908 59324
rect 15908 59268 15912 59324
rect 15848 59264 15912 59268
rect 15928 59324 15992 59328
rect 15928 59268 15932 59324
rect 15932 59268 15988 59324
rect 15988 59268 15992 59324
rect 15928 59264 15992 59268
rect 16008 59324 16072 59328
rect 16008 59268 16012 59324
rect 16012 59268 16068 59324
rect 16068 59268 16072 59324
rect 16008 59264 16072 59268
rect 16088 59324 16152 59328
rect 16088 59268 16092 59324
rect 16092 59268 16148 59324
rect 16148 59268 16152 59324
rect 16088 59264 16152 59268
rect 25778 59324 25842 59328
rect 25778 59268 25782 59324
rect 25782 59268 25838 59324
rect 25838 59268 25842 59324
rect 25778 59264 25842 59268
rect 25858 59324 25922 59328
rect 25858 59268 25862 59324
rect 25862 59268 25918 59324
rect 25918 59268 25922 59324
rect 25858 59264 25922 59268
rect 25938 59324 26002 59328
rect 25938 59268 25942 59324
rect 25942 59268 25998 59324
rect 25998 59268 26002 59324
rect 25938 59264 26002 59268
rect 26018 59324 26082 59328
rect 26018 59268 26022 59324
rect 26022 59268 26078 59324
rect 26078 59268 26082 59324
rect 26018 59264 26082 59268
rect 27108 59196 27172 59260
rect 28764 58788 28828 58852
rect 10882 58780 10946 58784
rect 10882 58724 10886 58780
rect 10886 58724 10942 58780
rect 10942 58724 10946 58780
rect 10882 58720 10946 58724
rect 10962 58780 11026 58784
rect 10962 58724 10966 58780
rect 10966 58724 11022 58780
rect 11022 58724 11026 58780
rect 10962 58720 11026 58724
rect 11042 58780 11106 58784
rect 11042 58724 11046 58780
rect 11046 58724 11102 58780
rect 11102 58724 11106 58780
rect 11042 58720 11106 58724
rect 11122 58780 11186 58784
rect 11122 58724 11126 58780
rect 11126 58724 11182 58780
rect 11182 58724 11186 58780
rect 11122 58720 11186 58724
rect 20813 58780 20877 58784
rect 20813 58724 20817 58780
rect 20817 58724 20873 58780
rect 20873 58724 20877 58780
rect 20813 58720 20877 58724
rect 20893 58780 20957 58784
rect 20893 58724 20897 58780
rect 20897 58724 20953 58780
rect 20953 58724 20957 58780
rect 20893 58720 20957 58724
rect 20973 58780 21037 58784
rect 20973 58724 20977 58780
rect 20977 58724 21033 58780
rect 21033 58724 21037 58780
rect 20973 58720 21037 58724
rect 21053 58780 21117 58784
rect 21053 58724 21057 58780
rect 21057 58724 21113 58780
rect 21113 58724 21117 58780
rect 21053 58720 21117 58724
rect 28764 58652 28828 58716
rect 27844 58516 27908 58580
rect 5917 58236 5981 58240
rect 5917 58180 5921 58236
rect 5921 58180 5977 58236
rect 5977 58180 5981 58236
rect 5917 58176 5981 58180
rect 5997 58236 6061 58240
rect 5997 58180 6001 58236
rect 6001 58180 6057 58236
rect 6057 58180 6061 58236
rect 5997 58176 6061 58180
rect 6077 58236 6141 58240
rect 6077 58180 6081 58236
rect 6081 58180 6137 58236
rect 6137 58180 6141 58236
rect 6077 58176 6141 58180
rect 6157 58236 6221 58240
rect 6157 58180 6161 58236
rect 6161 58180 6217 58236
rect 6217 58180 6221 58236
rect 6157 58176 6221 58180
rect 15848 58236 15912 58240
rect 15848 58180 15852 58236
rect 15852 58180 15908 58236
rect 15908 58180 15912 58236
rect 15848 58176 15912 58180
rect 15928 58236 15992 58240
rect 15928 58180 15932 58236
rect 15932 58180 15988 58236
rect 15988 58180 15992 58236
rect 15928 58176 15992 58180
rect 16008 58236 16072 58240
rect 16008 58180 16012 58236
rect 16012 58180 16068 58236
rect 16068 58180 16072 58236
rect 16008 58176 16072 58180
rect 16088 58236 16152 58240
rect 16088 58180 16092 58236
rect 16092 58180 16148 58236
rect 16148 58180 16152 58236
rect 16088 58176 16152 58180
rect 25778 58236 25842 58240
rect 25778 58180 25782 58236
rect 25782 58180 25838 58236
rect 25838 58180 25842 58236
rect 25778 58176 25842 58180
rect 25858 58236 25922 58240
rect 25858 58180 25862 58236
rect 25862 58180 25918 58236
rect 25918 58180 25922 58236
rect 25858 58176 25922 58180
rect 25938 58236 26002 58240
rect 25938 58180 25942 58236
rect 25942 58180 25998 58236
rect 25998 58180 26002 58236
rect 25938 58176 26002 58180
rect 26018 58236 26082 58240
rect 26018 58180 26022 58236
rect 26022 58180 26078 58236
rect 26078 58180 26082 58236
rect 26018 58176 26082 58180
rect 27476 57836 27540 57900
rect 29868 57836 29932 57900
rect 27476 57760 27540 57764
rect 27476 57704 27490 57760
rect 27490 57704 27540 57760
rect 27476 57700 27540 57704
rect 10882 57692 10946 57696
rect 10882 57636 10886 57692
rect 10886 57636 10942 57692
rect 10942 57636 10946 57692
rect 10882 57632 10946 57636
rect 10962 57692 11026 57696
rect 10962 57636 10966 57692
rect 10966 57636 11022 57692
rect 11022 57636 11026 57692
rect 10962 57632 11026 57636
rect 11042 57692 11106 57696
rect 11042 57636 11046 57692
rect 11046 57636 11102 57692
rect 11102 57636 11106 57692
rect 11042 57632 11106 57636
rect 11122 57692 11186 57696
rect 11122 57636 11126 57692
rect 11126 57636 11182 57692
rect 11182 57636 11186 57692
rect 11122 57632 11186 57636
rect 20813 57692 20877 57696
rect 20813 57636 20817 57692
rect 20817 57636 20873 57692
rect 20873 57636 20877 57692
rect 20813 57632 20877 57636
rect 20893 57692 20957 57696
rect 20893 57636 20897 57692
rect 20897 57636 20953 57692
rect 20953 57636 20957 57692
rect 20893 57632 20957 57636
rect 20973 57692 21037 57696
rect 20973 57636 20977 57692
rect 20977 57636 21033 57692
rect 21033 57636 21037 57692
rect 20973 57632 21037 57636
rect 21053 57692 21117 57696
rect 21053 57636 21057 57692
rect 21057 57636 21113 57692
rect 21113 57636 21117 57692
rect 21053 57632 21117 57636
rect 26188 57564 26252 57628
rect 26924 57564 26988 57628
rect 23980 57292 24044 57356
rect 26372 57292 26436 57356
rect 27660 57156 27724 57220
rect 30052 57156 30116 57220
rect 30604 57216 30668 57220
rect 30604 57160 30654 57216
rect 30654 57160 30668 57216
rect 30604 57156 30668 57160
rect 5917 57148 5981 57152
rect 5917 57092 5921 57148
rect 5921 57092 5977 57148
rect 5977 57092 5981 57148
rect 5917 57088 5981 57092
rect 5997 57148 6061 57152
rect 5997 57092 6001 57148
rect 6001 57092 6057 57148
rect 6057 57092 6061 57148
rect 5997 57088 6061 57092
rect 6077 57148 6141 57152
rect 6077 57092 6081 57148
rect 6081 57092 6137 57148
rect 6137 57092 6141 57148
rect 6077 57088 6141 57092
rect 6157 57148 6221 57152
rect 6157 57092 6161 57148
rect 6161 57092 6217 57148
rect 6217 57092 6221 57148
rect 6157 57088 6221 57092
rect 15848 57148 15912 57152
rect 15848 57092 15852 57148
rect 15852 57092 15908 57148
rect 15908 57092 15912 57148
rect 15848 57088 15912 57092
rect 15928 57148 15992 57152
rect 15928 57092 15932 57148
rect 15932 57092 15988 57148
rect 15988 57092 15992 57148
rect 15928 57088 15992 57092
rect 16008 57148 16072 57152
rect 16008 57092 16012 57148
rect 16012 57092 16068 57148
rect 16068 57092 16072 57148
rect 16008 57088 16072 57092
rect 16088 57148 16152 57152
rect 16088 57092 16092 57148
rect 16092 57092 16148 57148
rect 16148 57092 16152 57148
rect 16088 57088 16152 57092
rect 25778 57148 25842 57152
rect 25778 57092 25782 57148
rect 25782 57092 25838 57148
rect 25838 57092 25842 57148
rect 25778 57088 25842 57092
rect 25858 57148 25922 57152
rect 25858 57092 25862 57148
rect 25862 57092 25918 57148
rect 25918 57092 25922 57148
rect 25858 57088 25922 57092
rect 25938 57148 26002 57152
rect 25938 57092 25942 57148
rect 25942 57092 25998 57148
rect 25998 57092 26002 57148
rect 25938 57088 26002 57092
rect 26018 57148 26082 57152
rect 26018 57092 26022 57148
rect 26022 57092 26078 57148
rect 26078 57092 26082 57148
rect 26018 57088 26082 57092
rect 23428 56884 23492 56948
rect 29500 56884 29564 56948
rect 17356 56748 17420 56812
rect 29132 56748 29196 56812
rect 23612 56672 23676 56676
rect 23612 56616 23626 56672
rect 23626 56616 23676 56672
rect 23612 56612 23676 56616
rect 25084 56612 25148 56676
rect 10882 56604 10946 56608
rect 10882 56548 10886 56604
rect 10886 56548 10942 56604
rect 10942 56548 10946 56604
rect 10882 56544 10946 56548
rect 10962 56604 11026 56608
rect 10962 56548 10966 56604
rect 10966 56548 11022 56604
rect 11022 56548 11026 56604
rect 10962 56544 11026 56548
rect 11042 56604 11106 56608
rect 11042 56548 11046 56604
rect 11046 56548 11102 56604
rect 11102 56548 11106 56604
rect 11042 56544 11106 56548
rect 11122 56604 11186 56608
rect 11122 56548 11126 56604
rect 11126 56548 11182 56604
rect 11182 56548 11186 56604
rect 11122 56544 11186 56548
rect 20813 56604 20877 56608
rect 20813 56548 20817 56604
rect 20817 56548 20873 56604
rect 20873 56548 20877 56604
rect 20813 56544 20877 56548
rect 20893 56604 20957 56608
rect 20893 56548 20897 56604
rect 20897 56548 20953 56604
rect 20953 56548 20957 56604
rect 20893 56544 20957 56548
rect 20973 56604 21037 56608
rect 20973 56548 20977 56604
rect 20977 56548 21033 56604
rect 21033 56548 21037 56604
rect 20973 56544 21037 56548
rect 21053 56604 21117 56608
rect 21053 56548 21057 56604
rect 21057 56548 21113 56604
rect 21113 56548 21117 56604
rect 21053 56544 21117 56548
rect 5917 56060 5981 56064
rect 5917 56004 5921 56060
rect 5921 56004 5977 56060
rect 5977 56004 5981 56060
rect 5917 56000 5981 56004
rect 5997 56060 6061 56064
rect 5997 56004 6001 56060
rect 6001 56004 6057 56060
rect 6057 56004 6061 56060
rect 5997 56000 6061 56004
rect 6077 56060 6141 56064
rect 6077 56004 6081 56060
rect 6081 56004 6137 56060
rect 6137 56004 6141 56060
rect 6077 56000 6141 56004
rect 6157 56060 6221 56064
rect 6157 56004 6161 56060
rect 6161 56004 6217 56060
rect 6217 56004 6221 56060
rect 6157 56000 6221 56004
rect 15848 56060 15912 56064
rect 15848 56004 15852 56060
rect 15852 56004 15908 56060
rect 15908 56004 15912 56060
rect 15848 56000 15912 56004
rect 15928 56060 15992 56064
rect 15928 56004 15932 56060
rect 15932 56004 15988 56060
rect 15988 56004 15992 56060
rect 15928 56000 15992 56004
rect 16008 56060 16072 56064
rect 16008 56004 16012 56060
rect 16012 56004 16068 56060
rect 16068 56004 16072 56060
rect 16008 56000 16072 56004
rect 16088 56060 16152 56064
rect 16088 56004 16092 56060
rect 16092 56004 16148 56060
rect 16148 56004 16152 56060
rect 16088 56000 16152 56004
rect 25778 56060 25842 56064
rect 25778 56004 25782 56060
rect 25782 56004 25838 56060
rect 25838 56004 25842 56060
rect 25778 56000 25842 56004
rect 25858 56060 25922 56064
rect 25858 56004 25862 56060
rect 25862 56004 25918 56060
rect 25918 56004 25922 56060
rect 25858 56000 25922 56004
rect 25938 56060 26002 56064
rect 25938 56004 25942 56060
rect 25942 56004 25998 56060
rect 25998 56004 26002 56060
rect 25938 56000 26002 56004
rect 26018 56060 26082 56064
rect 26018 56004 26022 56060
rect 26022 56004 26078 56060
rect 26078 56004 26082 56060
rect 26018 56000 26082 56004
rect 23796 55856 23860 55860
rect 23796 55800 23846 55856
rect 23846 55800 23860 55856
rect 23796 55796 23860 55800
rect 24900 55796 24964 55860
rect 30788 55660 30852 55724
rect 10882 55516 10946 55520
rect 10882 55460 10886 55516
rect 10886 55460 10942 55516
rect 10942 55460 10946 55516
rect 10882 55456 10946 55460
rect 10962 55516 11026 55520
rect 10962 55460 10966 55516
rect 10966 55460 11022 55516
rect 11022 55460 11026 55516
rect 10962 55456 11026 55460
rect 11042 55516 11106 55520
rect 11042 55460 11046 55516
rect 11046 55460 11102 55516
rect 11102 55460 11106 55516
rect 11042 55456 11106 55460
rect 11122 55516 11186 55520
rect 11122 55460 11126 55516
rect 11126 55460 11182 55516
rect 11182 55460 11186 55516
rect 11122 55456 11186 55460
rect 20813 55516 20877 55520
rect 20813 55460 20817 55516
rect 20817 55460 20873 55516
rect 20873 55460 20877 55516
rect 20813 55456 20877 55460
rect 20893 55516 20957 55520
rect 20893 55460 20897 55516
rect 20897 55460 20953 55516
rect 20953 55460 20957 55516
rect 20893 55456 20957 55460
rect 20973 55516 21037 55520
rect 20973 55460 20977 55516
rect 20977 55460 21033 55516
rect 21033 55460 21037 55516
rect 20973 55456 21037 55460
rect 21053 55516 21117 55520
rect 21053 55460 21057 55516
rect 21057 55460 21113 55516
rect 21113 55460 21117 55516
rect 21053 55456 21117 55460
rect 27292 55388 27356 55452
rect 25084 54980 25148 55044
rect 5917 54972 5981 54976
rect 5917 54916 5921 54972
rect 5921 54916 5977 54972
rect 5977 54916 5981 54972
rect 5917 54912 5981 54916
rect 5997 54972 6061 54976
rect 5997 54916 6001 54972
rect 6001 54916 6057 54972
rect 6057 54916 6061 54972
rect 5997 54912 6061 54916
rect 6077 54972 6141 54976
rect 6077 54916 6081 54972
rect 6081 54916 6137 54972
rect 6137 54916 6141 54972
rect 6077 54912 6141 54916
rect 6157 54972 6221 54976
rect 6157 54916 6161 54972
rect 6161 54916 6217 54972
rect 6217 54916 6221 54972
rect 6157 54912 6221 54916
rect 15848 54972 15912 54976
rect 15848 54916 15852 54972
rect 15852 54916 15908 54972
rect 15908 54916 15912 54972
rect 15848 54912 15912 54916
rect 15928 54972 15992 54976
rect 15928 54916 15932 54972
rect 15932 54916 15988 54972
rect 15988 54916 15992 54972
rect 15928 54912 15992 54916
rect 16008 54972 16072 54976
rect 16008 54916 16012 54972
rect 16012 54916 16068 54972
rect 16068 54916 16072 54972
rect 16008 54912 16072 54916
rect 16088 54972 16152 54976
rect 16088 54916 16092 54972
rect 16092 54916 16148 54972
rect 16148 54916 16152 54972
rect 16088 54912 16152 54916
rect 25778 54972 25842 54976
rect 25778 54916 25782 54972
rect 25782 54916 25838 54972
rect 25838 54916 25842 54972
rect 25778 54912 25842 54916
rect 25858 54972 25922 54976
rect 25858 54916 25862 54972
rect 25862 54916 25918 54972
rect 25918 54916 25922 54972
rect 25858 54912 25922 54916
rect 25938 54972 26002 54976
rect 25938 54916 25942 54972
rect 25942 54916 25998 54972
rect 25998 54916 26002 54972
rect 25938 54912 26002 54916
rect 26018 54972 26082 54976
rect 26018 54916 26022 54972
rect 26022 54916 26078 54972
rect 26078 54916 26082 54972
rect 26018 54912 26082 54916
rect 24532 54844 24596 54908
rect 24716 54844 24780 54908
rect 28212 55252 28276 55316
rect 27108 54708 27172 54772
rect 28580 54572 28644 54636
rect 30052 54980 30116 55044
rect 31524 54436 31588 54500
rect 10882 54428 10946 54432
rect 10882 54372 10886 54428
rect 10886 54372 10942 54428
rect 10942 54372 10946 54428
rect 10882 54368 10946 54372
rect 10962 54428 11026 54432
rect 10962 54372 10966 54428
rect 10966 54372 11022 54428
rect 11022 54372 11026 54428
rect 10962 54368 11026 54372
rect 11042 54428 11106 54432
rect 11042 54372 11046 54428
rect 11046 54372 11102 54428
rect 11102 54372 11106 54428
rect 11042 54368 11106 54372
rect 11122 54428 11186 54432
rect 11122 54372 11126 54428
rect 11126 54372 11182 54428
rect 11182 54372 11186 54428
rect 11122 54368 11186 54372
rect 20813 54428 20877 54432
rect 20813 54372 20817 54428
rect 20817 54372 20873 54428
rect 20873 54372 20877 54428
rect 20813 54368 20877 54372
rect 20893 54428 20957 54432
rect 20893 54372 20897 54428
rect 20897 54372 20953 54428
rect 20953 54372 20957 54428
rect 20893 54368 20957 54372
rect 20973 54428 21037 54432
rect 20973 54372 20977 54428
rect 20977 54372 21033 54428
rect 21033 54372 21037 54428
rect 20973 54368 21037 54372
rect 21053 54428 21117 54432
rect 21053 54372 21057 54428
rect 21057 54372 21113 54428
rect 21113 54372 21117 54428
rect 21053 54368 21117 54372
rect 26372 54300 26436 54364
rect 26372 54164 26436 54228
rect 25268 54088 25332 54092
rect 25268 54032 25282 54088
rect 25282 54032 25332 54088
rect 25268 54028 25332 54032
rect 28764 54028 28828 54092
rect 5917 53884 5981 53888
rect 5917 53828 5921 53884
rect 5921 53828 5977 53884
rect 5977 53828 5981 53884
rect 5917 53824 5981 53828
rect 5997 53884 6061 53888
rect 5997 53828 6001 53884
rect 6001 53828 6057 53884
rect 6057 53828 6061 53884
rect 5997 53824 6061 53828
rect 6077 53884 6141 53888
rect 6077 53828 6081 53884
rect 6081 53828 6137 53884
rect 6137 53828 6141 53884
rect 6077 53824 6141 53828
rect 6157 53884 6221 53888
rect 6157 53828 6161 53884
rect 6161 53828 6217 53884
rect 6217 53828 6221 53884
rect 6157 53824 6221 53828
rect 15848 53884 15912 53888
rect 15848 53828 15852 53884
rect 15852 53828 15908 53884
rect 15908 53828 15912 53884
rect 15848 53824 15912 53828
rect 15928 53884 15992 53888
rect 15928 53828 15932 53884
rect 15932 53828 15988 53884
rect 15988 53828 15992 53884
rect 15928 53824 15992 53828
rect 16008 53884 16072 53888
rect 16008 53828 16012 53884
rect 16012 53828 16068 53884
rect 16068 53828 16072 53884
rect 16008 53824 16072 53828
rect 16088 53884 16152 53888
rect 16088 53828 16092 53884
rect 16092 53828 16148 53884
rect 16148 53828 16152 53884
rect 16088 53824 16152 53828
rect 25778 53884 25842 53888
rect 25778 53828 25782 53884
rect 25782 53828 25838 53884
rect 25838 53828 25842 53884
rect 25778 53824 25842 53828
rect 25858 53884 25922 53888
rect 25858 53828 25862 53884
rect 25862 53828 25918 53884
rect 25918 53828 25922 53884
rect 25858 53824 25922 53828
rect 25938 53884 26002 53888
rect 25938 53828 25942 53884
rect 25942 53828 25998 53884
rect 25998 53828 26002 53884
rect 25938 53824 26002 53828
rect 26018 53884 26082 53888
rect 26018 53828 26022 53884
rect 26022 53828 26078 53884
rect 26078 53828 26082 53884
rect 26018 53824 26082 53828
rect 19196 53756 19260 53820
rect 23612 53756 23676 53820
rect 27844 53816 27908 53820
rect 27844 53760 27894 53816
rect 27894 53760 27908 53816
rect 27844 53756 27908 53760
rect 17540 53620 17604 53684
rect 29500 53620 29564 53684
rect 30236 53484 30300 53548
rect 28396 53348 28460 53412
rect 28948 53348 29012 53412
rect 10882 53340 10946 53344
rect 10882 53284 10886 53340
rect 10886 53284 10942 53340
rect 10942 53284 10946 53340
rect 10882 53280 10946 53284
rect 10962 53340 11026 53344
rect 10962 53284 10966 53340
rect 10966 53284 11022 53340
rect 11022 53284 11026 53340
rect 10962 53280 11026 53284
rect 11042 53340 11106 53344
rect 11042 53284 11046 53340
rect 11046 53284 11102 53340
rect 11102 53284 11106 53340
rect 11042 53280 11106 53284
rect 11122 53340 11186 53344
rect 11122 53284 11126 53340
rect 11126 53284 11182 53340
rect 11182 53284 11186 53340
rect 11122 53280 11186 53284
rect 20813 53340 20877 53344
rect 20813 53284 20817 53340
rect 20817 53284 20873 53340
rect 20873 53284 20877 53340
rect 20813 53280 20877 53284
rect 20893 53340 20957 53344
rect 20893 53284 20897 53340
rect 20897 53284 20953 53340
rect 20953 53284 20957 53340
rect 20893 53280 20957 53284
rect 20973 53340 21037 53344
rect 20973 53284 20977 53340
rect 20977 53284 21033 53340
rect 21033 53284 21037 53340
rect 20973 53280 21037 53284
rect 21053 53340 21117 53344
rect 21053 53284 21057 53340
rect 21057 53284 21113 53340
rect 21113 53284 21117 53340
rect 21053 53280 21117 53284
rect 28764 53076 28828 53140
rect 29316 53136 29380 53140
rect 29316 53080 29330 53136
rect 29330 53080 29380 53136
rect 29316 53076 29380 53080
rect 30788 53076 30852 53140
rect 24164 52940 24228 53004
rect 27108 52940 27172 53004
rect 28028 52940 28092 53004
rect 23244 52804 23308 52868
rect 5917 52796 5981 52800
rect 5917 52740 5921 52796
rect 5921 52740 5977 52796
rect 5977 52740 5981 52796
rect 5917 52736 5981 52740
rect 5997 52796 6061 52800
rect 5997 52740 6001 52796
rect 6001 52740 6057 52796
rect 6057 52740 6061 52796
rect 5997 52736 6061 52740
rect 6077 52796 6141 52800
rect 6077 52740 6081 52796
rect 6081 52740 6137 52796
rect 6137 52740 6141 52796
rect 6077 52736 6141 52740
rect 6157 52796 6221 52800
rect 6157 52740 6161 52796
rect 6161 52740 6217 52796
rect 6217 52740 6221 52796
rect 6157 52736 6221 52740
rect 15848 52796 15912 52800
rect 15848 52740 15852 52796
rect 15852 52740 15908 52796
rect 15908 52740 15912 52796
rect 15848 52736 15912 52740
rect 15928 52796 15992 52800
rect 15928 52740 15932 52796
rect 15932 52740 15988 52796
rect 15988 52740 15992 52796
rect 15928 52736 15992 52740
rect 16008 52796 16072 52800
rect 16008 52740 16012 52796
rect 16012 52740 16068 52796
rect 16068 52740 16072 52796
rect 16008 52736 16072 52740
rect 16088 52796 16152 52800
rect 16088 52740 16092 52796
rect 16092 52740 16148 52796
rect 16148 52740 16152 52796
rect 16088 52736 16152 52740
rect 25778 52796 25842 52800
rect 25778 52740 25782 52796
rect 25782 52740 25838 52796
rect 25838 52740 25842 52796
rect 25778 52736 25842 52740
rect 25858 52796 25922 52800
rect 25858 52740 25862 52796
rect 25862 52740 25918 52796
rect 25918 52740 25922 52796
rect 25858 52736 25922 52740
rect 25938 52796 26002 52800
rect 25938 52740 25942 52796
rect 25942 52740 25998 52796
rect 25998 52740 26002 52796
rect 25938 52736 26002 52740
rect 26018 52796 26082 52800
rect 26018 52740 26022 52796
rect 26022 52740 26078 52796
rect 26078 52740 26082 52796
rect 26018 52736 26082 52740
rect 28028 52728 28092 52732
rect 28028 52672 28042 52728
rect 28042 52672 28092 52728
rect 28028 52668 28092 52672
rect 28396 52668 28460 52732
rect 30420 52668 30484 52732
rect 29316 52592 29380 52596
rect 29316 52536 29366 52592
rect 29366 52536 29380 52592
rect 23612 52396 23676 52460
rect 26556 52260 26620 52324
rect 10882 52252 10946 52256
rect 10882 52196 10886 52252
rect 10886 52196 10942 52252
rect 10942 52196 10946 52252
rect 10882 52192 10946 52196
rect 10962 52252 11026 52256
rect 10962 52196 10966 52252
rect 10966 52196 11022 52252
rect 11022 52196 11026 52252
rect 10962 52192 11026 52196
rect 11042 52252 11106 52256
rect 11042 52196 11046 52252
rect 11046 52196 11102 52252
rect 11102 52196 11106 52252
rect 11042 52192 11106 52196
rect 11122 52252 11186 52256
rect 11122 52196 11126 52252
rect 11126 52196 11182 52252
rect 11182 52196 11186 52252
rect 11122 52192 11186 52196
rect 20813 52252 20877 52256
rect 20813 52196 20817 52252
rect 20817 52196 20873 52252
rect 20873 52196 20877 52252
rect 20813 52192 20877 52196
rect 20893 52252 20957 52256
rect 20893 52196 20897 52252
rect 20897 52196 20953 52252
rect 20953 52196 20957 52252
rect 20893 52192 20957 52196
rect 20973 52252 21037 52256
rect 20973 52196 20977 52252
rect 20977 52196 21033 52252
rect 21033 52196 21037 52252
rect 20973 52192 21037 52196
rect 21053 52252 21117 52256
rect 21053 52196 21057 52252
rect 21057 52196 21113 52252
rect 21113 52196 21117 52252
rect 21053 52192 21117 52196
rect 26556 52124 26620 52188
rect 27292 52124 27356 52188
rect 27292 51988 27356 52052
rect 27660 51988 27724 52052
rect 29316 52532 29380 52536
rect 28764 52396 28828 52460
rect 28948 52124 29012 52188
rect 30236 52124 30300 52188
rect 26924 51852 26988 51916
rect 27660 51852 27724 51916
rect 29868 51716 29932 51780
rect 5917 51708 5981 51712
rect 5917 51652 5921 51708
rect 5921 51652 5977 51708
rect 5977 51652 5981 51708
rect 5917 51648 5981 51652
rect 5997 51708 6061 51712
rect 5997 51652 6001 51708
rect 6001 51652 6057 51708
rect 6057 51652 6061 51708
rect 5997 51648 6061 51652
rect 6077 51708 6141 51712
rect 6077 51652 6081 51708
rect 6081 51652 6137 51708
rect 6137 51652 6141 51708
rect 6077 51648 6141 51652
rect 6157 51708 6221 51712
rect 6157 51652 6161 51708
rect 6161 51652 6217 51708
rect 6217 51652 6221 51708
rect 6157 51648 6221 51652
rect 15848 51708 15912 51712
rect 15848 51652 15852 51708
rect 15852 51652 15908 51708
rect 15908 51652 15912 51708
rect 15848 51648 15912 51652
rect 15928 51708 15992 51712
rect 15928 51652 15932 51708
rect 15932 51652 15988 51708
rect 15988 51652 15992 51708
rect 15928 51648 15992 51652
rect 16008 51708 16072 51712
rect 16008 51652 16012 51708
rect 16012 51652 16068 51708
rect 16068 51652 16072 51708
rect 16008 51648 16072 51652
rect 16088 51708 16152 51712
rect 16088 51652 16092 51708
rect 16092 51652 16148 51708
rect 16148 51652 16152 51708
rect 16088 51648 16152 51652
rect 25778 51708 25842 51712
rect 25778 51652 25782 51708
rect 25782 51652 25838 51708
rect 25838 51652 25842 51708
rect 25778 51648 25842 51652
rect 25858 51708 25922 51712
rect 25858 51652 25862 51708
rect 25862 51652 25918 51708
rect 25918 51652 25922 51708
rect 25858 51648 25922 51652
rect 25938 51708 26002 51712
rect 25938 51652 25942 51708
rect 25942 51652 25998 51708
rect 25998 51652 26002 51708
rect 25938 51648 26002 51652
rect 26018 51708 26082 51712
rect 26018 51652 26022 51708
rect 26022 51652 26078 51708
rect 26078 51652 26082 51708
rect 26018 51648 26082 51652
rect 24348 51580 24412 51644
rect 29868 51640 29932 51644
rect 29868 51584 29918 51640
rect 29918 51584 29932 51640
rect 29868 51580 29932 51584
rect 23980 51444 24044 51508
rect 23428 51368 23492 51372
rect 23428 51312 23478 51368
rect 23478 51312 23492 51368
rect 23428 51308 23492 51312
rect 23612 51308 23676 51372
rect 10882 51164 10946 51168
rect 10882 51108 10886 51164
rect 10886 51108 10942 51164
rect 10942 51108 10946 51164
rect 10882 51104 10946 51108
rect 10962 51164 11026 51168
rect 10962 51108 10966 51164
rect 10966 51108 11022 51164
rect 11022 51108 11026 51164
rect 10962 51104 11026 51108
rect 11042 51164 11106 51168
rect 11042 51108 11046 51164
rect 11046 51108 11102 51164
rect 11102 51108 11106 51164
rect 11042 51104 11106 51108
rect 11122 51164 11186 51168
rect 11122 51108 11126 51164
rect 11126 51108 11182 51164
rect 11182 51108 11186 51164
rect 11122 51104 11186 51108
rect 20813 51164 20877 51168
rect 20813 51108 20817 51164
rect 20817 51108 20873 51164
rect 20873 51108 20877 51164
rect 20813 51104 20877 51108
rect 20893 51164 20957 51168
rect 20893 51108 20897 51164
rect 20897 51108 20953 51164
rect 20953 51108 20957 51164
rect 20893 51104 20957 51108
rect 20973 51164 21037 51168
rect 20973 51108 20977 51164
rect 20977 51108 21033 51164
rect 21033 51108 21037 51164
rect 20973 51104 21037 51108
rect 21053 51164 21117 51168
rect 21053 51108 21057 51164
rect 21057 51108 21113 51164
rect 21113 51108 21117 51164
rect 21053 51104 21117 51108
rect 24532 51096 24596 51100
rect 25636 51172 25700 51236
rect 26372 51308 26436 51372
rect 27108 51308 27172 51372
rect 29316 51368 29380 51372
rect 29316 51312 29366 51368
rect 29366 51312 29380 51368
rect 29316 51308 29380 51312
rect 29684 51368 29748 51372
rect 29684 51312 29698 51368
rect 29698 51312 29748 51368
rect 29684 51308 29748 51312
rect 26372 51232 26436 51236
rect 26372 51176 26422 51232
rect 26422 51176 26436 51232
rect 26372 51172 26436 51176
rect 27844 51232 27908 51236
rect 27844 51176 27858 51232
rect 27858 51176 27908 51232
rect 27844 51172 27908 51176
rect 28396 51172 28460 51236
rect 30052 51172 30116 51236
rect 30788 51172 30852 51236
rect 31156 51172 31220 51236
rect 24532 51040 24546 51096
rect 24546 51040 24596 51096
rect 24532 51036 24596 51040
rect 29132 51096 29196 51100
rect 29132 51040 29146 51096
rect 29146 51040 29196 51096
rect 29132 51036 29196 51040
rect 21404 50900 21468 50964
rect 24164 50900 24228 50964
rect 24532 50900 24596 50964
rect 27660 50900 27724 50964
rect 30420 50960 30484 50964
rect 30420 50904 30470 50960
rect 30470 50904 30484 50960
rect 30420 50900 30484 50904
rect 30972 50960 31036 50964
rect 30972 50904 30986 50960
rect 30986 50904 31036 50960
rect 30972 50900 31036 50904
rect 17724 50764 17788 50828
rect 24716 50628 24780 50692
rect 29868 50688 29932 50692
rect 29868 50632 29882 50688
rect 29882 50632 29932 50688
rect 29868 50628 29932 50632
rect 30788 50628 30852 50692
rect 5917 50620 5981 50624
rect 5917 50564 5921 50620
rect 5921 50564 5977 50620
rect 5977 50564 5981 50620
rect 5917 50560 5981 50564
rect 5997 50620 6061 50624
rect 5997 50564 6001 50620
rect 6001 50564 6057 50620
rect 6057 50564 6061 50620
rect 5997 50560 6061 50564
rect 6077 50620 6141 50624
rect 6077 50564 6081 50620
rect 6081 50564 6137 50620
rect 6137 50564 6141 50620
rect 6077 50560 6141 50564
rect 6157 50620 6221 50624
rect 6157 50564 6161 50620
rect 6161 50564 6217 50620
rect 6217 50564 6221 50620
rect 6157 50560 6221 50564
rect 15848 50620 15912 50624
rect 15848 50564 15852 50620
rect 15852 50564 15908 50620
rect 15908 50564 15912 50620
rect 15848 50560 15912 50564
rect 15928 50620 15992 50624
rect 15928 50564 15932 50620
rect 15932 50564 15988 50620
rect 15988 50564 15992 50620
rect 15928 50560 15992 50564
rect 16008 50620 16072 50624
rect 16008 50564 16012 50620
rect 16012 50564 16068 50620
rect 16068 50564 16072 50620
rect 16008 50560 16072 50564
rect 16088 50620 16152 50624
rect 16088 50564 16092 50620
rect 16092 50564 16148 50620
rect 16148 50564 16152 50620
rect 16088 50560 16152 50564
rect 25778 50620 25842 50624
rect 25778 50564 25782 50620
rect 25782 50564 25838 50620
rect 25838 50564 25842 50620
rect 25778 50560 25842 50564
rect 25858 50620 25922 50624
rect 25858 50564 25862 50620
rect 25862 50564 25918 50620
rect 25918 50564 25922 50620
rect 25858 50560 25922 50564
rect 25938 50620 26002 50624
rect 25938 50564 25942 50620
rect 25942 50564 25998 50620
rect 25998 50564 26002 50620
rect 25938 50560 26002 50564
rect 26018 50620 26082 50624
rect 26018 50564 26022 50620
rect 26022 50564 26078 50620
rect 26078 50564 26082 50620
rect 26018 50560 26082 50564
rect 24532 50492 24596 50556
rect 23612 50356 23676 50420
rect 25452 50356 25516 50420
rect 30052 50356 30116 50420
rect 30604 50220 30668 50284
rect 10882 50076 10946 50080
rect 10882 50020 10886 50076
rect 10886 50020 10942 50076
rect 10942 50020 10946 50076
rect 10882 50016 10946 50020
rect 10962 50076 11026 50080
rect 10962 50020 10966 50076
rect 10966 50020 11022 50076
rect 11022 50020 11026 50076
rect 10962 50016 11026 50020
rect 11042 50076 11106 50080
rect 11042 50020 11046 50076
rect 11046 50020 11102 50076
rect 11102 50020 11106 50076
rect 11042 50016 11106 50020
rect 11122 50076 11186 50080
rect 11122 50020 11126 50076
rect 11126 50020 11182 50076
rect 11182 50020 11186 50076
rect 11122 50016 11186 50020
rect 20813 50076 20877 50080
rect 20813 50020 20817 50076
rect 20817 50020 20873 50076
rect 20873 50020 20877 50076
rect 20813 50016 20877 50020
rect 20893 50076 20957 50080
rect 20893 50020 20897 50076
rect 20897 50020 20953 50076
rect 20953 50020 20957 50076
rect 20893 50016 20957 50020
rect 20973 50076 21037 50080
rect 20973 50020 20977 50076
rect 20977 50020 21033 50076
rect 21033 50020 21037 50076
rect 20973 50016 21037 50020
rect 21053 50076 21117 50080
rect 21053 50020 21057 50076
rect 21057 50020 21113 50076
rect 21113 50020 21117 50076
rect 21053 50016 21117 50020
rect 27660 50084 27724 50148
rect 23796 49948 23860 50012
rect 23980 50008 24044 50012
rect 23980 49952 23994 50008
rect 23994 49952 24044 50008
rect 23980 49948 24044 49952
rect 24716 50008 24780 50012
rect 24716 49952 24766 50008
rect 24766 49952 24780 50008
rect 24716 49948 24780 49952
rect 26924 49948 26988 50012
rect 23244 49812 23308 49876
rect 24348 49676 24412 49740
rect 5917 49532 5981 49536
rect 5917 49476 5921 49532
rect 5921 49476 5977 49532
rect 5977 49476 5981 49532
rect 5917 49472 5981 49476
rect 5997 49532 6061 49536
rect 5997 49476 6001 49532
rect 6001 49476 6057 49532
rect 6057 49476 6061 49532
rect 5997 49472 6061 49476
rect 6077 49532 6141 49536
rect 6077 49476 6081 49532
rect 6081 49476 6137 49532
rect 6137 49476 6141 49532
rect 6077 49472 6141 49476
rect 6157 49532 6221 49536
rect 6157 49476 6161 49532
rect 6161 49476 6217 49532
rect 6217 49476 6221 49532
rect 6157 49472 6221 49476
rect 15848 49532 15912 49536
rect 15848 49476 15852 49532
rect 15852 49476 15908 49532
rect 15908 49476 15912 49532
rect 15848 49472 15912 49476
rect 15928 49532 15992 49536
rect 15928 49476 15932 49532
rect 15932 49476 15988 49532
rect 15988 49476 15992 49532
rect 15928 49472 15992 49476
rect 16008 49532 16072 49536
rect 16008 49476 16012 49532
rect 16012 49476 16068 49532
rect 16068 49476 16072 49532
rect 16008 49472 16072 49476
rect 16088 49532 16152 49536
rect 16088 49476 16092 49532
rect 16092 49476 16148 49532
rect 16148 49476 16152 49532
rect 16088 49472 16152 49476
rect 25778 49532 25842 49536
rect 25778 49476 25782 49532
rect 25782 49476 25838 49532
rect 25838 49476 25842 49532
rect 25778 49472 25842 49476
rect 25858 49532 25922 49536
rect 25858 49476 25862 49532
rect 25862 49476 25918 49532
rect 25918 49476 25922 49532
rect 25858 49472 25922 49476
rect 25938 49532 26002 49536
rect 25938 49476 25942 49532
rect 25942 49476 25998 49532
rect 25998 49476 26002 49532
rect 25938 49472 26002 49476
rect 26018 49532 26082 49536
rect 26018 49476 26022 49532
rect 26022 49476 26078 49532
rect 26078 49476 26082 49532
rect 26018 49472 26082 49476
rect 26924 49464 26988 49468
rect 26924 49408 26974 49464
rect 26974 49408 26988 49464
rect 26924 49404 26988 49408
rect 27476 49464 27540 49468
rect 27476 49408 27490 49464
rect 27490 49408 27540 49464
rect 27476 49404 27540 49408
rect 10882 48988 10946 48992
rect 10882 48932 10886 48988
rect 10886 48932 10942 48988
rect 10942 48932 10946 48988
rect 10882 48928 10946 48932
rect 10962 48988 11026 48992
rect 10962 48932 10966 48988
rect 10966 48932 11022 48988
rect 11022 48932 11026 48988
rect 10962 48928 11026 48932
rect 11042 48988 11106 48992
rect 11042 48932 11046 48988
rect 11046 48932 11102 48988
rect 11102 48932 11106 48988
rect 11042 48928 11106 48932
rect 11122 48988 11186 48992
rect 11122 48932 11126 48988
rect 11126 48932 11182 48988
rect 11182 48932 11186 48988
rect 11122 48928 11186 48932
rect 20813 48988 20877 48992
rect 20813 48932 20817 48988
rect 20817 48932 20873 48988
rect 20873 48932 20877 48988
rect 20813 48928 20877 48932
rect 20893 48988 20957 48992
rect 20893 48932 20897 48988
rect 20897 48932 20953 48988
rect 20953 48932 20957 48988
rect 20893 48928 20957 48932
rect 20973 48988 21037 48992
rect 20973 48932 20977 48988
rect 20977 48932 21033 48988
rect 21033 48932 21037 48988
rect 20973 48928 21037 48932
rect 21053 48988 21117 48992
rect 21053 48932 21057 48988
rect 21057 48932 21113 48988
rect 21113 48932 21117 48988
rect 21053 48928 21117 48932
rect 24532 48860 24596 48924
rect 24164 48724 24228 48788
rect 24900 48452 24964 48516
rect 5917 48444 5981 48448
rect 5917 48388 5921 48444
rect 5921 48388 5977 48444
rect 5977 48388 5981 48444
rect 5917 48384 5981 48388
rect 5997 48444 6061 48448
rect 5997 48388 6001 48444
rect 6001 48388 6057 48444
rect 6057 48388 6061 48444
rect 5997 48384 6061 48388
rect 6077 48444 6141 48448
rect 6077 48388 6081 48444
rect 6081 48388 6137 48444
rect 6137 48388 6141 48444
rect 6077 48384 6141 48388
rect 6157 48444 6221 48448
rect 6157 48388 6161 48444
rect 6161 48388 6217 48444
rect 6217 48388 6221 48444
rect 6157 48384 6221 48388
rect 15848 48444 15912 48448
rect 15848 48388 15852 48444
rect 15852 48388 15908 48444
rect 15908 48388 15912 48444
rect 15848 48384 15912 48388
rect 15928 48444 15992 48448
rect 15928 48388 15932 48444
rect 15932 48388 15988 48444
rect 15988 48388 15992 48444
rect 15928 48384 15992 48388
rect 16008 48444 16072 48448
rect 16008 48388 16012 48444
rect 16012 48388 16068 48444
rect 16068 48388 16072 48444
rect 16008 48384 16072 48388
rect 16088 48444 16152 48448
rect 16088 48388 16092 48444
rect 16092 48388 16148 48444
rect 16148 48388 16152 48444
rect 16088 48384 16152 48388
rect 25778 48444 25842 48448
rect 25778 48388 25782 48444
rect 25782 48388 25838 48444
rect 25838 48388 25842 48444
rect 25778 48384 25842 48388
rect 25858 48444 25922 48448
rect 25858 48388 25862 48444
rect 25862 48388 25918 48444
rect 25918 48388 25922 48444
rect 25858 48384 25922 48388
rect 25938 48444 26002 48448
rect 25938 48388 25942 48444
rect 25942 48388 25998 48444
rect 25998 48388 26002 48444
rect 25938 48384 26002 48388
rect 26018 48444 26082 48448
rect 26018 48388 26022 48444
rect 26022 48388 26078 48444
rect 26078 48388 26082 48444
rect 26018 48384 26082 48388
rect 30420 49404 30484 49468
rect 31156 49268 31220 49332
rect 27476 48860 27540 48924
rect 27476 48724 27540 48788
rect 27844 48588 27908 48652
rect 28028 48452 28092 48516
rect 25268 48044 25332 48108
rect 26924 48328 26988 48380
rect 26924 48316 26938 48328
rect 26938 48316 26988 48328
rect 28948 48452 29012 48516
rect 29684 48452 29748 48516
rect 28764 48316 28828 48380
rect 29316 48316 29380 48380
rect 31524 48316 31588 48380
rect 27292 48104 27356 48108
rect 27292 48048 27306 48104
rect 27306 48048 27356 48104
rect 27292 48044 27356 48048
rect 27476 47908 27540 47972
rect 10882 47900 10946 47904
rect 10882 47844 10886 47900
rect 10886 47844 10942 47900
rect 10942 47844 10946 47900
rect 10882 47840 10946 47844
rect 10962 47900 11026 47904
rect 10962 47844 10966 47900
rect 10966 47844 11022 47900
rect 11022 47844 11026 47900
rect 10962 47840 11026 47844
rect 11042 47900 11106 47904
rect 11042 47844 11046 47900
rect 11046 47844 11102 47900
rect 11102 47844 11106 47900
rect 11042 47840 11106 47844
rect 11122 47900 11186 47904
rect 11122 47844 11126 47900
rect 11126 47844 11182 47900
rect 11182 47844 11186 47900
rect 11122 47840 11186 47844
rect 20813 47900 20877 47904
rect 20813 47844 20817 47900
rect 20817 47844 20873 47900
rect 20873 47844 20877 47900
rect 20813 47840 20877 47844
rect 20893 47900 20957 47904
rect 20893 47844 20897 47900
rect 20897 47844 20953 47900
rect 20953 47844 20957 47900
rect 20893 47840 20957 47844
rect 20973 47900 21037 47904
rect 20973 47844 20977 47900
rect 20977 47844 21033 47900
rect 21033 47844 21037 47900
rect 20973 47840 21037 47844
rect 21053 47900 21117 47904
rect 21053 47844 21057 47900
rect 21057 47844 21113 47900
rect 21113 47844 21117 47900
rect 21053 47840 21117 47844
rect 26188 47772 26252 47836
rect 28764 47908 28828 47972
rect 30052 47364 30116 47428
rect 31892 47364 31956 47428
rect 5917 47356 5981 47360
rect 5917 47300 5921 47356
rect 5921 47300 5977 47356
rect 5977 47300 5981 47356
rect 5917 47296 5981 47300
rect 5997 47356 6061 47360
rect 5997 47300 6001 47356
rect 6001 47300 6057 47356
rect 6057 47300 6061 47356
rect 5997 47296 6061 47300
rect 6077 47356 6141 47360
rect 6077 47300 6081 47356
rect 6081 47300 6137 47356
rect 6137 47300 6141 47356
rect 6077 47296 6141 47300
rect 6157 47356 6221 47360
rect 6157 47300 6161 47356
rect 6161 47300 6217 47356
rect 6217 47300 6221 47356
rect 6157 47296 6221 47300
rect 15848 47356 15912 47360
rect 15848 47300 15852 47356
rect 15852 47300 15908 47356
rect 15908 47300 15912 47356
rect 15848 47296 15912 47300
rect 15928 47356 15992 47360
rect 15928 47300 15932 47356
rect 15932 47300 15988 47356
rect 15988 47300 15992 47356
rect 15928 47296 15992 47300
rect 16008 47356 16072 47360
rect 16008 47300 16012 47356
rect 16012 47300 16068 47356
rect 16068 47300 16072 47356
rect 16008 47296 16072 47300
rect 16088 47356 16152 47360
rect 16088 47300 16092 47356
rect 16092 47300 16148 47356
rect 16148 47300 16152 47356
rect 16088 47296 16152 47300
rect 25778 47356 25842 47360
rect 25778 47300 25782 47356
rect 25782 47300 25838 47356
rect 25838 47300 25842 47356
rect 25778 47296 25842 47300
rect 25858 47356 25922 47360
rect 25858 47300 25862 47356
rect 25862 47300 25918 47356
rect 25918 47300 25922 47356
rect 25858 47296 25922 47300
rect 25938 47356 26002 47360
rect 25938 47300 25942 47356
rect 25942 47300 25998 47356
rect 25998 47300 26002 47356
rect 25938 47296 26002 47300
rect 26018 47356 26082 47360
rect 26018 47300 26022 47356
rect 26022 47300 26078 47356
rect 26078 47300 26082 47356
rect 26018 47296 26082 47300
rect 30788 47228 30852 47292
rect 26372 46820 26436 46884
rect 10882 46812 10946 46816
rect 10882 46756 10886 46812
rect 10886 46756 10942 46812
rect 10942 46756 10946 46812
rect 10882 46752 10946 46756
rect 10962 46812 11026 46816
rect 10962 46756 10966 46812
rect 10966 46756 11022 46812
rect 11022 46756 11026 46812
rect 10962 46752 11026 46756
rect 11042 46812 11106 46816
rect 11042 46756 11046 46812
rect 11046 46756 11102 46812
rect 11102 46756 11106 46812
rect 11042 46752 11106 46756
rect 11122 46812 11186 46816
rect 11122 46756 11126 46812
rect 11126 46756 11182 46812
rect 11182 46756 11186 46812
rect 11122 46752 11186 46756
rect 20813 46812 20877 46816
rect 20813 46756 20817 46812
rect 20817 46756 20873 46812
rect 20873 46756 20877 46812
rect 20813 46752 20877 46756
rect 20893 46812 20957 46816
rect 20893 46756 20897 46812
rect 20897 46756 20953 46812
rect 20953 46756 20957 46812
rect 20893 46752 20957 46756
rect 20973 46812 21037 46816
rect 20973 46756 20977 46812
rect 20977 46756 21033 46812
rect 21033 46756 21037 46812
rect 20973 46752 21037 46756
rect 21053 46812 21117 46816
rect 21053 46756 21057 46812
rect 21057 46756 21113 46812
rect 21113 46756 21117 46812
rect 21053 46752 21117 46756
rect 25268 46684 25332 46748
rect 23244 46412 23308 46476
rect 24900 46412 24964 46476
rect 26188 46412 26252 46476
rect 30604 46412 30668 46476
rect 31524 46412 31588 46476
rect 5917 46268 5981 46272
rect 5917 46212 5921 46268
rect 5921 46212 5977 46268
rect 5977 46212 5981 46268
rect 5917 46208 5981 46212
rect 5997 46268 6061 46272
rect 5997 46212 6001 46268
rect 6001 46212 6057 46268
rect 6057 46212 6061 46268
rect 5997 46208 6061 46212
rect 6077 46268 6141 46272
rect 6077 46212 6081 46268
rect 6081 46212 6137 46268
rect 6137 46212 6141 46268
rect 6077 46208 6141 46212
rect 6157 46268 6221 46272
rect 6157 46212 6161 46268
rect 6161 46212 6217 46268
rect 6217 46212 6221 46268
rect 6157 46208 6221 46212
rect 15848 46268 15912 46272
rect 15848 46212 15852 46268
rect 15852 46212 15908 46268
rect 15908 46212 15912 46268
rect 15848 46208 15912 46212
rect 15928 46268 15992 46272
rect 15928 46212 15932 46268
rect 15932 46212 15988 46268
rect 15988 46212 15992 46268
rect 15928 46208 15992 46212
rect 16008 46268 16072 46272
rect 16008 46212 16012 46268
rect 16012 46212 16068 46268
rect 16068 46212 16072 46268
rect 16008 46208 16072 46212
rect 16088 46268 16152 46272
rect 16088 46212 16092 46268
rect 16092 46212 16148 46268
rect 16148 46212 16152 46268
rect 16088 46208 16152 46212
rect 25778 46268 25842 46272
rect 25778 46212 25782 46268
rect 25782 46212 25838 46268
rect 25838 46212 25842 46268
rect 25778 46208 25842 46212
rect 25858 46268 25922 46272
rect 25858 46212 25862 46268
rect 25862 46212 25918 46268
rect 25918 46212 25922 46268
rect 25858 46208 25922 46212
rect 25938 46268 26002 46272
rect 25938 46212 25942 46268
rect 25942 46212 25998 46268
rect 25998 46212 26002 46268
rect 25938 46208 26002 46212
rect 26018 46268 26082 46272
rect 26018 46212 26022 46268
rect 26022 46212 26078 46268
rect 26078 46212 26082 46268
rect 26018 46208 26082 46212
rect 25084 46140 25148 46204
rect 27844 46140 27908 46204
rect 28948 46140 29012 46204
rect 30236 46004 30300 46068
rect 28212 45868 28276 45932
rect 10882 45724 10946 45728
rect 10882 45668 10886 45724
rect 10886 45668 10942 45724
rect 10942 45668 10946 45724
rect 10882 45664 10946 45668
rect 10962 45724 11026 45728
rect 10962 45668 10966 45724
rect 10966 45668 11022 45724
rect 11022 45668 11026 45724
rect 10962 45664 11026 45668
rect 11042 45724 11106 45728
rect 11042 45668 11046 45724
rect 11046 45668 11102 45724
rect 11102 45668 11106 45724
rect 11042 45664 11106 45668
rect 11122 45724 11186 45728
rect 11122 45668 11126 45724
rect 11126 45668 11182 45724
rect 11182 45668 11186 45724
rect 11122 45664 11186 45668
rect 20813 45724 20877 45728
rect 20813 45668 20817 45724
rect 20817 45668 20873 45724
rect 20873 45668 20877 45724
rect 20813 45664 20877 45668
rect 20893 45724 20957 45728
rect 20893 45668 20897 45724
rect 20897 45668 20953 45724
rect 20953 45668 20957 45724
rect 20893 45664 20957 45668
rect 20973 45724 21037 45728
rect 20973 45668 20977 45724
rect 20977 45668 21033 45724
rect 21033 45668 21037 45724
rect 20973 45664 21037 45668
rect 21053 45724 21117 45728
rect 21053 45668 21057 45724
rect 21057 45668 21113 45724
rect 21113 45668 21117 45724
rect 21053 45664 21117 45668
rect 28948 45596 29012 45660
rect 26924 45460 26988 45524
rect 5917 45180 5981 45184
rect 5917 45124 5921 45180
rect 5921 45124 5977 45180
rect 5977 45124 5981 45180
rect 5917 45120 5981 45124
rect 5997 45180 6061 45184
rect 5997 45124 6001 45180
rect 6001 45124 6057 45180
rect 6057 45124 6061 45180
rect 5997 45120 6061 45124
rect 6077 45180 6141 45184
rect 6077 45124 6081 45180
rect 6081 45124 6137 45180
rect 6137 45124 6141 45180
rect 6077 45120 6141 45124
rect 6157 45180 6221 45184
rect 6157 45124 6161 45180
rect 6161 45124 6217 45180
rect 6217 45124 6221 45180
rect 6157 45120 6221 45124
rect 15848 45180 15912 45184
rect 15848 45124 15852 45180
rect 15852 45124 15908 45180
rect 15908 45124 15912 45180
rect 15848 45120 15912 45124
rect 15928 45180 15992 45184
rect 15928 45124 15932 45180
rect 15932 45124 15988 45180
rect 15988 45124 15992 45180
rect 15928 45120 15992 45124
rect 16008 45180 16072 45184
rect 16008 45124 16012 45180
rect 16012 45124 16068 45180
rect 16068 45124 16072 45180
rect 16008 45120 16072 45124
rect 16088 45180 16152 45184
rect 16088 45124 16092 45180
rect 16092 45124 16148 45180
rect 16148 45124 16152 45180
rect 16088 45120 16152 45124
rect 25778 45180 25842 45184
rect 25778 45124 25782 45180
rect 25782 45124 25838 45180
rect 25838 45124 25842 45180
rect 25778 45120 25842 45124
rect 25858 45180 25922 45184
rect 25858 45124 25862 45180
rect 25862 45124 25918 45180
rect 25918 45124 25922 45180
rect 25858 45120 25922 45124
rect 25938 45180 26002 45184
rect 25938 45124 25942 45180
rect 25942 45124 25998 45180
rect 25998 45124 26002 45180
rect 25938 45120 26002 45124
rect 26018 45180 26082 45184
rect 26018 45124 26022 45180
rect 26022 45124 26078 45180
rect 26078 45124 26082 45180
rect 26018 45120 26082 45124
rect 24348 45052 24412 45116
rect 26372 45112 26436 45116
rect 26372 45056 26386 45112
rect 26386 45056 26436 45112
rect 26372 45052 26436 45056
rect 31524 45052 31588 45116
rect 27476 44644 27540 44708
rect 10882 44636 10946 44640
rect 10882 44580 10886 44636
rect 10886 44580 10942 44636
rect 10942 44580 10946 44636
rect 10882 44576 10946 44580
rect 10962 44636 11026 44640
rect 10962 44580 10966 44636
rect 10966 44580 11022 44636
rect 11022 44580 11026 44636
rect 10962 44576 11026 44580
rect 11042 44636 11106 44640
rect 11042 44580 11046 44636
rect 11046 44580 11102 44636
rect 11102 44580 11106 44636
rect 11042 44576 11106 44580
rect 11122 44636 11186 44640
rect 11122 44580 11126 44636
rect 11126 44580 11182 44636
rect 11182 44580 11186 44636
rect 11122 44576 11186 44580
rect 20813 44636 20877 44640
rect 20813 44580 20817 44636
rect 20817 44580 20873 44636
rect 20873 44580 20877 44636
rect 20813 44576 20877 44580
rect 20893 44636 20957 44640
rect 20893 44580 20897 44636
rect 20897 44580 20953 44636
rect 20953 44580 20957 44636
rect 20893 44576 20957 44580
rect 20973 44636 21037 44640
rect 20973 44580 20977 44636
rect 20977 44580 21033 44636
rect 21033 44580 21037 44636
rect 20973 44576 21037 44580
rect 21053 44636 21117 44640
rect 21053 44580 21057 44636
rect 21057 44580 21113 44636
rect 21113 44580 21117 44636
rect 21053 44576 21117 44580
rect 27292 44508 27356 44572
rect 27660 44372 27724 44436
rect 28764 44508 28828 44572
rect 30236 44508 30300 44572
rect 28764 44236 28828 44300
rect 29684 44236 29748 44300
rect 31708 44100 31772 44164
rect 5917 44092 5981 44096
rect 5917 44036 5921 44092
rect 5921 44036 5977 44092
rect 5977 44036 5981 44092
rect 5917 44032 5981 44036
rect 5997 44092 6061 44096
rect 5997 44036 6001 44092
rect 6001 44036 6057 44092
rect 6057 44036 6061 44092
rect 5997 44032 6061 44036
rect 6077 44092 6141 44096
rect 6077 44036 6081 44092
rect 6081 44036 6137 44092
rect 6137 44036 6141 44092
rect 6077 44032 6141 44036
rect 6157 44092 6221 44096
rect 6157 44036 6161 44092
rect 6161 44036 6217 44092
rect 6217 44036 6221 44092
rect 6157 44032 6221 44036
rect 15848 44092 15912 44096
rect 15848 44036 15852 44092
rect 15852 44036 15908 44092
rect 15908 44036 15912 44092
rect 15848 44032 15912 44036
rect 15928 44092 15992 44096
rect 15928 44036 15932 44092
rect 15932 44036 15988 44092
rect 15988 44036 15992 44092
rect 15928 44032 15992 44036
rect 16008 44092 16072 44096
rect 16008 44036 16012 44092
rect 16012 44036 16068 44092
rect 16068 44036 16072 44092
rect 16008 44032 16072 44036
rect 16088 44092 16152 44096
rect 16088 44036 16092 44092
rect 16092 44036 16148 44092
rect 16148 44036 16152 44092
rect 16088 44032 16152 44036
rect 25778 44092 25842 44096
rect 25778 44036 25782 44092
rect 25782 44036 25838 44092
rect 25838 44036 25842 44092
rect 25778 44032 25842 44036
rect 25858 44092 25922 44096
rect 25858 44036 25862 44092
rect 25862 44036 25918 44092
rect 25918 44036 25922 44092
rect 25858 44032 25922 44036
rect 25938 44092 26002 44096
rect 25938 44036 25942 44092
rect 25942 44036 25998 44092
rect 25998 44036 26002 44092
rect 25938 44032 26002 44036
rect 26018 44092 26082 44096
rect 26018 44036 26022 44092
rect 26022 44036 26078 44092
rect 26078 44036 26082 44092
rect 26018 44032 26082 44036
rect 30972 43556 31036 43620
rect 10882 43548 10946 43552
rect 10882 43492 10886 43548
rect 10886 43492 10942 43548
rect 10942 43492 10946 43548
rect 10882 43488 10946 43492
rect 10962 43548 11026 43552
rect 10962 43492 10966 43548
rect 10966 43492 11022 43548
rect 11022 43492 11026 43548
rect 10962 43488 11026 43492
rect 11042 43548 11106 43552
rect 11042 43492 11046 43548
rect 11046 43492 11102 43548
rect 11102 43492 11106 43548
rect 11042 43488 11106 43492
rect 11122 43548 11186 43552
rect 11122 43492 11126 43548
rect 11126 43492 11182 43548
rect 11182 43492 11186 43548
rect 11122 43488 11186 43492
rect 20813 43548 20877 43552
rect 20813 43492 20817 43548
rect 20817 43492 20873 43548
rect 20873 43492 20877 43548
rect 20813 43488 20877 43492
rect 20893 43548 20957 43552
rect 20893 43492 20897 43548
rect 20897 43492 20953 43548
rect 20953 43492 20957 43548
rect 20893 43488 20957 43492
rect 20973 43548 21037 43552
rect 20973 43492 20977 43548
rect 20977 43492 21033 43548
rect 21033 43492 21037 43548
rect 20973 43488 21037 43492
rect 21053 43548 21117 43552
rect 21053 43492 21057 43548
rect 21057 43492 21113 43548
rect 21113 43492 21117 43548
rect 21053 43488 21117 43492
rect 21404 43284 21468 43348
rect 23980 43208 24044 43212
rect 23980 43152 24030 43208
rect 24030 43152 24044 43208
rect 23980 43148 24044 43152
rect 24716 43208 24780 43212
rect 24716 43152 24766 43208
rect 24766 43152 24780 43208
rect 24716 43148 24780 43152
rect 27660 43148 27724 43212
rect 5917 43004 5981 43008
rect 5917 42948 5921 43004
rect 5921 42948 5977 43004
rect 5977 42948 5981 43004
rect 5917 42944 5981 42948
rect 5997 43004 6061 43008
rect 5997 42948 6001 43004
rect 6001 42948 6057 43004
rect 6057 42948 6061 43004
rect 5997 42944 6061 42948
rect 6077 43004 6141 43008
rect 6077 42948 6081 43004
rect 6081 42948 6137 43004
rect 6137 42948 6141 43004
rect 6077 42944 6141 42948
rect 6157 43004 6221 43008
rect 6157 42948 6161 43004
rect 6161 42948 6217 43004
rect 6217 42948 6221 43004
rect 6157 42944 6221 42948
rect 15848 43004 15912 43008
rect 15848 42948 15852 43004
rect 15852 42948 15908 43004
rect 15908 42948 15912 43004
rect 15848 42944 15912 42948
rect 15928 43004 15992 43008
rect 15928 42948 15932 43004
rect 15932 42948 15988 43004
rect 15988 42948 15992 43004
rect 15928 42944 15992 42948
rect 16008 43004 16072 43008
rect 16008 42948 16012 43004
rect 16012 42948 16068 43004
rect 16068 42948 16072 43004
rect 16008 42944 16072 42948
rect 16088 43004 16152 43008
rect 16088 42948 16092 43004
rect 16092 42948 16148 43004
rect 16148 42948 16152 43004
rect 16088 42944 16152 42948
rect 25778 43004 25842 43008
rect 25778 42948 25782 43004
rect 25782 42948 25838 43004
rect 25838 42948 25842 43004
rect 25778 42944 25842 42948
rect 25858 43004 25922 43008
rect 25858 42948 25862 43004
rect 25862 42948 25918 43004
rect 25918 42948 25922 43004
rect 25858 42944 25922 42948
rect 25938 43004 26002 43008
rect 25938 42948 25942 43004
rect 25942 42948 25998 43004
rect 25998 42948 26002 43004
rect 25938 42944 26002 42948
rect 26018 43004 26082 43008
rect 26018 42948 26022 43004
rect 26022 42948 26078 43004
rect 26078 42948 26082 43004
rect 26018 42944 26082 42948
rect 25268 42876 25332 42940
rect 26188 42740 26252 42804
rect 25268 42604 25332 42668
rect 27108 42604 27172 42668
rect 10882 42460 10946 42464
rect 10882 42404 10886 42460
rect 10886 42404 10942 42460
rect 10942 42404 10946 42460
rect 10882 42400 10946 42404
rect 10962 42460 11026 42464
rect 10962 42404 10966 42460
rect 10966 42404 11022 42460
rect 11022 42404 11026 42460
rect 10962 42400 11026 42404
rect 11042 42460 11106 42464
rect 11042 42404 11046 42460
rect 11046 42404 11102 42460
rect 11102 42404 11106 42460
rect 11042 42400 11106 42404
rect 11122 42460 11186 42464
rect 11122 42404 11126 42460
rect 11126 42404 11182 42460
rect 11182 42404 11186 42460
rect 11122 42400 11186 42404
rect 20813 42460 20877 42464
rect 20813 42404 20817 42460
rect 20817 42404 20873 42460
rect 20873 42404 20877 42460
rect 20813 42400 20877 42404
rect 20893 42460 20957 42464
rect 20893 42404 20897 42460
rect 20897 42404 20953 42460
rect 20953 42404 20957 42460
rect 20893 42400 20957 42404
rect 20973 42460 21037 42464
rect 20973 42404 20977 42460
rect 20977 42404 21033 42460
rect 21033 42404 21037 42460
rect 20973 42400 21037 42404
rect 21053 42460 21117 42464
rect 21053 42404 21057 42460
rect 21057 42404 21113 42460
rect 21113 42404 21117 42460
rect 21053 42400 21117 42404
rect 23244 42392 23308 42396
rect 23244 42336 23294 42392
rect 23294 42336 23308 42392
rect 23244 42332 23308 42336
rect 26188 42332 26252 42396
rect 24716 42196 24780 42260
rect 5917 41916 5981 41920
rect 5917 41860 5921 41916
rect 5921 41860 5977 41916
rect 5977 41860 5981 41916
rect 5917 41856 5981 41860
rect 5997 41916 6061 41920
rect 5997 41860 6001 41916
rect 6001 41860 6057 41916
rect 6057 41860 6061 41916
rect 5997 41856 6061 41860
rect 6077 41916 6141 41920
rect 6077 41860 6081 41916
rect 6081 41860 6137 41916
rect 6137 41860 6141 41916
rect 6077 41856 6141 41860
rect 6157 41916 6221 41920
rect 6157 41860 6161 41916
rect 6161 41860 6217 41916
rect 6217 41860 6221 41916
rect 6157 41856 6221 41860
rect 15848 41916 15912 41920
rect 15848 41860 15852 41916
rect 15852 41860 15908 41916
rect 15908 41860 15912 41916
rect 15848 41856 15912 41860
rect 15928 41916 15992 41920
rect 15928 41860 15932 41916
rect 15932 41860 15988 41916
rect 15988 41860 15992 41916
rect 15928 41856 15992 41860
rect 16008 41916 16072 41920
rect 16008 41860 16012 41916
rect 16012 41860 16068 41916
rect 16068 41860 16072 41916
rect 16008 41856 16072 41860
rect 16088 41916 16152 41920
rect 16088 41860 16092 41916
rect 16092 41860 16148 41916
rect 16148 41860 16152 41916
rect 16088 41856 16152 41860
rect 25778 41916 25842 41920
rect 25778 41860 25782 41916
rect 25782 41860 25838 41916
rect 25838 41860 25842 41916
rect 25778 41856 25842 41860
rect 25858 41916 25922 41920
rect 25858 41860 25862 41916
rect 25862 41860 25918 41916
rect 25918 41860 25922 41916
rect 25858 41856 25922 41860
rect 25938 41916 26002 41920
rect 25938 41860 25942 41916
rect 25942 41860 25998 41916
rect 25998 41860 26002 41916
rect 25938 41856 26002 41860
rect 26018 41916 26082 41920
rect 26018 41860 26022 41916
rect 26022 41860 26078 41916
rect 26078 41860 26082 41916
rect 26018 41856 26082 41860
rect 29868 43012 29932 43076
rect 30052 43012 30116 43076
rect 30420 43284 30484 43348
rect 30788 43148 30852 43212
rect 31340 43148 31404 43212
rect 30420 43012 30484 43076
rect 29868 42740 29932 42804
rect 30972 42604 31036 42668
rect 29132 42332 29196 42396
rect 29132 42256 29196 42260
rect 29132 42200 29182 42256
rect 29182 42200 29196 42256
rect 29132 42196 29196 42200
rect 10882 41372 10946 41376
rect 10882 41316 10886 41372
rect 10886 41316 10942 41372
rect 10942 41316 10946 41372
rect 10882 41312 10946 41316
rect 10962 41372 11026 41376
rect 10962 41316 10966 41372
rect 10966 41316 11022 41372
rect 11022 41316 11026 41372
rect 10962 41312 11026 41316
rect 11042 41372 11106 41376
rect 11042 41316 11046 41372
rect 11046 41316 11102 41372
rect 11102 41316 11106 41372
rect 11042 41312 11106 41316
rect 11122 41372 11186 41376
rect 11122 41316 11126 41372
rect 11126 41316 11182 41372
rect 11182 41316 11186 41372
rect 11122 41312 11186 41316
rect 20813 41372 20877 41376
rect 20813 41316 20817 41372
rect 20817 41316 20873 41372
rect 20873 41316 20877 41372
rect 20813 41312 20877 41316
rect 20893 41372 20957 41376
rect 20893 41316 20897 41372
rect 20897 41316 20953 41372
rect 20953 41316 20957 41372
rect 20893 41312 20957 41316
rect 20973 41372 21037 41376
rect 20973 41316 20977 41372
rect 20977 41316 21033 41372
rect 21033 41316 21037 41372
rect 20973 41312 21037 41316
rect 21053 41372 21117 41376
rect 21053 41316 21057 41372
rect 21057 41316 21113 41372
rect 21113 41316 21117 41372
rect 21053 41312 21117 41316
rect 24164 41516 24228 41580
rect 25268 41576 25332 41580
rect 25268 41520 25318 41576
rect 25318 41520 25332 41576
rect 25268 41516 25332 41520
rect 26372 41516 26436 41580
rect 26924 41576 26988 41580
rect 26924 41520 26938 41576
rect 26938 41520 26988 41576
rect 26924 41516 26988 41520
rect 24348 41380 24412 41444
rect 26372 41380 26436 41444
rect 26740 41380 26804 41444
rect 24900 41244 24964 41308
rect 28212 41712 28276 41716
rect 28212 41656 28226 41712
rect 28226 41656 28276 41712
rect 28212 41652 28276 41656
rect 24348 41108 24412 41172
rect 25452 41168 25516 41172
rect 25452 41112 25466 41168
rect 25466 41112 25516 41168
rect 25452 41108 25516 41112
rect 26924 41168 26988 41172
rect 26924 41112 26974 41168
rect 26974 41112 26988 41168
rect 26924 41108 26988 41112
rect 30052 41652 30116 41716
rect 30788 41712 30852 41716
rect 30788 41656 30802 41712
rect 30802 41656 30852 41712
rect 30788 41652 30852 41656
rect 30788 41576 30852 41580
rect 30788 41520 30838 41576
rect 30838 41520 30852 41576
rect 30788 41516 30852 41520
rect 28028 41244 28092 41308
rect 30604 41108 30668 41172
rect 25452 40836 25516 40900
rect 5917 40828 5981 40832
rect 5917 40772 5921 40828
rect 5921 40772 5977 40828
rect 5977 40772 5981 40828
rect 5917 40768 5981 40772
rect 5997 40828 6061 40832
rect 5997 40772 6001 40828
rect 6001 40772 6057 40828
rect 6057 40772 6061 40828
rect 5997 40768 6061 40772
rect 6077 40828 6141 40832
rect 6077 40772 6081 40828
rect 6081 40772 6137 40828
rect 6137 40772 6141 40828
rect 6077 40768 6141 40772
rect 6157 40828 6221 40832
rect 6157 40772 6161 40828
rect 6161 40772 6217 40828
rect 6217 40772 6221 40828
rect 6157 40768 6221 40772
rect 15848 40828 15912 40832
rect 15848 40772 15852 40828
rect 15852 40772 15908 40828
rect 15908 40772 15912 40828
rect 15848 40768 15912 40772
rect 15928 40828 15992 40832
rect 15928 40772 15932 40828
rect 15932 40772 15988 40828
rect 15988 40772 15992 40828
rect 15928 40768 15992 40772
rect 16008 40828 16072 40832
rect 16008 40772 16012 40828
rect 16012 40772 16068 40828
rect 16068 40772 16072 40828
rect 16008 40768 16072 40772
rect 16088 40828 16152 40832
rect 16088 40772 16092 40828
rect 16092 40772 16148 40828
rect 16148 40772 16152 40828
rect 16088 40768 16152 40772
rect 27660 41032 27724 41036
rect 27660 40976 27710 41032
rect 27710 40976 27724 41032
rect 27660 40972 27724 40976
rect 27292 40836 27356 40900
rect 27660 40836 27724 40900
rect 29132 40972 29196 41036
rect 25778 40828 25842 40832
rect 25778 40772 25782 40828
rect 25782 40772 25838 40828
rect 25838 40772 25842 40828
rect 25778 40768 25842 40772
rect 25858 40828 25922 40832
rect 25858 40772 25862 40828
rect 25862 40772 25918 40828
rect 25918 40772 25922 40828
rect 25858 40768 25922 40772
rect 25938 40828 26002 40832
rect 25938 40772 25942 40828
rect 25942 40772 25998 40828
rect 25998 40772 26002 40828
rect 25938 40768 26002 40772
rect 26018 40828 26082 40832
rect 26018 40772 26022 40828
rect 26022 40772 26078 40828
rect 26078 40772 26082 40828
rect 26018 40768 26082 40772
rect 30788 40700 30852 40764
rect 25636 40292 25700 40356
rect 10882 40284 10946 40288
rect 10882 40228 10886 40284
rect 10886 40228 10942 40284
rect 10942 40228 10946 40284
rect 10882 40224 10946 40228
rect 10962 40284 11026 40288
rect 10962 40228 10966 40284
rect 10966 40228 11022 40284
rect 11022 40228 11026 40284
rect 10962 40224 11026 40228
rect 11042 40284 11106 40288
rect 11042 40228 11046 40284
rect 11046 40228 11102 40284
rect 11102 40228 11106 40284
rect 11042 40224 11106 40228
rect 11122 40284 11186 40288
rect 11122 40228 11126 40284
rect 11126 40228 11182 40284
rect 11182 40228 11186 40284
rect 11122 40224 11186 40228
rect 20813 40284 20877 40288
rect 20813 40228 20817 40284
rect 20817 40228 20873 40284
rect 20873 40228 20877 40284
rect 20813 40224 20877 40228
rect 20893 40284 20957 40288
rect 20893 40228 20897 40284
rect 20897 40228 20953 40284
rect 20953 40228 20957 40284
rect 20893 40224 20957 40228
rect 20973 40284 21037 40288
rect 20973 40228 20977 40284
rect 20977 40228 21033 40284
rect 21033 40228 21037 40284
rect 20973 40224 21037 40228
rect 21053 40284 21117 40288
rect 21053 40228 21057 40284
rect 21057 40228 21113 40284
rect 21113 40228 21117 40284
rect 21053 40224 21117 40228
rect 30052 40428 30116 40492
rect 27476 40020 27540 40084
rect 24164 39884 24228 39948
rect 30788 39884 30852 39948
rect 31892 39884 31956 39948
rect 27108 39748 27172 39812
rect 5917 39740 5981 39744
rect 5917 39684 5921 39740
rect 5921 39684 5977 39740
rect 5977 39684 5981 39740
rect 5917 39680 5981 39684
rect 5997 39740 6061 39744
rect 5997 39684 6001 39740
rect 6001 39684 6057 39740
rect 6057 39684 6061 39740
rect 5997 39680 6061 39684
rect 6077 39740 6141 39744
rect 6077 39684 6081 39740
rect 6081 39684 6137 39740
rect 6137 39684 6141 39740
rect 6077 39680 6141 39684
rect 6157 39740 6221 39744
rect 6157 39684 6161 39740
rect 6161 39684 6217 39740
rect 6217 39684 6221 39740
rect 6157 39680 6221 39684
rect 15848 39740 15912 39744
rect 15848 39684 15852 39740
rect 15852 39684 15908 39740
rect 15908 39684 15912 39740
rect 15848 39680 15912 39684
rect 15928 39740 15992 39744
rect 15928 39684 15932 39740
rect 15932 39684 15988 39740
rect 15988 39684 15992 39740
rect 15928 39680 15992 39684
rect 16008 39740 16072 39744
rect 16008 39684 16012 39740
rect 16012 39684 16068 39740
rect 16068 39684 16072 39740
rect 16008 39680 16072 39684
rect 16088 39740 16152 39744
rect 16088 39684 16092 39740
rect 16092 39684 16148 39740
rect 16148 39684 16152 39740
rect 16088 39680 16152 39684
rect 25778 39740 25842 39744
rect 25778 39684 25782 39740
rect 25782 39684 25838 39740
rect 25838 39684 25842 39740
rect 25778 39680 25842 39684
rect 25858 39740 25922 39744
rect 25858 39684 25862 39740
rect 25862 39684 25918 39740
rect 25918 39684 25922 39740
rect 25858 39680 25922 39684
rect 25938 39740 26002 39744
rect 25938 39684 25942 39740
rect 25942 39684 25998 39740
rect 25998 39684 26002 39740
rect 25938 39680 26002 39684
rect 26018 39740 26082 39744
rect 26018 39684 26022 39740
rect 26022 39684 26078 39740
rect 26078 39684 26082 39740
rect 26018 39680 26082 39684
rect 26188 39536 26252 39540
rect 26188 39480 26202 39536
rect 26202 39480 26252 39536
rect 26188 39476 26252 39480
rect 26372 39340 26436 39404
rect 29132 39340 29196 39404
rect 30420 39340 30484 39404
rect 26372 39264 26436 39268
rect 26372 39208 26422 39264
rect 26422 39208 26436 39264
rect 26372 39204 26436 39208
rect 10882 39196 10946 39200
rect 10882 39140 10886 39196
rect 10886 39140 10942 39196
rect 10942 39140 10946 39196
rect 10882 39136 10946 39140
rect 10962 39196 11026 39200
rect 10962 39140 10966 39196
rect 10966 39140 11022 39196
rect 11022 39140 11026 39196
rect 10962 39136 11026 39140
rect 11042 39196 11106 39200
rect 11042 39140 11046 39196
rect 11046 39140 11102 39196
rect 11102 39140 11106 39196
rect 11042 39136 11106 39140
rect 11122 39196 11186 39200
rect 11122 39140 11126 39196
rect 11126 39140 11182 39196
rect 11182 39140 11186 39196
rect 11122 39136 11186 39140
rect 20813 39196 20877 39200
rect 20813 39140 20817 39196
rect 20817 39140 20873 39196
rect 20873 39140 20877 39196
rect 20813 39136 20877 39140
rect 20893 39196 20957 39200
rect 20893 39140 20897 39196
rect 20897 39140 20953 39196
rect 20953 39140 20957 39196
rect 20893 39136 20957 39140
rect 20973 39196 21037 39200
rect 20973 39140 20977 39196
rect 20977 39140 21033 39196
rect 21033 39140 21037 39196
rect 20973 39136 21037 39140
rect 21053 39196 21117 39200
rect 21053 39140 21057 39196
rect 21057 39140 21113 39196
rect 21113 39140 21117 39196
rect 21053 39136 21117 39140
rect 23612 38932 23676 38996
rect 26188 38932 26252 38996
rect 25636 38796 25700 38860
rect 5917 38652 5981 38656
rect 5917 38596 5921 38652
rect 5921 38596 5977 38652
rect 5977 38596 5981 38652
rect 5917 38592 5981 38596
rect 5997 38652 6061 38656
rect 5997 38596 6001 38652
rect 6001 38596 6057 38652
rect 6057 38596 6061 38652
rect 5997 38592 6061 38596
rect 6077 38652 6141 38656
rect 6077 38596 6081 38652
rect 6081 38596 6137 38652
rect 6137 38596 6141 38652
rect 6077 38592 6141 38596
rect 6157 38652 6221 38656
rect 6157 38596 6161 38652
rect 6161 38596 6217 38652
rect 6217 38596 6221 38652
rect 6157 38592 6221 38596
rect 15848 38652 15912 38656
rect 15848 38596 15852 38652
rect 15852 38596 15908 38652
rect 15908 38596 15912 38652
rect 15848 38592 15912 38596
rect 15928 38652 15992 38656
rect 15928 38596 15932 38652
rect 15932 38596 15988 38652
rect 15988 38596 15992 38652
rect 15928 38592 15992 38596
rect 16008 38652 16072 38656
rect 16008 38596 16012 38652
rect 16012 38596 16068 38652
rect 16068 38596 16072 38652
rect 16008 38592 16072 38596
rect 16088 38652 16152 38656
rect 16088 38596 16092 38652
rect 16092 38596 16148 38652
rect 16148 38596 16152 38652
rect 16088 38592 16152 38596
rect 30420 38932 30484 38996
rect 31708 38932 31772 38996
rect 25778 38652 25842 38656
rect 25778 38596 25782 38652
rect 25782 38596 25838 38652
rect 25838 38596 25842 38652
rect 25778 38592 25842 38596
rect 25858 38652 25922 38656
rect 25858 38596 25862 38652
rect 25862 38596 25918 38652
rect 25918 38596 25922 38652
rect 25858 38592 25922 38596
rect 25938 38652 26002 38656
rect 25938 38596 25942 38652
rect 25942 38596 25998 38652
rect 25998 38596 26002 38652
rect 25938 38592 26002 38596
rect 26018 38652 26082 38656
rect 26018 38596 26022 38652
rect 26022 38596 26078 38652
rect 26078 38596 26082 38652
rect 26018 38592 26082 38596
rect 25268 38524 25332 38588
rect 26372 38584 26436 38588
rect 26372 38528 26422 38584
rect 26422 38528 26436 38584
rect 26372 38524 26436 38528
rect 24900 38388 24964 38452
rect 28028 38448 28092 38452
rect 28028 38392 28042 38448
rect 28042 38392 28092 38448
rect 28028 38388 28092 38392
rect 24532 38252 24596 38316
rect 10882 38108 10946 38112
rect 10882 38052 10886 38108
rect 10886 38052 10942 38108
rect 10942 38052 10946 38108
rect 10882 38048 10946 38052
rect 10962 38108 11026 38112
rect 10962 38052 10966 38108
rect 10966 38052 11022 38108
rect 11022 38052 11026 38108
rect 10962 38048 11026 38052
rect 11042 38108 11106 38112
rect 11042 38052 11046 38108
rect 11046 38052 11102 38108
rect 11102 38052 11106 38108
rect 11042 38048 11106 38052
rect 11122 38108 11186 38112
rect 11122 38052 11126 38108
rect 11126 38052 11182 38108
rect 11182 38052 11186 38108
rect 11122 38048 11186 38052
rect 20813 38108 20877 38112
rect 20813 38052 20817 38108
rect 20817 38052 20873 38108
rect 20873 38052 20877 38108
rect 20813 38048 20877 38052
rect 20893 38108 20957 38112
rect 20893 38052 20897 38108
rect 20897 38052 20953 38108
rect 20953 38052 20957 38108
rect 20893 38048 20957 38052
rect 20973 38108 21037 38112
rect 20973 38052 20977 38108
rect 20977 38052 21033 38108
rect 21033 38052 21037 38108
rect 20973 38048 21037 38052
rect 21053 38108 21117 38112
rect 21053 38052 21057 38108
rect 21057 38052 21113 38108
rect 21113 38052 21117 38108
rect 21053 38048 21117 38052
rect 23612 38040 23676 38044
rect 23612 37984 23626 38040
rect 23626 37984 23676 38040
rect 23612 37980 23676 37984
rect 25084 38116 25148 38180
rect 25452 38116 25516 38180
rect 26924 38116 26988 38180
rect 28028 38116 28092 38180
rect 31156 37980 31220 38044
rect 31340 37980 31404 38044
rect 25452 37844 25516 37908
rect 26188 37844 26252 37908
rect 23980 37768 24044 37772
rect 23980 37712 24030 37768
rect 24030 37712 24044 37768
rect 23980 37708 24044 37712
rect 27476 37708 27540 37772
rect 24900 37632 24964 37636
rect 24900 37576 24914 37632
rect 24914 37576 24964 37632
rect 24900 37572 24964 37576
rect 5917 37564 5981 37568
rect 5917 37508 5921 37564
rect 5921 37508 5977 37564
rect 5977 37508 5981 37564
rect 5917 37504 5981 37508
rect 5997 37564 6061 37568
rect 5997 37508 6001 37564
rect 6001 37508 6057 37564
rect 6057 37508 6061 37564
rect 5997 37504 6061 37508
rect 6077 37564 6141 37568
rect 6077 37508 6081 37564
rect 6081 37508 6137 37564
rect 6137 37508 6141 37564
rect 6077 37504 6141 37508
rect 6157 37564 6221 37568
rect 6157 37508 6161 37564
rect 6161 37508 6217 37564
rect 6217 37508 6221 37564
rect 6157 37504 6221 37508
rect 15848 37564 15912 37568
rect 15848 37508 15852 37564
rect 15852 37508 15908 37564
rect 15908 37508 15912 37564
rect 15848 37504 15912 37508
rect 15928 37564 15992 37568
rect 15928 37508 15932 37564
rect 15932 37508 15988 37564
rect 15988 37508 15992 37564
rect 15928 37504 15992 37508
rect 16008 37564 16072 37568
rect 16008 37508 16012 37564
rect 16012 37508 16068 37564
rect 16068 37508 16072 37564
rect 16008 37504 16072 37508
rect 16088 37564 16152 37568
rect 16088 37508 16092 37564
rect 16092 37508 16148 37564
rect 16148 37508 16152 37564
rect 16088 37504 16152 37508
rect 25778 37564 25842 37568
rect 25778 37508 25782 37564
rect 25782 37508 25838 37564
rect 25838 37508 25842 37564
rect 25778 37504 25842 37508
rect 25858 37564 25922 37568
rect 25858 37508 25862 37564
rect 25862 37508 25918 37564
rect 25918 37508 25922 37564
rect 25858 37504 25922 37508
rect 25938 37564 26002 37568
rect 25938 37508 25942 37564
rect 25942 37508 25998 37564
rect 25998 37508 26002 37564
rect 25938 37504 26002 37508
rect 26018 37564 26082 37568
rect 26018 37508 26022 37564
rect 26022 37508 26078 37564
rect 26078 37508 26082 37564
rect 26018 37504 26082 37508
rect 24716 37436 24780 37500
rect 26924 37436 26988 37500
rect 26372 37300 26436 37364
rect 25268 37164 25332 37228
rect 30420 37164 30484 37228
rect 26740 37028 26804 37092
rect 31156 37028 31220 37092
rect 10882 37020 10946 37024
rect 10882 36964 10886 37020
rect 10886 36964 10942 37020
rect 10942 36964 10946 37020
rect 10882 36960 10946 36964
rect 10962 37020 11026 37024
rect 10962 36964 10966 37020
rect 10966 36964 11022 37020
rect 11022 36964 11026 37020
rect 10962 36960 11026 36964
rect 11042 37020 11106 37024
rect 11042 36964 11046 37020
rect 11046 36964 11102 37020
rect 11102 36964 11106 37020
rect 11042 36960 11106 36964
rect 11122 37020 11186 37024
rect 11122 36964 11126 37020
rect 11126 36964 11182 37020
rect 11182 36964 11186 37020
rect 11122 36960 11186 36964
rect 20813 37020 20877 37024
rect 20813 36964 20817 37020
rect 20817 36964 20873 37020
rect 20873 36964 20877 37020
rect 20813 36960 20877 36964
rect 20893 37020 20957 37024
rect 20893 36964 20897 37020
rect 20897 36964 20953 37020
rect 20953 36964 20957 37020
rect 20893 36960 20957 36964
rect 20973 37020 21037 37024
rect 20973 36964 20977 37020
rect 20977 36964 21033 37020
rect 21033 36964 21037 37020
rect 20973 36960 21037 36964
rect 21053 37020 21117 37024
rect 21053 36964 21057 37020
rect 21057 36964 21113 37020
rect 21113 36964 21117 37020
rect 21053 36960 21117 36964
rect 24900 36620 24964 36684
rect 26556 36620 26620 36684
rect 30052 36680 30116 36684
rect 30052 36624 30066 36680
rect 30066 36624 30116 36680
rect 30052 36620 30116 36624
rect 5917 36476 5981 36480
rect 5917 36420 5921 36476
rect 5921 36420 5977 36476
rect 5977 36420 5981 36476
rect 5917 36416 5981 36420
rect 5997 36476 6061 36480
rect 5997 36420 6001 36476
rect 6001 36420 6057 36476
rect 6057 36420 6061 36476
rect 5997 36416 6061 36420
rect 6077 36476 6141 36480
rect 6077 36420 6081 36476
rect 6081 36420 6137 36476
rect 6137 36420 6141 36476
rect 6077 36416 6141 36420
rect 6157 36476 6221 36480
rect 6157 36420 6161 36476
rect 6161 36420 6217 36476
rect 6217 36420 6221 36476
rect 6157 36416 6221 36420
rect 15848 36476 15912 36480
rect 15848 36420 15852 36476
rect 15852 36420 15908 36476
rect 15908 36420 15912 36476
rect 15848 36416 15912 36420
rect 15928 36476 15992 36480
rect 15928 36420 15932 36476
rect 15932 36420 15988 36476
rect 15988 36420 15992 36476
rect 15928 36416 15992 36420
rect 16008 36476 16072 36480
rect 16008 36420 16012 36476
rect 16012 36420 16068 36476
rect 16068 36420 16072 36476
rect 16008 36416 16072 36420
rect 16088 36476 16152 36480
rect 16088 36420 16092 36476
rect 16092 36420 16148 36476
rect 16148 36420 16152 36476
rect 16088 36416 16152 36420
rect 25778 36476 25842 36480
rect 25778 36420 25782 36476
rect 25782 36420 25838 36476
rect 25838 36420 25842 36476
rect 25778 36416 25842 36420
rect 25858 36476 25922 36480
rect 25858 36420 25862 36476
rect 25862 36420 25918 36476
rect 25918 36420 25922 36476
rect 25858 36416 25922 36420
rect 25938 36476 26002 36480
rect 25938 36420 25942 36476
rect 25942 36420 25998 36476
rect 25998 36420 26002 36476
rect 25938 36416 26002 36420
rect 26018 36476 26082 36480
rect 26018 36420 26022 36476
rect 26022 36420 26078 36476
rect 26078 36420 26082 36476
rect 26018 36416 26082 36420
rect 30972 36212 31036 36276
rect 25452 36076 25516 36140
rect 31524 36076 31588 36140
rect 25452 35940 25516 36004
rect 10882 35932 10946 35936
rect 10882 35876 10886 35932
rect 10886 35876 10942 35932
rect 10942 35876 10946 35932
rect 10882 35872 10946 35876
rect 10962 35932 11026 35936
rect 10962 35876 10966 35932
rect 10966 35876 11022 35932
rect 11022 35876 11026 35932
rect 10962 35872 11026 35876
rect 11042 35932 11106 35936
rect 11042 35876 11046 35932
rect 11046 35876 11102 35932
rect 11102 35876 11106 35932
rect 11042 35872 11106 35876
rect 11122 35932 11186 35936
rect 11122 35876 11126 35932
rect 11126 35876 11182 35932
rect 11182 35876 11186 35932
rect 11122 35872 11186 35876
rect 20813 35932 20877 35936
rect 20813 35876 20817 35932
rect 20817 35876 20873 35932
rect 20873 35876 20877 35932
rect 20813 35872 20877 35876
rect 20893 35932 20957 35936
rect 20893 35876 20897 35932
rect 20897 35876 20953 35932
rect 20953 35876 20957 35932
rect 20893 35872 20957 35876
rect 20973 35932 21037 35936
rect 20973 35876 20977 35932
rect 20977 35876 21033 35932
rect 21033 35876 21037 35932
rect 20973 35872 21037 35876
rect 21053 35932 21117 35936
rect 21053 35876 21057 35932
rect 21057 35876 21113 35932
rect 21113 35876 21117 35932
rect 21053 35872 21117 35876
rect 25084 35804 25148 35868
rect 25268 35668 25332 35732
rect 5917 35388 5981 35392
rect 5917 35332 5921 35388
rect 5921 35332 5977 35388
rect 5977 35332 5981 35388
rect 5917 35328 5981 35332
rect 5997 35388 6061 35392
rect 5997 35332 6001 35388
rect 6001 35332 6057 35388
rect 6057 35332 6061 35388
rect 5997 35328 6061 35332
rect 6077 35388 6141 35392
rect 6077 35332 6081 35388
rect 6081 35332 6137 35388
rect 6137 35332 6141 35388
rect 6077 35328 6141 35332
rect 6157 35388 6221 35392
rect 6157 35332 6161 35388
rect 6161 35332 6217 35388
rect 6217 35332 6221 35388
rect 6157 35328 6221 35332
rect 15848 35388 15912 35392
rect 15848 35332 15852 35388
rect 15852 35332 15908 35388
rect 15908 35332 15912 35388
rect 15848 35328 15912 35332
rect 15928 35388 15992 35392
rect 15928 35332 15932 35388
rect 15932 35332 15988 35388
rect 15988 35332 15992 35388
rect 15928 35328 15992 35332
rect 16008 35388 16072 35392
rect 16008 35332 16012 35388
rect 16012 35332 16068 35388
rect 16068 35332 16072 35388
rect 16008 35328 16072 35332
rect 16088 35388 16152 35392
rect 16088 35332 16092 35388
rect 16092 35332 16148 35388
rect 16148 35332 16152 35388
rect 16088 35328 16152 35332
rect 25778 35388 25842 35392
rect 25778 35332 25782 35388
rect 25782 35332 25838 35388
rect 25838 35332 25842 35388
rect 25778 35328 25842 35332
rect 25858 35388 25922 35392
rect 25858 35332 25862 35388
rect 25862 35332 25918 35388
rect 25918 35332 25922 35388
rect 25858 35328 25922 35332
rect 25938 35388 26002 35392
rect 25938 35332 25942 35388
rect 25942 35332 25998 35388
rect 25998 35332 26002 35388
rect 25938 35328 26002 35332
rect 26018 35388 26082 35392
rect 26018 35332 26022 35388
rect 26022 35332 26078 35388
rect 26078 35332 26082 35388
rect 26018 35328 26082 35332
rect 24164 35320 24228 35324
rect 24164 35264 24178 35320
rect 24178 35264 24228 35320
rect 24164 35260 24228 35264
rect 10882 34844 10946 34848
rect 10882 34788 10886 34844
rect 10886 34788 10942 34844
rect 10942 34788 10946 34844
rect 10882 34784 10946 34788
rect 10962 34844 11026 34848
rect 10962 34788 10966 34844
rect 10966 34788 11022 34844
rect 11022 34788 11026 34844
rect 10962 34784 11026 34788
rect 11042 34844 11106 34848
rect 11042 34788 11046 34844
rect 11046 34788 11102 34844
rect 11102 34788 11106 34844
rect 11042 34784 11106 34788
rect 11122 34844 11186 34848
rect 11122 34788 11126 34844
rect 11126 34788 11182 34844
rect 11182 34788 11186 34844
rect 11122 34784 11186 34788
rect 20813 34844 20877 34848
rect 20813 34788 20817 34844
rect 20817 34788 20873 34844
rect 20873 34788 20877 34844
rect 20813 34784 20877 34788
rect 20893 34844 20957 34848
rect 20893 34788 20897 34844
rect 20897 34788 20953 34844
rect 20953 34788 20957 34844
rect 20893 34784 20957 34788
rect 20973 34844 21037 34848
rect 20973 34788 20977 34844
rect 20977 34788 21033 34844
rect 21033 34788 21037 34844
rect 20973 34784 21037 34788
rect 21053 34844 21117 34848
rect 21053 34788 21057 34844
rect 21057 34788 21113 34844
rect 21113 34788 21117 34844
rect 21053 34784 21117 34788
rect 5917 34300 5981 34304
rect 5917 34244 5921 34300
rect 5921 34244 5977 34300
rect 5977 34244 5981 34300
rect 5917 34240 5981 34244
rect 5997 34300 6061 34304
rect 5997 34244 6001 34300
rect 6001 34244 6057 34300
rect 6057 34244 6061 34300
rect 5997 34240 6061 34244
rect 6077 34300 6141 34304
rect 6077 34244 6081 34300
rect 6081 34244 6137 34300
rect 6137 34244 6141 34300
rect 6077 34240 6141 34244
rect 6157 34300 6221 34304
rect 6157 34244 6161 34300
rect 6161 34244 6217 34300
rect 6217 34244 6221 34300
rect 6157 34240 6221 34244
rect 15848 34300 15912 34304
rect 15848 34244 15852 34300
rect 15852 34244 15908 34300
rect 15908 34244 15912 34300
rect 15848 34240 15912 34244
rect 15928 34300 15992 34304
rect 15928 34244 15932 34300
rect 15932 34244 15988 34300
rect 15988 34244 15992 34300
rect 15928 34240 15992 34244
rect 16008 34300 16072 34304
rect 16008 34244 16012 34300
rect 16012 34244 16068 34300
rect 16068 34244 16072 34300
rect 16008 34240 16072 34244
rect 16088 34300 16152 34304
rect 16088 34244 16092 34300
rect 16092 34244 16148 34300
rect 16148 34244 16152 34300
rect 16088 34240 16152 34244
rect 25778 34300 25842 34304
rect 25778 34244 25782 34300
rect 25782 34244 25838 34300
rect 25838 34244 25842 34300
rect 25778 34240 25842 34244
rect 25858 34300 25922 34304
rect 25858 34244 25862 34300
rect 25862 34244 25918 34300
rect 25918 34244 25922 34300
rect 25858 34240 25922 34244
rect 25938 34300 26002 34304
rect 25938 34244 25942 34300
rect 25942 34244 25998 34300
rect 25998 34244 26002 34300
rect 25938 34240 26002 34244
rect 26018 34300 26082 34304
rect 26018 34244 26022 34300
rect 26022 34244 26078 34300
rect 26078 34244 26082 34300
rect 26018 34240 26082 34244
rect 30236 34172 30300 34236
rect 17356 34036 17420 34100
rect 24348 33764 24412 33828
rect 10882 33756 10946 33760
rect 10882 33700 10886 33756
rect 10886 33700 10942 33756
rect 10942 33700 10946 33756
rect 10882 33696 10946 33700
rect 10962 33756 11026 33760
rect 10962 33700 10966 33756
rect 10966 33700 11022 33756
rect 11022 33700 11026 33756
rect 10962 33696 11026 33700
rect 11042 33756 11106 33760
rect 11042 33700 11046 33756
rect 11046 33700 11102 33756
rect 11102 33700 11106 33756
rect 11042 33696 11106 33700
rect 11122 33756 11186 33760
rect 11122 33700 11126 33756
rect 11126 33700 11182 33756
rect 11182 33700 11186 33756
rect 11122 33696 11186 33700
rect 20813 33756 20877 33760
rect 20813 33700 20817 33756
rect 20817 33700 20873 33756
rect 20873 33700 20877 33756
rect 20813 33696 20877 33700
rect 20893 33756 20957 33760
rect 20893 33700 20897 33756
rect 20897 33700 20953 33756
rect 20953 33700 20957 33756
rect 20893 33696 20957 33700
rect 20973 33756 21037 33760
rect 20973 33700 20977 33756
rect 20977 33700 21033 33756
rect 21033 33700 21037 33756
rect 20973 33696 21037 33700
rect 21053 33756 21117 33760
rect 21053 33700 21057 33756
rect 21057 33700 21113 33756
rect 21113 33700 21117 33756
rect 21053 33696 21117 33700
rect 27108 33552 27172 33556
rect 27108 33496 27158 33552
rect 27158 33496 27172 33552
rect 27108 33492 27172 33496
rect 5917 33212 5981 33216
rect 5917 33156 5921 33212
rect 5921 33156 5977 33212
rect 5977 33156 5981 33212
rect 5917 33152 5981 33156
rect 5997 33212 6061 33216
rect 5997 33156 6001 33212
rect 6001 33156 6057 33212
rect 6057 33156 6061 33212
rect 5997 33152 6061 33156
rect 6077 33212 6141 33216
rect 6077 33156 6081 33212
rect 6081 33156 6137 33212
rect 6137 33156 6141 33212
rect 6077 33152 6141 33156
rect 6157 33212 6221 33216
rect 6157 33156 6161 33212
rect 6161 33156 6217 33212
rect 6217 33156 6221 33212
rect 6157 33152 6221 33156
rect 15848 33212 15912 33216
rect 15848 33156 15852 33212
rect 15852 33156 15908 33212
rect 15908 33156 15912 33212
rect 15848 33152 15912 33156
rect 15928 33212 15992 33216
rect 15928 33156 15932 33212
rect 15932 33156 15988 33212
rect 15988 33156 15992 33212
rect 15928 33152 15992 33156
rect 16008 33212 16072 33216
rect 16008 33156 16012 33212
rect 16012 33156 16068 33212
rect 16068 33156 16072 33212
rect 16008 33152 16072 33156
rect 16088 33212 16152 33216
rect 16088 33156 16092 33212
rect 16092 33156 16148 33212
rect 16148 33156 16152 33212
rect 16088 33152 16152 33156
rect 25778 33212 25842 33216
rect 25778 33156 25782 33212
rect 25782 33156 25838 33212
rect 25838 33156 25842 33212
rect 25778 33152 25842 33156
rect 25858 33212 25922 33216
rect 25858 33156 25862 33212
rect 25862 33156 25918 33212
rect 25918 33156 25922 33212
rect 25858 33152 25922 33156
rect 25938 33212 26002 33216
rect 25938 33156 25942 33212
rect 25942 33156 25998 33212
rect 25998 33156 26002 33212
rect 25938 33152 26002 33156
rect 26018 33212 26082 33216
rect 26018 33156 26022 33212
rect 26022 33156 26078 33212
rect 26078 33156 26082 33212
rect 26018 33152 26082 33156
rect 25636 32948 25700 33012
rect 25636 32812 25700 32876
rect 29132 32812 29196 32876
rect 10882 32668 10946 32672
rect 10882 32612 10886 32668
rect 10886 32612 10942 32668
rect 10942 32612 10946 32668
rect 10882 32608 10946 32612
rect 10962 32668 11026 32672
rect 10962 32612 10966 32668
rect 10966 32612 11022 32668
rect 11022 32612 11026 32668
rect 10962 32608 11026 32612
rect 11042 32668 11106 32672
rect 11042 32612 11046 32668
rect 11046 32612 11102 32668
rect 11102 32612 11106 32668
rect 11042 32608 11106 32612
rect 11122 32668 11186 32672
rect 11122 32612 11126 32668
rect 11126 32612 11182 32668
rect 11182 32612 11186 32668
rect 11122 32608 11186 32612
rect 20813 32668 20877 32672
rect 20813 32612 20817 32668
rect 20817 32612 20873 32668
rect 20873 32612 20877 32668
rect 20813 32608 20877 32612
rect 20893 32668 20957 32672
rect 20893 32612 20897 32668
rect 20897 32612 20953 32668
rect 20953 32612 20957 32668
rect 20893 32608 20957 32612
rect 20973 32668 21037 32672
rect 20973 32612 20977 32668
rect 20977 32612 21033 32668
rect 21033 32612 21037 32668
rect 20973 32608 21037 32612
rect 21053 32668 21117 32672
rect 21053 32612 21057 32668
rect 21057 32612 21113 32668
rect 21113 32612 21117 32668
rect 21053 32608 21117 32612
rect 26188 32540 26252 32604
rect 26924 32540 26988 32604
rect 26924 32404 26988 32468
rect 29132 32676 29196 32740
rect 27292 32268 27356 32332
rect 23244 32192 23308 32196
rect 23244 32136 23258 32192
rect 23258 32136 23308 32192
rect 23244 32132 23308 32136
rect 26556 32132 26620 32196
rect 5917 32124 5981 32128
rect 5917 32068 5921 32124
rect 5921 32068 5977 32124
rect 5977 32068 5981 32124
rect 5917 32064 5981 32068
rect 5997 32124 6061 32128
rect 5997 32068 6001 32124
rect 6001 32068 6057 32124
rect 6057 32068 6061 32124
rect 5997 32064 6061 32068
rect 6077 32124 6141 32128
rect 6077 32068 6081 32124
rect 6081 32068 6137 32124
rect 6137 32068 6141 32124
rect 6077 32064 6141 32068
rect 6157 32124 6221 32128
rect 6157 32068 6161 32124
rect 6161 32068 6217 32124
rect 6217 32068 6221 32124
rect 6157 32064 6221 32068
rect 15848 32124 15912 32128
rect 15848 32068 15852 32124
rect 15852 32068 15908 32124
rect 15908 32068 15912 32124
rect 15848 32064 15912 32068
rect 15928 32124 15992 32128
rect 15928 32068 15932 32124
rect 15932 32068 15988 32124
rect 15988 32068 15992 32124
rect 15928 32064 15992 32068
rect 16008 32124 16072 32128
rect 16008 32068 16012 32124
rect 16012 32068 16068 32124
rect 16068 32068 16072 32124
rect 16008 32064 16072 32068
rect 16088 32124 16152 32128
rect 16088 32068 16092 32124
rect 16092 32068 16148 32124
rect 16148 32068 16152 32124
rect 16088 32064 16152 32068
rect 25778 32124 25842 32128
rect 25778 32068 25782 32124
rect 25782 32068 25838 32124
rect 25838 32068 25842 32124
rect 25778 32064 25842 32068
rect 25858 32124 25922 32128
rect 25858 32068 25862 32124
rect 25862 32068 25918 32124
rect 25918 32068 25922 32124
rect 25858 32064 25922 32068
rect 25938 32124 26002 32128
rect 25938 32068 25942 32124
rect 25942 32068 25998 32124
rect 25998 32068 26002 32124
rect 25938 32064 26002 32068
rect 26018 32124 26082 32128
rect 26018 32068 26022 32124
rect 26022 32068 26078 32124
rect 26078 32068 26082 32124
rect 26018 32064 26082 32068
rect 24716 31996 24780 32060
rect 25268 31724 25332 31788
rect 27108 31724 27172 31788
rect 27660 32132 27724 32196
rect 27660 32056 27724 32060
rect 30972 32268 31036 32332
rect 27660 32000 27710 32056
rect 27710 32000 27724 32056
rect 27660 31996 27724 32000
rect 28212 31860 28276 31924
rect 30420 31860 30484 31924
rect 30604 31724 30668 31788
rect 10882 31580 10946 31584
rect 10882 31524 10886 31580
rect 10886 31524 10942 31580
rect 10942 31524 10946 31580
rect 10882 31520 10946 31524
rect 10962 31580 11026 31584
rect 10962 31524 10966 31580
rect 10966 31524 11022 31580
rect 11022 31524 11026 31580
rect 10962 31520 11026 31524
rect 11042 31580 11106 31584
rect 11042 31524 11046 31580
rect 11046 31524 11102 31580
rect 11102 31524 11106 31580
rect 11042 31520 11106 31524
rect 11122 31580 11186 31584
rect 11122 31524 11126 31580
rect 11126 31524 11182 31580
rect 11182 31524 11186 31580
rect 11122 31520 11186 31524
rect 20813 31580 20877 31584
rect 20813 31524 20817 31580
rect 20817 31524 20873 31580
rect 20873 31524 20877 31580
rect 20813 31520 20877 31524
rect 20893 31580 20957 31584
rect 20893 31524 20897 31580
rect 20897 31524 20953 31580
rect 20953 31524 20957 31580
rect 20893 31520 20957 31524
rect 20973 31580 21037 31584
rect 20973 31524 20977 31580
rect 20977 31524 21033 31580
rect 21033 31524 21037 31580
rect 20973 31520 21037 31524
rect 21053 31580 21117 31584
rect 21053 31524 21057 31580
rect 21057 31524 21113 31580
rect 21113 31524 21117 31580
rect 21053 31520 21117 31524
rect 26372 31588 26436 31652
rect 31156 31860 31220 31924
rect 23244 31512 23308 31516
rect 23244 31456 23294 31512
rect 23294 31456 23308 31512
rect 23244 31452 23308 31456
rect 27660 31452 27724 31516
rect 25084 31316 25148 31380
rect 27660 31316 27724 31380
rect 30420 31316 30484 31380
rect 25452 31180 25516 31244
rect 5917 31036 5981 31040
rect 5917 30980 5921 31036
rect 5921 30980 5977 31036
rect 5977 30980 5981 31036
rect 5917 30976 5981 30980
rect 5997 31036 6061 31040
rect 5997 30980 6001 31036
rect 6001 30980 6057 31036
rect 6057 30980 6061 31036
rect 5997 30976 6061 30980
rect 6077 31036 6141 31040
rect 6077 30980 6081 31036
rect 6081 30980 6137 31036
rect 6137 30980 6141 31036
rect 6077 30976 6141 30980
rect 6157 31036 6221 31040
rect 6157 30980 6161 31036
rect 6161 30980 6217 31036
rect 6217 30980 6221 31036
rect 6157 30976 6221 30980
rect 15848 31036 15912 31040
rect 15848 30980 15852 31036
rect 15852 30980 15908 31036
rect 15908 30980 15912 31036
rect 15848 30976 15912 30980
rect 15928 31036 15992 31040
rect 15928 30980 15932 31036
rect 15932 30980 15988 31036
rect 15988 30980 15992 31036
rect 15928 30976 15992 30980
rect 16008 31036 16072 31040
rect 16008 30980 16012 31036
rect 16012 30980 16068 31036
rect 16068 30980 16072 31036
rect 16008 30976 16072 30980
rect 16088 31036 16152 31040
rect 16088 30980 16092 31036
rect 16092 30980 16148 31036
rect 16148 30980 16152 31036
rect 16088 30976 16152 30980
rect 25778 31036 25842 31040
rect 25778 30980 25782 31036
rect 25782 30980 25838 31036
rect 25838 30980 25842 31036
rect 25778 30976 25842 30980
rect 25858 31036 25922 31040
rect 25858 30980 25862 31036
rect 25862 30980 25918 31036
rect 25918 30980 25922 31036
rect 25858 30976 25922 30980
rect 25938 31036 26002 31040
rect 25938 30980 25942 31036
rect 25942 30980 25998 31036
rect 25998 30980 26002 31036
rect 25938 30976 26002 30980
rect 26018 31036 26082 31040
rect 26018 30980 26022 31036
rect 26022 30980 26078 31036
rect 26078 30980 26082 31036
rect 26018 30976 26082 30980
rect 27476 31044 27540 31108
rect 30604 31044 30668 31108
rect 27476 30968 27540 30972
rect 27476 30912 27526 30968
rect 27526 30912 27540 30968
rect 27476 30908 27540 30912
rect 28948 30908 29012 30972
rect 31156 30908 31220 30972
rect 28948 30772 29012 30836
rect 25268 30636 25332 30700
rect 10882 30492 10946 30496
rect 10882 30436 10886 30492
rect 10886 30436 10942 30492
rect 10942 30436 10946 30492
rect 10882 30432 10946 30436
rect 10962 30492 11026 30496
rect 10962 30436 10966 30492
rect 10966 30436 11022 30492
rect 11022 30436 11026 30492
rect 10962 30432 11026 30436
rect 11042 30492 11106 30496
rect 11042 30436 11046 30492
rect 11046 30436 11102 30492
rect 11102 30436 11106 30492
rect 11042 30432 11106 30436
rect 11122 30492 11186 30496
rect 11122 30436 11126 30492
rect 11126 30436 11182 30492
rect 11182 30436 11186 30492
rect 11122 30432 11186 30436
rect 20813 30492 20877 30496
rect 20813 30436 20817 30492
rect 20817 30436 20873 30492
rect 20873 30436 20877 30492
rect 20813 30432 20877 30436
rect 20893 30492 20957 30496
rect 20893 30436 20897 30492
rect 20897 30436 20953 30492
rect 20953 30436 20957 30492
rect 20893 30432 20957 30436
rect 20973 30492 21037 30496
rect 20973 30436 20977 30492
rect 20977 30436 21033 30492
rect 21033 30436 21037 30492
rect 20973 30432 21037 30436
rect 21053 30492 21117 30496
rect 21053 30436 21057 30492
rect 21057 30436 21113 30492
rect 21113 30436 21117 30492
rect 21053 30432 21117 30436
rect 26372 30364 26436 30428
rect 30788 30364 30852 30428
rect 24164 30228 24228 30292
rect 25268 30092 25332 30156
rect 26188 30092 26252 30156
rect 5917 29948 5981 29952
rect 5917 29892 5921 29948
rect 5921 29892 5977 29948
rect 5977 29892 5981 29948
rect 5917 29888 5981 29892
rect 5997 29948 6061 29952
rect 5997 29892 6001 29948
rect 6001 29892 6057 29948
rect 6057 29892 6061 29948
rect 5997 29888 6061 29892
rect 6077 29948 6141 29952
rect 6077 29892 6081 29948
rect 6081 29892 6137 29948
rect 6137 29892 6141 29948
rect 6077 29888 6141 29892
rect 6157 29948 6221 29952
rect 6157 29892 6161 29948
rect 6161 29892 6217 29948
rect 6217 29892 6221 29948
rect 6157 29888 6221 29892
rect 15848 29948 15912 29952
rect 15848 29892 15852 29948
rect 15852 29892 15908 29948
rect 15908 29892 15912 29948
rect 15848 29888 15912 29892
rect 15928 29948 15992 29952
rect 15928 29892 15932 29948
rect 15932 29892 15988 29948
rect 15988 29892 15992 29948
rect 15928 29888 15992 29892
rect 16008 29948 16072 29952
rect 16008 29892 16012 29948
rect 16012 29892 16068 29948
rect 16068 29892 16072 29948
rect 16008 29888 16072 29892
rect 16088 29948 16152 29952
rect 16088 29892 16092 29948
rect 16092 29892 16148 29948
rect 16148 29892 16152 29948
rect 16088 29888 16152 29892
rect 25778 29948 25842 29952
rect 25778 29892 25782 29948
rect 25782 29892 25838 29948
rect 25838 29892 25842 29948
rect 25778 29888 25842 29892
rect 25858 29948 25922 29952
rect 25858 29892 25862 29948
rect 25862 29892 25918 29948
rect 25918 29892 25922 29948
rect 25858 29888 25922 29892
rect 25938 29948 26002 29952
rect 25938 29892 25942 29948
rect 25942 29892 25998 29948
rect 25998 29892 26002 29948
rect 25938 29888 26002 29892
rect 26018 29948 26082 29952
rect 26018 29892 26022 29948
rect 26022 29892 26078 29948
rect 26078 29892 26082 29948
rect 26018 29888 26082 29892
rect 22140 29880 22204 29884
rect 22140 29824 22154 29880
rect 22154 29824 22204 29880
rect 22140 29820 22204 29824
rect 27108 29880 27172 29884
rect 27108 29824 27122 29880
rect 27122 29824 27172 29880
rect 27108 29820 27172 29824
rect 24900 29684 24964 29748
rect 26740 29744 26804 29748
rect 26740 29688 26790 29744
rect 26790 29688 26804 29744
rect 26740 29684 26804 29688
rect 26740 29548 26804 29612
rect 30604 29956 30668 30020
rect 28212 29820 28276 29884
rect 10882 29404 10946 29408
rect 10882 29348 10886 29404
rect 10886 29348 10942 29404
rect 10942 29348 10946 29404
rect 10882 29344 10946 29348
rect 10962 29404 11026 29408
rect 10962 29348 10966 29404
rect 10966 29348 11022 29404
rect 11022 29348 11026 29404
rect 10962 29344 11026 29348
rect 11042 29404 11106 29408
rect 11042 29348 11046 29404
rect 11046 29348 11102 29404
rect 11102 29348 11106 29404
rect 11042 29344 11106 29348
rect 11122 29404 11186 29408
rect 11122 29348 11126 29404
rect 11126 29348 11182 29404
rect 11182 29348 11186 29404
rect 11122 29344 11186 29348
rect 20813 29404 20877 29408
rect 20813 29348 20817 29404
rect 20817 29348 20873 29404
rect 20873 29348 20877 29404
rect 20813 29344 20877 29348
rect 20893 29404 20957 29408
rect 20893 29348 20897 29404
rect 20897 29348 20953 29404
rect 20953 29348 20957 29404
rect 20893 29344 20957 29348
rect 20973 29404 21037 29408
rect 20973 29348 20977 29404
rect 20977 29348 21033 29404
rect 21033 29348 21037 29404
rect 20973 29344 21037 29348
rect 21053 29404 21117 29408
rect 21053 29348 21057 29404
rect 21057 29348 21113 29404
rect 21113 29348 21117 29404
rect 21053 29344 21117 29348
rect 26188 29276 26252 29340
rect 27292 29140 27356 29204
rect 28028 28868 28092 28932
rect 5917 28860 5981 28864
rect 5917 28804 5921 28860
rect 5921 28804 5977 28860
rect 5977 28804 5981 28860
rect 5917 28800 5981 28804
rect 5997 28860 6061 28864
rect 5997 28804 6001 28860
rect 6001 28804 6057 28860
rect 6057 28804 6061 28860
rect 5997 28800 6061 28804
rect 6077 28860 6141 28864
rect 6077 28804 6081 28860
rect 6081 28804 6137 28860
rect 6137 28804 6141 28860
rect 6077 28800 6141 28804
rect 6157 28860 6221 28864
rect 6157 28804 6161 28860
rect 6161 28804 6217 28860
rect 6217 28804 6221 28860
rect 6157 28800 6221 28804
rect 15848 28860 15912 28864
rect 15848 28804 15852 28860
rect 15852 28804 15908 28860
rect 15908 28804 15912 28860
rect 15848 28800 15912 28804
rect 15928 28860 15992 28864
rect 15928 28804 15932 28860
rect 15932 28804 15988 28860
rect 15988 28804 15992 28860
rect 15928 28800 15992 28804
rect 16008 28860 16072 28864
rect 16008 28804 16012 28860
rect 16012 28804 16068 28860
rect 16068 28804 16072 28860
rect 16008 28800 16072 28804
rect 16088 28860 16152 28864
rect 16088 28804 16092 28860
rect 16092 28804 16148 28860
rect 16148 28804 16152 28860
rect 16088 28800 16152 28804
rect 25778 28860 25842 28864
rect 25778 28804 25782 28860
rect 25782 28804 25838 28860
rect 25838 28804 25842 28860
rect 25778 28800 25842 28804
rect 25858 28860 25922 28864
rect 25858 28804 25862 28860
rect 25862 28804 25918 28860
rect 25918 28804 25922 28860
rect 25858 28800 25922 28804
rect 25938 28860 26002 28864
rect 25938 28804 25942 28860
rect 25942 28804 25998 28860
rect 25998 28804 26002 28860
rect 25938 28800 26002 28804
rect 26018 28860 26082 28864
rect 26018 28804 26022 28860
rect 26022 28804 26078 28860
rect 26078 28804 26082 28860
rect 26018 28800 26082 28804
rect 30604 28732 30668 28796
rect 25084 28656 25148 28660
rect 25084 28600 25098 28656
rect 25098 28600 25148 28656
rect 25084 28596 25148 28600
rect 10882 28316 10946 28320
rect 10882 28260 10886 28316
rect 10886 28260 10942 28316
rect 10942 28260 10946 28316
rect 10882 28256 10946 28260
rect 10962 28316 11026 28320
rect 10962 28260 10966 28316
rect 10966 28260 11022 28316
rect 11022 28260 11026 28316
rect 10962 28256 11026 28260
rect 11042 28316 11106 28320
rect 11042 28260 11046 28316
rect 11046 28260 11102 28316
rect 11102 28260 11106 28316
rect 11042 28256 11106 28260
rect 11122 28316 11186 28320
rect 11122 28260 11126 28316
rect 11126 28260 11182 28316
rect 11182 28260 11186 28316
rect 11122 28256 11186 28260
rect 20813 28316 20877 28320
rect 20813 28260 20817 28316
rect 20817 28260 20873 28316
rect 20873 28260 20877 28316
rect 20813 28256 20877 28260
rect 20893 28316 20957 28320
rect 20893 28260 20897 28316
rect 20897 28260 20953 28316
rect 20953 28260 20957 28316
rect 20893 28256 20957 28260
rect 20973 28316 21037 28320
rect 20973 28260 20977 28316
rect 20977 28260 21033 28316
rect 21033 28260 21037 28316
rect 20973 28256 21037 28260
rect 21053 28316 21117 28320
rect 21053 28260 21057 28316
rect 21057 28260 21113 28316
rect 21113 28260 21117 28316
rect 21053 28256 21117 28260
rect 15516 28188 15580 28252
rect 5917 27772 5981 27776
rect 5917 27716 5921 27772
rect 5921 27716 5977 27772
rect 5977 27716 5981 27772
rect 5917 27712 5981 27716
rect 5997 27772 6061 27776
rect 5997 27716 6001 27772
rect 6001 27716 6057 27772
rect 6057 27716 6061 27772
rect 5997 27712 6061 27716
rect 6077 27772 6141 27776
rect 6077 27716 6081 27772
rect 6081 27716 6137 27772
rect 6137 27716 6141 27772
rect 6077 27712 6141 27716
rect 6157 27772 6221 27776
rect 6157 27716 6161 27772
rect 6161 27716 6217 27772
rect 6217 27716 6221 27772
rect 6157 27712 6221 27716
rect 19196 28052 19260 28116
rect 25452 27916 25516 27980
rect 26372 27916 26436 27980
rect 15516 27840 15580 27844
rect 15516 27784 15530 27840
rect 15530 27784 15580 27840
rect 15516 27780 15580 27784
rect 29132 27780 29196 27844
rect 15848 27772 15912 27776
rect 15848 27716 15852 27772
rect 15852 27716 15908 27772
rect 15908 27716 15912 27772
rect 15848 27712 15912 27716
rect 15928 27772 15992 27776
rect 15928 27716 15932 27772
rect 15932 27716 15988 27772
rect 15988 27716 15992 27772
rect 15928 27712 15992 27716
rect 16008 27772 16072 27776
rect 16008 27716 16012 27772
rect 16012 27716 16068 27772
rect 16068 27716 16072 27772
rect 16008 27712 16072 27716
rect 16088 27772 16152 27776
rect 16088 27716 16092 27772
rect 16092 27716 16148 27772
rect 16148 27716 16152 27772
rect 16088 27712 16152 27716
rect 25778 27772 25842 27776
rect 25778 27716 25782 27772
rect 25782 27716 25838 27772
rect 25838 27716 25842 27772
rect 25778 27712 25842 27716
rect 25858 27772 25922 27776
rect 25858 27716 25862 27772
rect 25862 27716 25918 27772
rect 25918 27716 25922 27772
rect 25858 27712 25922 27716
rect 25938 27772 26002 27776
rect 25938 27716 25942 27772
rect 25942 27716 25998 27772
rect 25998 27716 26002 27772
rect 25938 27712 26002 27716
rect 26018 27772 26082 27776
rect 26018 27716 26022 27772
rect 26022 27716 26078 27772
rect 26078 27716 26082 27772
rect 26018 27712 26082 27716
rect 17540 27508 17604 27572
rect 26924 27372 26988 27436
rect 26372 27236 26436 27300
rect 10882 27228 10946 27232
rect 10882 27172 10886 27228
rect 10886 27172 10942 27228
rect 10942 27172 10946 27228
rect 10882 27168 10946 27172
rect 10962 27228 11026 27232
rect 10962 27172 10966 27228
rect 10966 27172 11022 27228
rect 11022 27172 11026 27228
rect 10962 27168 11026 27172
rect 11042 27228 11106 27232
rect 11042 27172 11046 27228
rect 11046 27172 11102 27228
rect 11102 27172 11106 27228
rect 11042 27168 11106 27172
rect 11122 27228 11186 27232
rect 11122 27172 11126 27228
rect 11126 27172 11182 27228
rect 11182 27172 11186 27228
rect 11122 27168 11186 27172
rect 20813 27228 20877 27232
rect 20813 27172 20817 27228
rect 20817 27172 20873 27228
rect 20873 27172 20877 27228
rect 20813 27168 20877 27172
rect 20893 27228 20957 27232
rect 20893 27172 20897 27228
rect 20897 27172 20953 27228
rect 20953 27172 20957 27228
rect 20893 27168 20957 27172
rect 20973 27228 21037 27232
rect 20973 27172 20977 27228
rect 20977 27172 21033 27228
rect 21033 27172 21037 27228
rect 20973 27168 21037 27172
rect 21053 27228 21117 27232
rect 21053 27172 21057 27228
rect 21057 27172 21113 27228
rect 21113 27172 21117 27228
rect 21053 27168 21117 27172
rect 25452 27160 25516 27164
rect 25452 27104 25466 27160
rect 25466 27104 25516 27160
rect 25452 27100 25516 27104
rect 27292 26964 27356 27028
rect 25636 26828 25700 26892
rect 28028 26692 28092 26756
rect 5917 26684 5981 26688
rect 5917 26628 5921 26684
rect 5921 26628 5977 26684
rect 5977 26628 5981 26684
rect 5917 26624 5981 26628
rect 5997 26684 6061 26688
rect 5997 26628 6001 26684
rect 6001 26628 6057 26684
rect 6057 26628 6061 26684
rect 5997 26624 6061 26628
rect 6077 26684 6141 26688
rect 6077 26628 6081 26684
rect 6081 26628 6137 26684
rect 6137 26628 6141 26684
rect 6077 26624 6141 26628
rect 6157 26684 6221 26688
rect 6157 26628 6161 26684
rect 6161 26628 6217 26684
rect 6217 26628 6221 26684
rect 6157 26624 6221 26628
rect 15848 26684 15912 26688
rect 15848 26628 15852 26684
rect 15852 26628 15908 26684
rect 15908 26628 15912 26684
rect 15848 26624 15912 26628
rect 15928 26684 15992 26688
rect 15928 26628 15932 26684
rect 15932 26628 15988 26684
rect 15988 26628 15992 26684
rect 15928 26624 15992 26628
rect 16008 26684 16072 26688
rect 16008 26628 16012 26684
rect 16012 26628 16068 26684
rect 16068 26628 16072 26684
rect 16008 26624 16072 26628
rect 16088 26684 16152 26688
rect 16088 26628 16092 26684
rect 16092 26628 16148 26684
rect 16148 26628 16152 26684
rect 16088 26624 16152 26628
rect 25778 26684 25842 26688
rect 25778 26628 25782 26684
rect 25782 26628 25838 26684
rect 25838 26628 25842 26684
rect 25778 26624 25842 26628
rect 25858 26684 25922 26688
rect 25858 26628 25862 26684
rect 25862 26628 25918 26684
rect 25918 26628 25922 26684
rect 25858 26624 25922 26628
rect 25938 26684 26002 26688
rect 25938 26628 25942 26684
rect 25942 26628 25998 26684
rect 25998 26628 26002 26684
rect 25938 26624 26002 26628
rect 26018 26684 26082 26688
rect 26018 26628 26022 26684
rect 26022 26628 26078 26684
rect 26078 26628 26082 26684
rect 26018 26624 26082 26628
rect 27660 26556 27724 26620
rect 10882 26140 10946 26144
rect 10882 26084 10886 26140
rect 10886 26084 10942 26140
rect 10942 26084 10946 26140
rect 10882 26080 10946 26084
rect 10962 26140 11026 26144
rect 10962 26084 10966 26140
rect 10966 26084 11022 26140
rect 11022 26084 11026 26140
rect 10962 26080 11026 26084
rect 11042 26140 11106 26144
rect 11042 26084 11046 26140
rect 11046 26084 11102 26140
rect 11102 26084 11106 26140
rect 11042 26080 11106 26084
rect 11122 26140 11186 26144
rect 11122 26084 11126 26140
rect 11126 26084 11182 26140
rect 11182 26084 11186 26140
rect 11122 26080 11186 26084
rect 20813 26140 20877 26144
rect 20813 26084 20817 26140
rect 20817 26084 20873 26140
rect 20873 26084 20877 26140
rect 20813 26080 20877 26084
rect 20893 26140 20957 26144
rect 20893 26084 20897 26140
rect 20897 26084 20953 26140
rect 20953 26084 20957 26140
rect 20893 26080 20957 26084
rect 20973 26140 21037 26144
rect 20973 26084 20977 26140
rect 20977 26084 21033 26140
rect 21033 26084 21037 26140
rect 20973 26080 21037 26084
rect 21053 26140 21117 26144
rect 21053 26084 21057 26140
rect 21057 26084 21113 26140
rect 21113 26084 21117 26140
rect 21053 26080 21117 26084
rect 28212 25876 28276 25940
rect 28948 25936 29012 25940
rect 28948 25880 28962 25936
rect 28962 25880 29012 25936
rect 28948 25876 29012 25880
rect 26556 25740 26620 25804
rect 5917 25596 5981 25600
rect 5917 25540 5921 25596
rect 5921 25540 5977 25596
rect 5977 25540 5981 25596
rect 5917 25536 5981 25540
rect 5997 25596 6061 25600
rect 5997 25540 6001 25596
rect 6001 25540 6057 25596
rect 6057 25540 6061 25596
rect 5997 25536 6061 25540
rect 6077 25596 6141 25600
rect 6077 25540 6081 25596
rect 6081 25540 6137 25596
rect 6137 25540 6141 25596
rect 6077 25536 6141 25540
rect 6157 25596 6221 25600
rect 6157 25540 6161 25596
rect 6161 25540 6217 25596
rect 6217 25540 6221 25596
rect 6157 25536 6221 25540
rect 15848 25596 15912 25600
rect 15848 25540 15852 25596
rect 15852 25540 15908 25596
rect 15908 25540 15912 25596
rect 15848 25536 15912 25540
rect 15928 25596 15992 25600
rect 15928 25540 15932 25596
rect 15932 25540 15988 25596
rect 15988 25540 15992 25596
rect 15928 25536 15992 25540
rect 16008 25596 16072 25600
rect 16008 25540 16012 25596
rect 16012 25540 16068 25596
rect 16068 25540 16072 25596
rect 16008 25536 16072 25540
rect 16088 25596 16152 25600
rect 16088 25540 16092 25596
rect 16092 25540 16148 25596
rect 16148 25540 16152 25596
rect 16088 25536 16152 25540
rect 25778 25596 25842 25600
rect 25778 25540 25782 25596
rect 25782 25540 25838 25596
rect 25838 25540 25842 25596
rect 25778 25536 25842 25540
rect 25858 25596 25922 25600
rect 25858 25540 25862 25596
rect 25862 25540 25918 25596
rect 25918 25540 25922 25596
rect 25858 25536 25922 25540
rect 25938 25596 26002 25600
rect 25938 25540 25942 25596
rect 25942 25540 25998 25596
rect 25998 25540 26002 25596
rect 25938 25536 26002 25540
rect 26018 25596 26082 25600
rect 26018 25540 26022 25596
rect 26022 25540 26078 25596
rect 26078 25540 26082 25596
rect 26018 25536 26082 25540
rect 24900 25392 24964 25396
rect 24900 25336 24914 25392
rect 24914 25336 24964 25392
rect 24900 25332 24964 25336
rect 25268 25256 25332 25260
rect 25268 25200 25318 25256
rect 25318 25200 25332 25256
rect 25268 25196 25332 25200
rect 10882 25052 10946 25056
rect 10882 24996 10886 25052
rect 10886 24996 10942 25052
rect 10942 24996 10946 25052
rect 10882 24992 10946 24996
rect 10962 25052 11026 25056
rect 10962 24996 10966 25052
rect 10966 24996 11022 25052
rect 11022 24996 11026 25052
rect 10962 24992 11026 24996
rect 11042 25052 11106 25056
rect 11042 24996 11046 25052
rect 11046 24996 11102 25052
rect 11102 24996 11106 25052
rect 11042 24992 11106 24996
rect 11122 25052 11186 25056
rect 11122 24996 11126 25052
rect 11126 24996 11182 25052
rect 11182 24996 11186 25052
rect 11122 24992 11186 24996
rect 20813 25052 20877 25056
rect 20813 24996 20817 25052
rect 20817 24996 20873 25052
rect 20873 24996 20877 25052
rect 20813 24992 20877 24996
rect 20893 25052 20957 25056
rect 20893 24996 20897 25052
rect 20897 24996 20953 25052
rect 20953 24996 20957 25052
rect 20893 24992 20957 24996
rect 20973 25052 21037 25056
rect 20973 24996 20977 25052
rect 20977 24996 21033 25052
rect 21033 24996 21037 25052
rect 20973 24992 21037 24996
rect 21053 25052 21117 25056
rect 21053 24996 21057 25052
rect 21057 24996 21113 25052
rect 21113 24996 21117 25052
rect 21053 24992 21117 24996
rect 27292 25196 27356 25260
rect 22140 24788 22204 24852
rect 30236 24788 30300 24852
rect 26188 24712 26252 24716
rect 26188 24656 26238 24712
rect 26238 24656 26252 24712
rect 26188 24652 26252 24656
rect 5917 24508 5981 24512
rect 5917 24452 5921 24508
rect 5921 24452 5977 24508
rect 5977 24452 5981 24508
rect 5917 24448 5981 24452
rect 5997 24508 6061 24512
rect 5997 24452 6001 24508
rect 6001 24452 6057 24508
rect 6057 24452 6061 24508
rect 5997 24448 6061 24452
rect 6077 24508 6141 24512
rect 6077 24452 6081 24508
rect 6081 24452 6137 24508
rect 6137 24452 6141 24508
rect 6077 24448 6141 24452
rect 6157 24508 6221 24512
rect 6157 24452 6161 24508
rect 6161 24452 6217 24508
rect 6217 24452 6221 24508
rect 6157 24448 6221 24452
rect 15848 24508 15912 24512
rect 15848 24452 15852 24508
rect 15852 24452 15908 24508
rect 15908 24452 15912 24508
rect 15848 24448 15912 24452
rect 15928 24508 15992 24512
rect 15928 24452 15932 24508
rect 15932 24452 15988 24508
rect 15988 24452 15992 24508
rect 15928 24448 15992 24452
rect 16008 24508 16072 24512
rect 16008 24452 16012 24508
rect 16012 24452 16068 24508
rect 16068 24452 16072 24508
rect 16008 24448 16072 24452
rect 16088 24508 16152 24512
rect 16088 24452 16092 24508
rect 16092 24452 16148 24508
rect 16148 24452 16152 24508
rect 16088 24448 16152 24452
rect 25778 24508 25842 24512
rect 25778 24452 25782 24508
rect 25782 24452 25838 24508
rect 25838 24452 25842 24508
rect 25778 24448 25842 24452
rect 25858 24508 25922 24512
rect 25858 24452 25862 24508
rect 25862 24452 25918 24508
rect 25918 24452 25922 24508
rect 25858 24448 25922 24452
rect 25938 24508 26002 24512
rect 25938 24452 25942 24508
rect 25942 24452 25998 24508
rect 25998 24452 26002 24508
rect 25938 24448 26002 24452
rect 26018 24508 26082 24512
rect 26018 24452 26022 24508
rect 26022 24452 26078 24508
rect 26078 24452 26082 24508
rect 26018 24448 26082 24452
rect 25268 24108 25332 24172
rect 26740 23972 26804 24036
rect 10882 23964 10946 23968
rect 10882 23908 10886 23964
rect 10886 23908 10942 23964
rect 10942 23908 10946 23964
rect 10882 23904 10946 23908
rect 10962 23964 11026 23968
rect 10962 23908 10966 23964
rect 10966 23908 11022 23964
rect 11022 23908 11026 23964
rect 10962 23904 11026 23908
rect 11042 23964 11106 23968
rect 11042 23908 11046 23964
rect 11046 23908 11102 23964
rect 11102 23908 11106 23964
rect 11042 23904 11106 23908
rect 11122 23964 11186 23968
rect 11122 23908 11126 23964
rect 11126 23908 11182 23964
rect 11182 23908 11186 23964
rect 11122 23904 11186 23908
rect 20813 23964 20877 23968
rect 20813 23908 20817 23964
rect 20817 23908 20873 23964
rect 20873 23908 20877 23964
rect 20813 23904 20877 23908
rect 20893 23964 20957 23968
rect 20893 23908 20897 23964
rect 20897 23908 20953 23964
rect 20953 23908 20957 23964
rect 20893 23904 20957 23908
rect 20973 23964 21037 23968
rect 20973 23908 20977 23964
rect 20977 23908 21033 23964
rect 21033 23908 21037 23964
rect 20973 23904 21037 23908
rect 21053 23964 21117 23968
rect 21053 23908 21057 23964
rect 21057 23908 21113 23964
rect 21113 23908 21117 23964
rect 21053 23904 21117 23908
rect 27476 23836 27540 23900
rect 28028 23700 28092 23764
rect 5917 23420 5981 23424
rect 5917 23364 5921 23420
rect 5921 23364 5977 23420
rect 5977 23364 5981 23420
rect 5917 23360 5981 23364
rect 5997 23420 6061 23424
rect 5997 23364 6001 23420
rect 6001 23364 6057 23420
rect 6057 23364 6061 23420
rect 5997 23360 6061 23364
rect 6077 23420 6141 23424
rect 6077 23364 6081 23420
rect 6081 23364 6137 23420
rect 6137 23364 6141 23420
rect 6077 23360 6141 23364
rect 6157 23420 6221 23424
rect 6157 23364 6161 23420
rect 6161 23364 6217 23420
rect 6217 23364 6221 23420
rect 6157 23360 6221 23364
rect 15848 23420 15912 23424
rect 15848 23364 15852 23420
rect 15852 23364 15908 23420
rect 15908 23364 15912 23420
rect 15848 23360 15912 23364
rect 15928 23420 15992 23424
rect 15928 23364 15932 23420
rect 15932 23364 15988 23420
rect 15988 23364 15992 23420
rect 15928 23360 15992 23364
rect 16008 23420 16072 23424
rect 16008 23364 16012 23420
rect 16012 23364 16068 23420
rect 16068 23364 16072 23420
rect 16008 23360 16072 23364
rect 16088 23420 16152 23424
rect 16088 23364 16092 23420
rect 16092 23364 16148 23420
rect 16148 23364 16152 23420
rect 16088 23360 16152 23364
rect 25778 23420 25842 23424
rect 25778 23364 25782 23420
rect 25782 23364 25838 23420
rect 25838 23364 25842 23420
rect 25778 23360 25842 23364
rect 25858 23420 25922 23424
rect 25858 23364 25862 23420
rect 25862 23364 25918 23420
rect 25918 23364 25922 23420
rect 25858 23360 25922 23364
rect 25938 23420 26002 23424
rect 25938 23364 25942 23420
rect 25942 23364 25998 23420
rect 25998 23364 26002 23420
rect 25938 23360 26002 23364
rect 26018 23420 26082 23424
rect 26018 23364 26022 23420
rect 26022 23364 26078 23420
rect 26078 23364 26082 23420
rect 26018 23360 26082 23364
rect 10882 22876 10946 22880
rect 10882 22820 10886 22876
rect 10886 22820 10942 22876
rect 10942 22820 10946 22876
rect 10882 22816 10946 22820
rect 10962 22876 11026 22880
rect 10962 22820 10966 22876
rect 10966 22820 11022 22876
rect 11022 22820 11026 22876
rect 10962 22816 11026 22820
rect 11042 22876 11106 22880
rect 11042 22820 11046 22876
rect 11046 22820 11102 22876
rect 11102 22820 11106 22876
rect 11042 22816 11106 22820
rect 11122 22876 11186 22880
rect 11122 22820 11126 22876
rect 11126 22820 11182 22876
rect 11182 22820 11186 22876
rect 11122 22816 11186 22820
rect 20813 22876 20877 22880
rect 20813 22820 20817 22876
rect 20817 22820 20873 22876
rect 20873 22820 20877 22876
rect 20813 22816 20877 22820
rect 20893 22876 20957 22880
rect 20893 22820 20897 22876
rect 20897 22820 20953 22876
rect 20953 22820 20957 22876
rect 20893 22816 20957 22820
rect 20973 22876 21037 22880
rect 20973 22820 20977 22876
rect 20977 22820 21033 22876
rect 21033 22820 21037 22876
rect 20973 22816 21037 22820
rect 21053 22876 21117 22880
rect 21053 22820 21057 22876
rect 21057 22820 21113 22876
rect 21113 22820 21117 22876
rect 21053 22816 21117 22820
rect 24900 23020 24964 23084
rect 24716 22748 24780 22812
rect 26188 22748 26252 22812
rect 25636 22340 25700 22404
rect 5917 22332 5981 22336
rect 5917 22276 5921 22332
rect 5921 22276 5977 22332
rect 5977 22276 5981 22332
rect 5917 22272 5981 22276
rect 5997 22332 6061 22336
rect 5997 22276 6001 22332
rect 6001 22276 6057 22332
rect 6057 22276 6061 22332
rect 5997 22272 6061 22276
rect 6077 22332 6141 22336
rect 6077 22276 6081 22332
rect 6081 22276 6137 22332
rect 6137 22276 6141 22332
rect 6077 22272 6141 22276
rect 6157 22332 6221 22336
rect 6157 22276 6161 22332
rect 6161 22276 6217 22332
rect 6217 22276 6221 22332
rect 6157 22272 6221 22276
rect 15848 22332 15912 22336
rect 15848 22276 15852 22332
rect 15852 22276 15908 22332
rect 15908 22276 15912 22332
rect 15848 22272 15912 22276
rect 15928 22332 15992 22336
rect 15928 22276 15932 22332
rect 15932 22276 15988 22332
rect 15988 22276 15992 22332
rect 15928 22272 15992 22276
rect 16008 22332 16072 22336
rect 16008 22276 16012 22332
rect 16012 22276 16068 22332
rect 16068 22276 16072 22332
rect 16008 22272 16072 22276
rect 16088 22332 16152 22336
rect 16088 22276 16092 22332
rect 16092 22276 16148 22332
rect 16148 22276 16152 22332
rect 16088 22272 16152 22276
rect 25778 22332 25842 22336
rect 25778 22276 25782 22332
rect 25782 22276 25838 22332
rect 25838 22276 25842 22332
rect 25778 22272 25842 22276
rect 25858 22332 25922 22336
rect 25858 22276 25862 22332
rect 25862 22276 25918 22332
rect 25918 22276 25922 22332
rect 25858 22272 25922 22276
rect 25938 22332 26002 22336
rect 25938 22276 25942 22332
rect 25942 22276 25998 22332
rect 25998 22276 26002 22332
rect 25938 22272 26002 22276
rect 26018 22332 26082 22336
rect 26018 22276 26022 22332
rect 26022 22276 26078 22332
rect 26078 22276 26082 22332
rect 26018 22272 26082 22276
rect 30420 22476 30484 22540
rect 25452 22068 25516 22132
rect 26740 22128 26804 22132
rect 26740 22072 26790 22128
rect 26790 22072 26804 22128
rect 26740 22068 26804 22072
rect 27108 22068 27172 22132
rect 27844 21992 27908 21996
rect 27844 21936 27858 21992
rect 27858 21936 27908 21992
rect 27844 21932 27908 21936
rect 29132 21932 29196 21996
rect 30236 22068 30300 22132
rect 10882 21788 10946 21792
rect 10882 21732 10886 21788
rect 10886 21732 10942 21788
rect 10942 21732 10946 21788
rect 10882 21728 10946 21732
rect 10962 21788 11026 21792
rect 10962 21732 10966 21788
rect 10966 21732 11022 21788
rect 11022 21732 11026 21788
rect 10962 21728 11026 21732
rect 11042 21788 11106 21792
rect 11042 21732 11046 21788
rect 11046 21732 11102 21788
rect 11102 21732 11106 21788
rect 11042 21728 11106 21732
rect 11122 21788 11186 21792
rect 11122 21732 11126 21788
rect 11126 21732 11182 21788
rect 11182 21732 11186 21788
rect 11122 21728 11186 21732
rect 20813 21788 20877 21792
rect 20813 21732 20817 21788
rect 20817 21732 20873 21788
rect 20873 21732 20877 21788
rect 20813 21728 20877 21732
rect 20893 21788 20957 21792
rect 20893 21732 20897 21788
rect 20897 21732 20953 21788
rect 20953 21732 20957 21788
rect 20893 21728 20957 21732
rect 20973 21788 21037 21792
rect 20973 21732 20977 21788
rect 20977 21732 21033 21788
rect 21033 21732 21037 21788
rect 20973 21728 21037 21732
rect 21053 21788 21117 21792
rect 21053 21732 21057 21788
rect 21057 21732 21113 21788
rect 21113 21732 21117 21788
rect 21053 21728 21117 21732
rect 24900 21720 24964 21724
rect 24900 21664 24950 21720
rect 24950 21664 24964 21720
rect 24900 21660 24964 21664
rect 25084 21448 25148 21452
rect 25084 21392 25134 21448
rect 25134 21392 25148 21448
rect 25084 21388 25148 21392
rect 5917 21244 5981 21248
rect 5917 21188 5921 21244
rect 5921 21188 5977 21244
rect 5977 21188 5981 21244
rect 5917 21184 5981 21188
rect 5997 21244 6061 21248
rect 5997 21188 6001 21244
rect 6001 21188 6057 21244
rect 6057 21188 6061 21244
rect 5997 21184 6061 21188
rect 6077 21244 6141 21248
rect 6077 21188 6081 21244
rect 6081 21188 6137 21244
rect 6137 21188 6141 21244
rect 6077 21184 6141 21188
rect 6157 21244 6221 21248
rect 6157 21188 6161 21244
rect 6161 21188 6217 21244
rect 6217 21188 6221 21244
rect 6157 21184 6221 21188
rect 15848 21244 15912 21248
rect 15848 21188 15852 21244
rect 15852 21188 15908 21244
rect 15908 21188 15912 21244
rect 15848 21184 15912 21188
rect 15928 21244 15992 21248
rect 15928 21188 15932 21244
rect 15932 21188 15988 21244
rect 15988 21188 15992 21244
rect 15928 21184 15992 21188
rect 16008 21244 16072 21248
rect 16008 21188 16012 21244
rect 16012 21188 16068 21244
rect 16068 21188 16072 21244
rect 16008 21184 16072 21188
rect 16088 21244 16152 21248
rect 16088 21188 16092 21244
rect 16092 21188 16148 21244
rect 16148 21188 16152 21244
rect 16088 21184 16152 21188
rect 25778 21244 25842 21248
rect 25778 21188 25782 21244
rect 25782 21188 25838 21244
rect 25838 21188 25842 21244
rect 25778 21184 25842 21188
rect 25858 21244 25922 21248
rect 25858 21188 25862 21244
rect 25862 21188 25918 21244
rect 25918 21188 25922 21244
rect 25858 21184 25922 21188
rect 25938 21244 26002 21248
rect 25938 21188 25942 21244
rect 25942 21188 25998 21244
rect 25998 21188 26002 21244
rect 25938 21184 26002 21188
rect 26018 21244 26082 21248
rect 26018 21188 26022 21244
rect 26022 21188 26078 21244
rect 26078 21188 26082 21244
rect 26018 21184 26082 21188
rect 25636 20980 25700 21044
rect 26372 20768 26436 20772
rect 26372 20712 26422 20768
rect 26422 20712 26436 20768
rect 26372 20708 26436 20712
rect 10882 20700 10946 20704
rect 10882 20644 10886 20700
rect 10886 20644 10942 20700
rect 10942 20644 10946 20700
rect 10882 20640 10946 20644
rect 10962 20700 11026 20704
rect 10962 20644 10966 20700
rect 10966 20644 11022 20700
rect 11022 20644 11026 20700
rect 10962 20640 11026 20644
rect 11042 20700 11106 20704
rect 11042 20644 11046 20700
rect 11046 20644 11102 20700
rect 11102 20644 11106 20700
rect 11042 20640 11106 20644
rect 11122 20700 11186 20704
rect 11122 20644 11126 20700
rect 11126 20644 11182 20700
rect 11182 20644 11186 20700
rect 11122 20640 11186 20644
rect 20813 20700 20877 20704
rect 20813 20644 20817 20700
rect 20817 20644 20873 20700
rect 20873 20644 20877 20700
rect 20813 20640 20877 20644
rect 20893 20700 20957 20704
rect 20893 20644 20897 20700
rect 20897 20644 20953 20700
rect 20953 20644 20957 20700
rect 20893 20640 20957 20644
rect 20973 20700 21037 20704
rect 20973 20644 20977 20700
rect 20977 20644 21033 20700
rect 21033 20644 21037 20700
rect 20973 20640 21037 20644
rect 21053 20700 21117 20704
rect 21053 20644 21057 20700
rect 21057 20644 21113 20700
rect 21113 20644 21117 20700
rect 21053 20640 21117 20644
rect 5917 20156 5981 20160
rect 5917 20100 5921 20156
rect 5921 20100 5977 20156
rect 5977 20100 5981 20156
rect 5917 20096 5981 20100
rect 5997 20156 6061 20160
rect 5997 20100 6001 20156
rect 6001 20100 6057 20156
rect 6057 20100 6061 20156
rect 5997 20096 6061 20100
rect 6077 20156 6141 20160
rect 6077 20100 6081 20156
rect 6081 20100 6137 20156
rect 6137 20100 6141 20156
rect 6077 20096 6141 20100
rect 6157 20156 6221 20160
rect 6157 20100 6161 20156
rect 6161 20100 6217 20156
rect 6217 20100 6221 20156
rect 6157 20096 6221 20100
rect 15848 20156 15912 20160
rect 15848 20100 15852 20156
rect 15852 20100 15908 20156
rect 15908 20100 15912 20156
rect 15848 20096 15912 20100
rect 15928 20156 15992 20160
rect 15928 20100 15932 20156
rect 15932 20100 15988 20156
rect 15988 20100 15992 20156
rect 15928 20096 15992 20100
rect 16008 20156 16072 20160
rect 16008 20100 16012 20156
rect 16012 20100 16068 20156
rect 16068 20100 16072 20156
rect 16008 20096 16072 20100
rect 16088 20156 16152 20160
rect 16088 20100 16092 20156
rect 16092 20100 16148 20156
rect 16148 20100 16152 20156
rect 16088 20096 16152 20100
rect 25778 20156 25842 20160
rect 25778 20100 25782 20156
rect 25782 20100 25838 20156
rect 25838 20100 25842 20156
rect 25778 20096 25842 20100
rect 25858 20156 25922 20160
rect 25858 20100 25862 20156
rect 25862 20100 25918 20156
rect 25918 20100 25922 20156
rect 25858 20096 25922 20100
rect 25938 20156 26002 20160
rect 25938 20100 25942 20156
rect 25942 20100 25998 20156
rect 25998 20100 26002 20156
rect 25938 20096 26002 20100
rect 26018 20156 26082 20160
rect 26018 20100 26022 20156
rect 26022 20100 26078 20156
rect 26078 20100 26082 20156
rect 26018 20096 26082 20100
rect 30420 19756 30484 19820
rect 25268 19620 25332 19684
rect 10882 19612 10946 19616
rect 10882 19556 10886 19612
rect 10886 19556 10942 19612
rect 10942 19556 10946 19612
rect 10882 19552 10946 19556
rect 10962 19612 11026 19616
rect 10962 19556 10966 19612
rect 10966 19556 11022 19612
rect 11022 19556 11026 19612
rect 10962 19552 11026 19556
rect 11042 19612 11106 19616
rect 11042 19556 11046 19612
rect 11046 19556 11102 19612
rect 11102 19556 11106 19612
rect 11042 19552 11106 19556
rect 11122 19612 11186 19616
rect 11122 19556 11126 19612
rect 11126 19556 11182 19612
rect 11182 19556 11186 19612
rect 11122 19552 11186 19556
rect 20813 19612 20877 19616
rect 20813 19556 20817 19612
rect 20817 19556 20873 19612
rect 20873 19556 20877 19612
rect 20813 19552 20877 19556
rect 20893 19612 20957 19616
rect 20893 19556 20897 19612
rect 20897 19556 20953 19612
rect 20953 19556 20957 19612
rect 20893 19552 20957 19556
rect 20973 19612 21037 19616
rect 20973 19556 20977 19612
rect 20977 19556 21033 19612
rect 21033 19556 21037 19612
rect 20973 19552 21037 19556
rect 21053 19612 21117 19616
rect 21053 19556 21057 19612
rect 21057 19556 21113 19612
rect 21113 19556 21117 19612
rect 21053 19552 21117 19556
rect 5917 19068 5981 19072
rect 5917 19012 5921 19068
rect 5921 19012 5977 19068
rect 5977 19012 5981 19068
rect 5917 19008 5981 19012
rect 5997 19068 6061 19072
rect 5997 19012 6001 19068
rect 6001 19012 6057 19068
rect 6057 19012 6061 19068
rect 5997 19008 6061 19012
rect 6077 19068 6141 19072
rect 6077 19012 6081 19068
rect 6081 19012 6137 19068
rect 6137 19012 6141 19068
rect 6077 19008 6141 19012
rect 6157 19068 6221 19072
rect 6157 19012 6161 19068
rect 6161 19012 6217 19068
rect 6217 19012 6221 19068
rect 6157 19008 6221 19012
rect 15848 19068 15912 19072
rect 15848 19012 15852 19068
rect 15852 19012 15908 19068
rect 15908 19012 15912 19068
rect 15848 19008 15912 19012
rect 15928 19068 15992 19072
rect 15928 19012 15932 19068
rect 15932 19012 15988 19068
rect 15988 19012 15992 19068
rect 15928 19008 15992 19012
rect 16008 19068 16072 19072
rect 16008 19012 16012 19068
rect 16012 19012 16068 19068
rect 16068 19012 16072 19068
rect 16008 19008 16072 19012
rect 16088 19068 16152 19072
rect 16088 19012 16092 19068
rect 16092 19012 16148 19068
rect 16148 19012 16152 19068
rect 16088 19008 16152 19012
rect 25778 19068 25842 19072
rect 25778 19012 25782 19068
rect 25782 19012 25838 19068
rect 25838 19012 25842 19068
rect 25778 19008 25842 19012
rect 25858 19068 25922 19072
rect 25858 19012 25862 19068
rect 25862 19012 25918 19068
rect 25918 19012 25922 19068
rect 25858 19008 25922 19012
rect 25938 19068 26002 19072
rect 25938 19012 25942 19068
rect 25942 19012 25998 19068
rect 25998 19012 26002 19068
rect 25938 19008 26002 19012
rect 26018 19068 26082 19072
rect 26018 19012 26022 19068
rect 26022 19012 26078 19068
rect 26078 19012 26082 19068
rect 26018 19008 26082 19012
rect 26188 18668 26252 18732
rect 28580 18668 28644 18732
rect 10882 18524 10946 18528
rect 10882 18468 10886 18524
rect 10886 18468 10942 18524
rect 10942 18468 10946 18524
rect 10882 18464 10946 18468
rect 10962 18524 11026 18528
rect 10962 18468 10966 18524
rect 10966 18468 11022 18524
rect 11022 18468 11026 18524
rect 10962 18464 11026 18468
rect 11042 18524 11106 18528
rect 11042 18468 11046 18524
rect 11046 18468 11102 18524
rect 11102 18468 11106 18524
rect 11042 18464 11106 18468
rect 11122 18524 11186 18528
rect 11122 18468 11126 18524
rect 11126 18468 11182 18524
rect 11182 18468 11186 18524
rect 11122 18464 11186 18468
rect 20813 18524 20877 18528
rect 20813 18468 20817 18524
rect 20817 18468 20873 18524
rect 20873 18468 20877 18524
rect 20813 18464 20877 18468
rect 20893 18524 20957 18528
rect 20893 18468 20897 18524
rect 20897 18468 20953 18524
rect 20953 18468 20957 18524
rect 20893 18464 20957 18468
rect 20973 18524 21037 18528
rect 20973 18468 20977 18524
rect 20977 18468 21033 18524
rect 21033 18468 21037 18524
rect 20973 18464 21037 18468
rect 21053 18524 21117 18528
rect 21053 18468 21057 18524
rect 21057 18468 21113 18524
rect 21113 18468 21117 18524
rect 21053 18464 21117 18468
rect 25636 18124 25700 18188
rect 5917 17980 5981 17984
rect 5917 17924 5921 17980
rect 5921 17924 5977 17980
rect 5977 17924 5981 17980
rect 5917 17920 5981 17924
rect 5997 17980 6061 17984
rect 5997 17924 6001 17980
rect 6001 17924 6057 17980
rect 6057 17924 6061 17980
rect 5997 17920 6061 17924
rect 6077 17980 6141 17984
rect 6077 17924 6081 17980
rect 6081 17924 6137 17980
rect 6137 17924 6141 17980
rect 6077 17920 6141 17924
rect 6157 17980 6221 17984
rect 6157 17924 6161 17980
rect 6161 17924 6217 17980
rect 6217 17924 6221 17980
rect 6157 17920 6221 17924
rect 15848 17980 15912 17984
rect 15848 17924 15852 17980
rect 15852 17924 15908 17980
rect 15908 17924 15912 17980
rect 15848 17920 15912 17924
rect 15928 17980 15992 17984
rect 15928 17924 15932 17980
rect 15932 17924 15988 17980
rect 15988 17924 15992 17980
rect 15928 17920 15992 17924
rect 16008 17980 16072 17984
rect 16008 17924 16012 17980
rect 16012 17924 16068 17980
rect 16068 17924 16072 17980
rect 16008 17920 16072 17924
rect 16088 17980 16152 17984
rect 16088 17924 16092 17980
rect 16092 17924 16148 17980
rect 16148 17924 16152 17980
rect 16088 17920 16152 17924
rect 25778 17980 25842 17984
rect 25778 17924 25782 17980
rect 25782 17924 25838 17980
rect 25838 17924 25842 17980
rect 25778 17920 25842 17924
rect 25858 17980 25922 17984
rect 25858 17924 25862 17980
rect 25862 17924 25918 17980
rect 25918 17924 25922 17980
rect 25858 17920 25922 17924
rect 25938 17980 26002 17984
rect 25938 17924 25942 17980
rect 25942 17924 25998 17980
rect 25998 17924 26002 17980
rect 25938 17920 26002 17924
rect 26018 17980 26082 17984
rect 26018 17924 26022 17980
rect 26022 17924 26078 17980
rect 26078 17924 26082 17980
rect 26018 17920 26082 17924
rect 26188 17580 26252 17644
rect 29132 18124 29196 18188
rect 10882 17436 10946 17440
rect 10882 17380 10886 17436
rect 10886 17380 10942 17436
rect 10942 17380 10946 17436
rect 10882 17376 10946 17380
rect 10962 17436 11026 17440
rect 10962 17380 10966 17436
rect 10966 17380 11022 17436
rect 11022 17380 11026 17436
rect 10962 17376 11026 17380
rect 11042 17436 11106 17440
rect 11042 17380 11046 17436
rect 11046 17380 11102 17436
rect 11102 17380 11106 17436
rect 11042 17376 11106 17380
rect 11122 17436 11186 17440
rect 11122 17380 11126 17436
rect 11126 17380 11182 17436
rect 11182 17380 11186 17436
rect 11122 17376 11186 17380
rect 20813 17436 20877 17440
rect 20813 17380 20817 17436
rect 20817 17380 20873 17436
rect 20873 17380 20877 17436
rect 20813 17376 20877 17380
rect 20893 17436 20957 17440
rect 20893 17380 20897 17436
rect 20897 17380 20953 17436
rect 20953 17380 20957 17436
rect 20893 17376 20957 17380
rect 20973 17436 21037 17440
rect 20973 17380 20977 17436
rect 20977 17380 21033 17436
rect 21033 17380 21037 17436
rect 20973 17376 21037 17380
rect 21053 17436 21117 17440
rect 21053 17380 21057 17436
rect 21057 17380 21113 17436
rect 21113 17380 21117 17436
rect 21053 17376 21117 17380
rect 5917 16892 5981 16896
rect 5917 16836 5921 16892
rect 5921 16836 5977 16892
rect 5977 16836 5981 16892
rect 5917 16832 5981 16836
rect 5997 16892 6061 16896
rect 5997 16836 6001 16892
rect 6001 16836 6057 16892
rect 6057 16836 6061 16892
rect 5997 16832 6061 16836
rect 6077 16892 6141 16896
rect 6077 16836 6081 16892
rect 6081 16836 6137 16892
rect 6137 16836 6141 16892
rect 6077 16832 6141 16836
rect 6157 16892 6221 16896
rect 6157 16836 6161 16892
rect 6161 16836 6217 16892
rect 6217 16836 6221 16892
rect 6157 16832 6221 16836
rect 15848 16892 15912 16896
rect 15848 16836 15852 16892
rect 15852 16836 15908 16892
rect 15908 16836 15912 16892
rect 15848 16832 15912 16836
rect 15928 16892 15992 16896
rect 15928 16836 15932 16892
rect 15932 16836 15988 16892
rect 15988 16836 15992 16892
rect 15928 16832 15992 16836
rect 16008 16892 16072 16896
rect 16008 16836 16012 16892
rect 16012 16836 16068 16892
rect 16068 16836 16072 16892
rect 16008 16832 16072 16836
rect 16088 16892 16152 16896
rect 16088 16836 16092 16892
rect 16092 16836 16148 16892
rect 16148 16836 16152 16892
rect 16088 16832 16152 16836
rect 25778 16892 25842 16896
rect 25778 16836 25782 16892
rect 25782 16836 25838 16892
rect 25838 16836 25842 16892
rect 25778 16832 25842 16836
rect 25858 16892 25922 16896
rect 25858 16836 25862 16892
rect 25862 16836 25918 16892
rect 25918 16836 25922 16892
rect 25858 16832 25922 16836
rect 25938 16892 26002 16896
rect 25938 16836 25942 16892
rect 25942 16836 25998 16892
rect 25998 16836 26002 16892
rect 25938 16832 26002 16836
rect 26018 16892 26082 16896
rect 26018 16836 26022 16892
rect 26022 16836 26078 16892
rect 26078 16836 26082 16892
rect 26018 16832 26082 16836
rect 10882 16348 10946 16352
rect 10882 16292 10886 16348
rect 10886 16292 10942 16348
rect 10942 16292 10946 16348
rect 10882 16288 10946 16292
rect 10962 16348 11026 16352
rect 10962 16292 10966 16348
rect 10966 16292 11022 16348
rect 11022 16292 11026 16348
rect 10962 16288 11026 16292
rect 11042 16348 11106 16352
rect 11042 16292 11046 16348
rect 11046 16292 11102 16348
rect 11102 16292 11106 16348
rect 11042 16288 11106 16292
rect 11122 16348 11186 16352
rect 11122 16292 11126 16348
rect 11126 16292 11182 16348
rect 11182 16292 11186 16348
rect 11122 16288 11186 16292
rect 20813 16348 20877 16352
rect 20813 16292 20817 16348
rect 20817 16292 20873 16348
rect 20873 16292 20877 16348
rect 20813 16288 20877 16292
rect 20893 16348 20957 16352
rect 20893 16292 20897 16348
rect 20897 16292 20953 16348
rect 20953 16292 20957 16348
rect 20893 16288 20957 16292
rect 20973 16348 21037 16352
rect 20973 16292 20977 16348
rect 20977 16292 21033 16348
rect 21033 16292 21037 16348
rect 20973 16288 21037 16292
rect 21053 16348 21117 16352
rect 21053 16292 21057 16348
rect 21057 16292 21113 16348
rect 21113 16292 21117 16348
rect 21053 16288 21117 16292
rect 17724 16084 17788 16148
rect 5917 15804 5981 15808
rect 5917 15748 5921 15804
rect 5921 15748 5977 15804
rect 5977 15748 5981 15804
rect 5917 15744 5981 15748
rect 5997 15804 6061 15808
rect 5997 15748 6001 15804
rect 6001 15748 6057 15804
rect 6057 15748 6061 15804
rect 5997 15744 6061 15748
rect 6077 15804 6141 15808
rect 6077 15748 6081 15804
rect 6081 15748 6137 15804
rect 6137 15748 6141 15804
rect 6077 15744 6141 15748
rect 6157 15804 6221 15808
rect 6157 15748 6161 15804
rect 6161 15748 6217 15804
rect 6217 15748 6221 15804
rect 6157 15744 6221 15748
rect 15848 15804 15912 15808
rect 15848 15748 15852 15804
rect 15852 15748 15908 15804
rect 15908 15748 15912 15804
rect 15848 15744 15912 15748
rect 15928 15804 15992 15808
rect 15928 15748 15932 15804
rect 15932 15748 15988 15804
rect 15988 15748 15992 15804
rect 15928 15744 15992 15748
rect 16008 15804 16072 15808
rect 16008 15748 16012 15804
rect 16012 15748 16068 15804
rect 16068 15748 16072 15804
rect 16008 15744 16072 15748
rect 16088 15804 16152 15808
rect 16088 15748 16092 15804
rect 16092 15748 16148 15804
rect 16148 15748 16152 15804
rect 16088 15744 16152 15748
rect 25778 15804 25842 15808
rect 25778 15748 25782 15804
rect 25782 15748 25838 15804
rect 25838 15748 25842 15804
rect 25778 15744 25842 15748
rect 25858 15804 25922 15808
rect 25858 15748 25862 15804
rect 25862 15748 25918 15804
rect 25918 15748 25922 15804
rect 25858 15744 25922 15748
rect 25938 15804 26002 15808
rect 25938 15748 25942 15804
rect 25942 15748 25998 15804
rect 25998 15748 26002 15804
rect 25938 15744 26002 15748
rect 26018 15804 26082 15808
rect 26018 15748 26022 15804
rect 26022 15748 26078 15804
rect 26078 15748 26082 15804
rect 26018 15744 26082 15748
rect 29500 15404 29564 15468
rect 25636 15328 25700 15332
rect 25636 15272 25650 15328
rect 25650 15272 25700 15328
rect 25636 15268 25700 15272
rect 10882 15260 10946 15264
rect 10882 15204 10886 15260
rect 10886 15204 10942 15260
rect 10942 15204 10946 15260
rect 10882 15200 10946 15204
rect 10962 15260 11026 15264
rect 10962 15204 10966 15260
rect 10966 15204 11022 15260
rect 11022 15204 11026 15260
rect 10962 15200 11026 15204
rect 11042 15260 11106 15264
rect 11042 15204 11046 15260
rect 11046 15204 11102 15260
rect 11102 15204 11106 15260
rect 11042 15200 11106 15204
rect 11122 15260 11186 15264
rect 11122 15204 11126 15260
rect 11126 15204 11182 15260
rect 11182 15204 11186 15260
rect 11122 15200 11186 15204
rect 20813 15260 20877 15264
rect 20813 15204 20817 15260
rect 20817 15204 20873 15260
rect 20873 15204 20877 15260
rect 20813 15200 20877 15204
rect 20893 15260 20957 15264
rect 20893 15204 20897 15260
rect 20897 15204 20953 15260
rect 20953 15204 20957 15260
rect 20893 15200 20957 15204
rect 20973 15260 21037 15264
rect 20973 15204 20977 15260
rect 20977 15204 21033 15260
rect 21033 15204 21037 15260
rect 20973 15200 21037 15204
rect 21053 15260 21117 15264
rect 21053 15204 21057 15260
rect 21057 15204 21113 15260
rect 21113 15204 21117 15260
rect 21053 15200 21117 15204
rect 28396 15132 28460 15196
rect 5917 14716 5981 14720
rect 5917 14660 5921 14716
rect 5921 14660 5977 14716
rect 5977 14660 5981 14716
rect 5917 14656 5981 14660
rect 5997 14716 6061 14720
rect 5997 14660 6001 14716
rect 6001 14660 6057 14716
rect 6057 14660 6061 14716
rect 5997 14656 6061 14660
rect 6077 14716 6141 14720
rect 6077 14660 6081 14716
rect 6081 14660 6137 14716
rect 6137 14660 6141 14716
rect 6077 14656 6141 14660
rect 6157 14716 6221 14720
rect 6157 14660 6161 14716
rect 6161 14660 6217 14716
rect 6217 14660 6221 14716
rect 6157 14656 6221 14660
rect 15848 14716 15912 14720
rect 15848 14660 15852 14716
rect 15852 14660 15908 14716
rect 15908 14660 15912 14716
rect 15848 14656 15912 14660
rect 15928 14716 15992 14720
rect 15928 14660 15932 14716
rect 15932 14660 15988 14716
rect 15988 14660 15992 14716
rect 15928 14656 15992 14660
rect 16008 14716 16072 14720
rect 16008 14660 16012 14716
rect 16012 14660 16068 14716
rect 16068 14660 16072 14716
rect 16008 14656 16072 14660
rect 16088 14716 16152 14720
rect 16088 14660 16092 14716
rect 16092 14660 16148 14716
rect 16148 14660 16152 14716
rect 16088 14656 16152 14660
rect 25778 14716 25842 14720
rect 25778 14660 25782 14716
rect 25782 14660 25838 14716
rect 25838 14660 25842 14716
rect 25778 14656 25842 14660
rect 25858 14716 25922 14720
rect 25858 14660 25862 14716
rect 25862 14660 25918 14716
rect 25918 14660 25922 14716
rect 25858 14656 25922 14660
rect 25938 14716 26002 14720
rect 25938 14660 25942 14716
rect 25942 14660 25998 14716
rect 25998 14660 26002 14716
rect 25938 14656 26002 14660
rect 26018 14716 26082 14720
rect 26018 14660 26022 14716
rect 26022 14660 26078 14716
rect 26078 14660 26082 14716
rect 26018 14656 26082 14660
rect 10882 14172 10946 14176
rect 10882 14116 10886 14172
rect 10886 14116 10942 14172
rect 10942 14116 10946 14172
rect 10882 14112 10946 14116
rect 10962 14172 11026 14176
rect 10962 14116 10966 14172
rect 10966 14116 11022 14172
rect 11022 14116 11026 14172
rect 10962 14112 11026 14116
rect 11042 14172 11106 14176
rect 11042 14116 11046 14172
rect 11046 14116 11102 14172
rect 11102 14116 11106 14172
rect 11042 14112 11106 14116
rect 11122 14172 11186 14176
rect 11122 14116 11126 14172
rect 11126 14116 11182 14172
rect 11182 14116 11186 14172
rect 11122 14112 11186 14116
rect 20813 14172 20877 14176
rect 20813 14116 20817 14172
rect 20817 14116 20873 14172
rect 20873 14116 20877 14172
rect 20813 14112 20877 14116
rect 20893 14172 20957 14176
rect 20893 14116 20897 14172
rect 20897 14116 20953 14172
rect 20953 14116 20957 14172
rect 20893 14112 20957 14116
rect 20973 14172 21037 14176
rect 20973 14116 20977 14172
rect 20977 14116 21033 14172
rect 21033 14116 21037 14172
rect 20973 14112 21037 14116
rect 21053 14172 21117 14176
rect 21053 14116 21057 14172
rect 21057 14116 21113 14172
rect 21113 14116 21117 14172
rect 21053 14112 21117 14116
rect 29316 14044 29380 14108
rect 5917 13628 5981 13632
rect 5917 13572 5921 13628
rect 5921 13572 5977 13628
rect 5977 13572 5981 13628
rect 5917 13568 5981 13572
rect 5997 13628 6061 13632
rect 5997 13572 6001 13628
rect 6001 13572 6057 13628
rect 6057 13572 6061 13628
rect 5997 13568 6061 13572
rect 6077 13628 6141 13632
rect 6077 13572 6081 13628
rect 6081 13572 6137 13628
rect 6137 13572 6141 13628
rect 6077 13568 6141 13572
rect 6157 13628 6221 13632
rect 6157 13572 6161 13628
rect 6161 13572 6217 13628
rect 6217 13572 6221 13628
rect 6157 13568 6221 13572
rect 15848 13628 15912 13632
rect 15848 13572 15852 13628
rect 15852 13572 15908 13628
rect 15908 13572 15912 13628
rect 15848 13568 15912 13572
rect 15928 13628 15992 13632
rect 15928 13572 15932 13628
rect 15932 13572 15988 13628
rect 15988 13572 15992 13628
rect 15928 13568 15992 13572
rect 16008 13628 16072 13632
rect 16008 13572 16012 13628
rect 16012 13572 16068 13628
rect 16068 13572 16072 13628
rect 16008 13568 16072 13572
rect 16088 13628 16152 13632
rect 16088 13572 16092 13628
rect 16092 13572 16148 13628
rect 16148 13572 16152 13628
rect 16088 13568 16152 13572
rect 25778 13628 25842 13632
rect 25778 13572 25782 13628
rect 25782 13572 25838 13628
rect 25838 13572 25842 13628
rect 25778 13568 25842 13572
rect 25858 13628 25922 13632
rect 25858 13572 25862 13628
rect 25862 13572 25918 13628
rect 25918 13572 25922 13628
rect 25858 13568 25922 13572
rect 25938 13628 26002 13632
rect 25938 13572 25942 13628
rect 25942 13572 25998 13628
rect 25998 13572 26002 13628
rect 25938 13568 26002 13572
rect 26018 13628 26082 13632
rect 26018 13572 26022 13628
rect 26022 13572 26078 13628
rect 26078 13572 26082 13628
rect 26018 13568 26082 13572
rect 10882 13084 10946 13088
rect 10882 13028 10886 13084
rect 10886 13028 10942 13084
rect 10942 13028 10946 13084
rect 10882 13024 10946 13028
rect 10962 13084 11026 13088
rect 10962 13028 10966 13084
rect 10966 13028 11022 13084
rect 11022 13028 11026 13084
rect 10962 13024 11026 13028
rect 11042 13084 11106 13088
rect 11042 13028 11046 13084
rect 11046 13028 11102 13084
rect 11102 13028 11106 13084
rect 11042 13024 11106 13028
rect 11122 13084 11186 13088
rect 11122 13028 11126 13084
rect 11126 13028 11182 13084
rect 11182 13028 11186 13084
rect 11122 13024 11186 13028
rect 20813 13084 20877 13088
rect 20813 13028 20817 13084
rect 20817 13028 20873 13084
rect 20873 13028 20877 13084
rect 20813 13024 20877 13028
rect 20893 13084 20957 13088
rect 20893 13028 20897 13084
rect 20897 13028 20953 13084
rect 20953 13028 20957 13084
rect 20893 13024 20957 13028
rect 20973 13084 21037 13088
rect 20973 13028 20977 13084
rect 20977 13028 21033 13084
rect 21033 13028 21037 13084
rect 20973 13024 21037 13028
rect 21053 13084 21117 13088
rect 21053 13028 21057 13084
rect 21057 13028 21113 13084
rect 21113 13028 21117 13084
rect 21053 13024 21117 13028
rect 5917 12540 5981 12544
rect 5917 12484 5921 12540
rect 5921 12484 5977 12540
rect 5977 12484 5981 12540
rect 5917 12480 5981 12484
rect 5997 12540 6061 12544
rect 5997 12484 6001 12540
rect 6001 12484 6057 12540
rect 6057 12484 6061 12540
rect 5997 12480 6061 12484
rect 6077 12540 6141 12544
rect 6077 12484 6081 12540
rect 6081 12484 6137 12540
rect 6137 12484 6141 12540
rect 6077 12480 6141 12484
rect 6157 12540 6221 12544
rect 6157 12484 6161 12540
rect 6161 12484 6217 12540
rect 6217 12484 6221 12540
rect 6157 12480 6221 12484
rect 15848 12540 15912 12544
rect 15848 12484 15852 12540
rect 15852 12484 15908 12540
rect 15908 12484 15912 12540
rect 15848 12480 15912 12484
rect 15928 12540 15992 12544
rect 15928 12484 15932 12540
rect 15932 12484 15988 12540
rect 15988 12484 15992 12540
rect 15928 12480 15992 12484
rect 16008 12540 16072 12544
rect 16008 12484 16012 12540
rect 16012 12484 16068 12540
rect 16068 12484 16072 12540
rect 16008 12480 16072 12484
rect 16088 12540 16152 12544
rect 16088 12484 16092 12540
rect 16092 12484 16148 12540
rect 16148 12484 16152 12540
rect 16088 12480 16152 12484
rect 25778 12540 25842 12544
rect 25778 12484 25782 12540
rect 25782 12484 25838 12540
rect 25838 12484 25842 12540
rect 25778 12480 25842 12484
rect 25858 12540 25922 12544
rect 25858 12484 25862 12540
rect 25862 12484 25918 12540
rect 25918 12484 25922 12540
rect 25858 12480 25922 12484
rect 25938 12540 26002 12544
rect 25938 12484 25942 12540
rect 25942 12484 25998 12540
rect 25998 12484 26002 12540
rect 25938 12480 26002 12484
rect 26018 12540 26082 12544
rect 26018 12484 26022 12540
rect 26022 12484 26078 12540
rect 26078 12484 26082 12540
rect 26018 12480 26082 12484
rect 26188 12064 26252 12068
rect 26188 12008 26202 12064
rect 26202 12008 26252 12064
rect 26188 12004 26252 12008
rect 10882 11996 10946 12000
rect 10882 11940 10886 11996
rect 10886 11940 10942 11996
rect 10942 11940 10946 11996
rect 10882 11936 10946 11940
rect 10962 11996 11026 12000
rect 10962 11940 10966 11996
rect 10966 11940 11022 11996
rect 11022 11940 11026 11996
rect 10962 11936 11026 11940
rect 11042 11996 11106 12000
rect 11042 11940 11046 11996
rect 11046 11940 11102 11996
rect 11102 11940 11106 11996
rect 11042 11936 11106 11940
rect 11122 11996 11186 12000
rect 11122 11940 11126 11996
rect 11126 11940 11182 11996
rect 11182 11940 11186 11996
rect 11122 11936 11186 11940
rect 20813 11996 20877 12000
rect 20813 11940 20817 11996
rect 20817 11940 20873 11996
rect 20873 11940 20877 11996
rect 20813 11936 20877 11940
rect 20893 11996 20957 12000
rect 20893 11940 20897 11996
rect 20897 11940 20953 11996
rect 20953 11940 20957 11996
rect 20893 11936 20957 11940
rect 20973 11996 21037 12000
rect 20973 11940 20977 11996
rect 20977 11940 21033 11996
rect 21033 11940 21037 11996
rect 20973 11936 21037 11940
rect 21053 11996 21117 12000
rect 21053 11940 21057 11996
rect 21057 11940 21113 11996
rect 21113 11940 21117 11996
rect 21053 11936 21117 11940
rect 5917 11452 5981 11456
rect 5917 11396 5921 11452
rect 5921 11396 5977 11452
rect 5977 11396 5981 11452
rect 5917 11392 5981 11396
rect 5997 11452 6061 11456
rect 5997 11396 6001 11452
rect 6001 11396 6057 11452
rect 6057 11396 6061 11452
rect 5997 11392 6061 11396
rect 6077 11452 6141 11456
rect 6077 11396 6081 11452
rect 6081 11396 6137 11452
rect 6137 11396 6141 11452
rect 6077 11392 6141 11396
rect 6157 11452 6221 11456
rect 6157 11396 6161 11452
rect 6161 11396 6217 11452
rect 6217 11396 6221 11452
rect 6157 11392 6221 11396
rect 15848 11452 15912 11456
rect 15848 11396 15852 11452
rect 15852 11396 15908 11452
rect 15908 11396 15912 11452
rect 15848 11392 15912 11396
rect 15928 11452 15992 11456
rect 15928 11396 15932 11452
rect 15932 11396 15988 11452
rect 15988 11396 15992 11452
rect 15928 11392 15992 11396
rect 16008 11452 16072 11456
rect 16008 11396 16012 11452
rect 16012 11396 16068 11452
rect 16068 11396 16072 11452
rect 16008 11392 16072 11396
rect 16088 11452 16152 11456
rect 16088 11396 16092 11452
rect 16092 11396 16148 11452
rect 16148 11396 16152 11452
rect 16088 11392 16152 11396
rect 25778 11452 25842 11456
rect 25778 11396 25782 11452
rect 25782 11396 25838 11452
rect 25838 11396 25842 11452
rect 25778 11392 25842 11396
rect 25858 11452 25922 11456
rect 25858 11396 25862 11452
rect 25862 11396 25918 11452
rect 25918 11396 25922 11452
rect 25858 11392 25922 11396
rect 25938 11452 26002 11456
rect 25938 11396 25942 11452
rect 25942 11396 25998 11452
rect 25998 11396 26002 11452
rect 25938 11392 26002 11396
rect 26018 11452 26082 11456
rect 26018 11396 26022 11452
rect 26022 11396 26078 11452
rect 26078 11396 26082 11452
rect 26018 11392 26082 11396
rect 10882 10908 10946 10912
rect 10882 10852 10886 10908
rect 10886 10852 10942 10908
rect 10942 10852 10946 10908
rect 10882 10848 10946 10852
rect 10962 10908 11026 10912
rect 10962 10852 10966 10908
rect 10966 10852 11022 10908
rect 11022 10852 11026 10908
rect 10962 10848 11026 10852
rect 11042 10908 11106 10912
rect 11042 10852 11046 10908
rect 11046 10852 11102 10908
rect 11102 10852 11106 10908
rect 11042 10848 11106 10852
rect 11122 10908 11186 10912
rect 11122 10852 11126 10908
rect 11126 10852 11182 10908
rect 11182 10852 11186 10908
rect 11122 10848 11186 10852
rect 20813 10908 20877 10912
rect 20813 10852 20817 10908
rect 20817 10852 20873 10908
rect 20873 10852 20877 10908
rect 20813 10848 20877 10852
rect 20893 10908 20957 10912
rect 20893 10852 20897 10908
rect 20897 10852 20953 10908
rect 20953 10852 20957 10908
rect 20893 10848 20957 10852
rect 20973 10908 21037 10912
rect 20973 10852 20977 10908
rect 20977 10852 21033 10908
rect 21033 10852 21037 10908
rect 20973 10848 21037 10852
rect 21053 10908 21117 10912
rect 21053 10852 21057 10908
rect 21057 10852 21113 10908
rect 21113 10852 21117 10908
rect 21053 10848 21117 10852
rect 5917 10364 5981 10368
rect 5917 10308 5921 10364
rect 5921 10308 5977 10364
rect 5977 10308 5981 10364
rect 5917 10304 5981 10308
rect 5997 10364 6061 10368
rect 5997 10308 6001 10364
rect 6001 10308 6057 10364
rect 6057 10308 6061 10364
rect 5997 10304 6061 10308
rect 6077 10364 6141 10368
rect 6077 10308 6081 10364
rect 6081 10308 6137 10364
rect 6137 10308 6141 10364
rect 6077 10304 6141 10308
rect 6157 10364 6221 10368
rect 6157 10308 6161 10364
rect 6161 10308 6217 10364
rect 6217 10308 6221 10364
rect 6157 10304 6221 10308
rect 15848 10364 15912 10368
rect 15848 10308 15852 10364
rect 15852 10308 15908 10364
rect 15908 10308 15912 10364
rect 15848 10304 15912 10308
rect 15928 10364 15992 10368
rect 15928 10308 15932 10364
rect 15932 10308 15988 10364
rect 15988 10308 15992 10364
rect 15928 10304 15992 10308
rect 16008 10364 16072 10368
rect 16008 10308 16012 10364
rect 16012 10308 16068 10364
rect 16068 10308 16072 10364
rect 16008 10304 16072 10308
rect 16088 10364 16152 10368
rect 16088 10308 16092 10364
rect 16092 10308 16148 10364
rect 16148 10308 16152 10364
rect 16088 10304 16152 10308
rect 25778 10364 25842 10368
rect 25778 10308 25782 10364
rect 25782 10308 25838 10364
rect 25838 10308 25842 10364
rect 25778 10304 25842 10308
rect 25858 10364 25922 10368
rect 25858 10308 25862 10364
rect 25862 10308 25918 10364
rect 25918 10308 25922 10364
rect 25858 10304 25922 10308
rect 25938 10364 26002 10368
rect 25938 10308 25942 10364
rect 25942 10308 25998 10364
rect 25998 10308 26002 10364
rect 25938 10304 26002 10308
rect 26018 10364 26082 10368
rect 26018 10308 26022 10364
rect 26022 10308 26078 10364
rect 26078 10308 26082 10364
rect 26018 10304 26082 10308
rect 10882 9820 10946 9824
rect 10882 9764 10886 9820
rect 10886 9764 10942 9820
rect 10942 9764 10946 9820
rect 10882 9760 10946 9764
rect 10962 9820 11026 9824
rect 10962 9764 10966 9820
rect 10966 9764 11022 9820
rect 11022 9764 11026 9820
rect 10962 9760 11026 9764
rect 11042 9820 11106 9824
rect 11042 9764 11046 9820
rect 11046 9764 11102 9820
rect 11102 9764 11106 9820
rect 11042 9760 11106 9764
rect 11122 9820 11186 9824
rect 11122 9764 11126 9820
rect 11126 9764 11182 9820
rect 11182 9764 11186 9820
rect 11122 9760 11186 9764
rect 20813 9820 20877 9824
rect 20813 9764 20817 9820
rect 20817 9764 20873 9820
rect 20873 9764 20877 9820
rect 20813 9760 20877 9764
rect 20893 9820 20957 9824
rect 20893 9764 20897 9820
rect 20897 9764 20953 9820
rect 20953 9764 20957 9820
rect 20893 9760 20957 9764
rect 20973 9820 21037 9824
rect 20973 9764 20977 9820
rect 20977 9764 21033 9820
rect 21033 9764 21037 9820
rect 20973 9760 21037 9764
rect 21053 9820 21117 9824
rect 21053 9764 21057 9820
rect 21057 9764 21113 9820
rect 21113 9764 21117 9820
rect 21053 9760 21117 9764
rect 5917 9276 5981 9280
rect 5917 9220 5921 9276
rect 5921 9220 5977 9276
rect 5977 9220 5981 9276
rect 5917 9216 5981 9220
rect 5997 9276 6061 9280
rect 5997 9220 6001 9276
rect 6001 9220 6057 9276
rect 6057 9220 6061 9276
rect 5997 9216 6061 9220
rect 6077 9276 6141 9280
rect 6077 9220 6081 9276
rect 6081 9220 6137 9276
rect 6137 9220 6141 9276
rect 6077 9216 6141 9220
rect 6157 9276 6221 9280
rect 6157 9220 6161 9276
rect 6161 9220 6217 9276
rect 6217 9220 6221 9276
rect 6157 9216 6221 9220
rect 15848 9276 15912 9280
rect 15848 9220 15852 9276
rect 15852 9220 15908 9276
rect 15908 9220 15912 9276
rect 15848 9216 15912 9220
rect 15928 9276 15992 9280
rect 15928 9220 15932 9276
rect 15932 9220 15988 9276
rect 15988 9220 15992 9276
rect 15928 9216 15992 9220
rect 16008 9276 16072 9280
rect 16008 9220 16012 9276
rect 16012 9220 16068 9276
rect 16068 9220 16072 9276
rect 16008 9216 16072 9220
rect 16088 9276 16152 9280
rect 16088 9220 16092 9276
rect 16092 9220 16148 9276
rect 16148 9220 16152 9276
rect 16088 9216 16152 9220
rect 25778 9276 25842 9280
rect 25778 9220 25782 9276
rect 25782 9220 25838 9276
rect 25838 9220 25842 9276
rect 25778 9216 25842 9220
rect 25858 9276 25922 9280
rect 25858 9220 25862 9276
rect 25862 9220 25918 9276
rect 25918 9220 25922 9276
rect 25858 9216 25922 9220
rect 25938 9276 26002 9280
rect 25938 9220 25942 9276
rect 25942 9220 25998 9276
rect 25998 9220 26002 9276
rect 25938 9216 26002 9220
rect 26018 9276 26082 9280
rect 26018 9220 26022 9276
rect 26022 9220 26078 9276
rect 26078 9220 26082 9276
rect 26018 9216 26082 9220
rect 10882 8732 10946 8736
rect 10882 8676 10886 8732
rect 10886 8676 10942 8732
rect 10942 8676 10946 8732
rect 10882 8672 10946 8676
rect 10962 8732 11026 8736
rect 10962 8676 10966 8732
rect 10966 8676 11022 8732
rect 11022 8676 11026 8732
rect 10962 8672 11026 8676
rect 11042 8732 11106 8736
rect 11042 8676 11046 8732
rect 11046 8676 11102 8732
rect 11102 8676 11106 8732
rect 11042 8672 11106 8676
rect 11122 8732 11186 8736
rect 11122 8676 11126 8732
rect 11126 8676 11182 8732
rect 11182 8676 11186 8732
rect 11122 8672 11186 8676
rect 20813 8732 20877 8736
rect 20813 8676 20817 8732
rect 20817 8676 20873 8732
rect 20873 8676 20877 8732
rect 20813 8672 20877 8676
rect 20893 8732 20957 8736
rect 20893 8676 20897 8732
rect 20897 8676 20953 8732
rect 20953 8676 20957 8732
rect 20893 8672 20957 8676
rect 20973 8732 21037 8736
rect 20973 8676 20977 8732
rect 20977 8676 21033 8732
rect 21033 8676 21037 8732
rect 20973 8672 21037 8676
rect 21053 8732 21117 8736
rect 21053 8676 21057 8732
rect 21057 8676 21113 8732
rect 21113 8676 21117 8732
rect 21053 8672 21117 8676
rect 5917 8188 5981 8192
rect 5917 8132 5921 8188
rect 5921 8132 5977 8188
rect 5977 8132 5981 8188
rect 5917 8128 5981 8132
rect 5997 8188 6061 8192
rect 5997 8132 6001 8188
rect 6001 8132 6057 8188
rect 6057 8132 6061 8188
rect 5997 8128 6061 8132
rect 6077 8188 6141 8192
rect 6077 8132 6081 8188
rect 6081 8132 6137 8188
rect 6137 8132 6141 8188
rect 6077 8128 6141 8132
rect 6157 8188 6221 8192
rect 6157 8132 6161 8188
rect 6161 8132 6217 8188
rect 6217 8132 6221 8188
rect 6157 8128 6221 8132
rect 15848 8188 15912 8192
rect 15848 8132 15852 8188
rect 15852 8132 15908 8188
rect 15908 8132 15912 8188
rect 15848 8128 15912 8132
rect 15928 8188 15992 8192
rect 15928 8132 15932 8188
rect 15932 8132 15988 8188
rect 15988 8132 15992 8188
rect 15928 8128 15992 8132
rect 16008 8188 16072 8192
rect 16008 8132 16012 8188
rect 16012 8132 16068 8188
rect 16068 8132 16072 8188
rect 16008 8128 16072 8132
rect 16088 8188 16152 8192
rect 16088 8132 16092 8188
rect 16092 8132 16148 8188
rect 16148 8132 16152 8188
rect 16088 8128 16152 8132
rect 25778 8188 25842 8192
rect 25778 8132 25782 8188
rect 25782 8132 25838 8188
rect 25838 8132 25842 8188
rect 25778 8128 25842 8132
rect 25858 8188 25922 8192
rect 25858 8132 25862 8188
rect 25862 8132 25918 8188
rect 25918 8132 25922 8188
rect 25858 8128 25922 8132
rect 25938 8188 26002 8192
rect 25938 8132 25942 8188
rect 25942 8132 25998 8188
rect 25998 8132 26002 8188
rect 25938 8128 26002 8132
rect 26018 8188 26082 8192
rect 26018 8132 26022 8188
rect 26022 8132 26078 8188
rect 26078 8132 26082 8188
rect 26018 8128 26082 8132
rect 10882 7644 10946 7648
rect 10882 7588 10886 7644
rect 10886 7588 10942 7644
rect 10942 7588 10946 7644
rect 10882 7584 10946 7588
rect 10962 7644 11026 7648
rect 10962 7588 10966 7644
rect 10966 7588 11022 7644
rect 11022 7588 11026 7644
rect 10962 7584 11026 7588
rect 11042 7644 11106 7648
rect 11042 7588 11046 7644
rect 11046 7588 11102 7644
rect 11102 7588 11106 7644
rect 11042 7584 11106 7588
rect 11122 7644 11186 7648
rect 11122 7588 11126 7644
rect 11126 7588 11182 7644
rect 11182 7588 11186 7644
rect 11122 7584 11186 7588
rect 20813 7644 20877 7648
rect 20813 7588 20817 7644
rect 20817 7588 20873 7644
rect 20873 7588 20877 7644
rect 20813 7584 20877 7588
rect 20893 7644 20957 7648
rect 20893 7588 20897 7644
rect 20897 7588 20953 7644
rect 20953 7588 20957 7644
rect 20893 7584 20957 7588
rect 20973 7644 21037 7648
rect 20973 7588 20977 7644
rect 20977 7588 21033 7644
rect 21033 7588 21037 7644
rect 20973 7584 21037 7588
rect 21053 7644 21117 7648
rect 21053 7588 21057 7644
rect 21057 7588 21113 7644
rect 21113 7588 21117 7644
rect 21053 7584 21117 7588
rect 5917 7100 5981 7104
rect 5917 7044 5921 7100
rect 5921 7044 5977 7100
rect 5977 7044 5981 7100
rect 5917 7040 5981 7044
rect 5997 7100 6061 7104
rect 5997 7044 6001 7100
rect 6001 7044 6057 7100
rect 6057 7044 6061 7100
rect 5997 7040 6061 7044
rect 6077 7100 6141 7104
rect 6077 7044 6081 7100
rect 6081 7044 6137 7100
rect 6137 7044 6141 7100
rect 6077 7040 6141 7044
rect 6157 7100 6221 7104
rect 6157 7044 6161 7100
rect 6161 7044 6217 7100
rect 6217 7044 6221 7100
rect 6157 7040 6221 7044
rect 15848 7100 15912 7104
rect 15848 7044 15852 7100
rect 15852 7044 15908 7100
rect 15908 7044 15912 7100
rect 15848 7040 15912 7044
rect 15928 7100 15992 7104
rect 15928 7044 15932 7100
rect 15932 7044 15988 7100
rect 15988 7044 15992 7100
rect 15928 7040 15992 7044
rect 16008 7100 16072 7104
rect 16008 7044 16012 7100
rect 16012 7044 16068 7100
rect 16068 7044 16072 7100
rect 16008 7040 16072 7044
rect 16088 7100 16152 7104
rect 16088 7044 16092 7100
rect 16092 7044 16148 7100
rect 16148 7044 16152 7100
rect 16088 7040 16152 7044
rect 25778 7100 25842 7104
rect 25778 7044 25782 7100
rect 25782 7044 25838 7100
rect 25838 7044 25842 7100
rect 25778 7040 25842 7044
rect 25858 7100 25922 7104
rect 25858 7044 25862 7100
rect 25862 7044 25918 7100
rect 25918 7044 25922 7100
rect 25858 7040 25922 7044
rect 25938 7100 26002 7104
rect 25938 7044 25942 7100
rect 25942 7044 25998 7100
rect 25998 7044 26002 7100
rect 25938 7040 26002 7044
rect 26018 7100 26082 7104
rect 26018 7044 26022 7100
rect 26022 7044 26078 7100
rect 26078 7044 26082 7100
rect 26018 7040 26082 7044
rect 10882 6556 10946 6560
rect 10882 6500 10886 6556
rect 10886 6500 10942 6556
rect 10942 6500 10946 6556
rect 10882 6496 10946 6500
rect 10962 6556 11026 6560
rect 10962 6500 10966 6556
rect 10966 6500 11022 6556
rect 11022 6500 11026 6556
rect 10962 6496 11026 6500
rect 11042 6556 11106 6560
rect 11042 6500 11046 6556
rect 11046 6500 11102 6556
rect 11102 6500 11106 6556
rect 11042 6496 11106 6500
rect 11122 6556 11186 6560
rect 11122 6500 11126 6556
rect 11126 6500 11182 6556
rect 11182 6500 11186 6556
rect 11122 6496 11186 6500
rect 20813 6556 20877 6560
rect 20813 6500 20817 6556
rect 20817 6500 20873 6556
rect 20873 6500 20877 6556
rect 20813 6496 20877 6500
rect 20893 6556 20957 6560
rect 20893 6500 20897 6556
rect 20897 6500 20953 6556
rect 20953 6500 20957 6556
rect 20893 6496 20957 6500
rect 20973 6556 21037 6560
rect 20973 6500 20977 6556
rect 20977 6500 21033 6556
rect 21033 6500 21037 6556
rect 20973 6496 21037 6500
rect 21053 6556 21117 6560
rect 21053 6500 21057 6556
rect 21057 6500 21113 6556
rect 21113 6500 21117 6556
rect 21053 6496 21117 6500
rect 30052 6428 30116 6492
rect 5917 6012 5981 6016
rect 5917 5956 5921 6012
rect 5921 5956 5977 6012
rect 5977 5956 5981 6012
rect 5917 5952 5981 5956
rect 5997 6012 6061 6016
rect 5997 5956 6001 6012
rect 6001 5956 6057 6012
rect 6057 5956 6061 6012
rect 5997 5952 6061 5956
rect 6077 6012 6141 6016
rect 6077 5956 6081 6012
rect 6081 5956 6137 6012
rect 6137 5956 6141 6012
rect 6077 5952 6141 5956
rect 6157 6012 6221 6016
rect 6157 5956 6161 6012
rect 6161 5956 6217 6012
rect 6217 5956 6221 6012
rect 6157 5952 6221 5956
rect 15848 6012 15912 6016
rect 15848 5956 15852 6012
rect 15852 5956 15908 6012
rect 15908 5956 15912 6012
rect 15848 5952 15912 5956
rect 15928 6012 15992 6016
rect 15928 5956 15932 6012
rect 15932 5956 15988 6012
rect 15988 5956 15992 6012
rect 15928 5952 15992 5956
rect 16008 6012 16072 6016
rect 16008 5956 16012 6012
rect 16012 5956 16068 6012
rect 16068 5956 16072 6012
rect 16008 5952 16072 5956
rect 16088 6012 16152 6016
rect 16088 5956 16092 6012
rect 16092 5956 16148 6012
rect 16148 5956 16152 6012
rect 16088 5952 16152 5956
rect 25778 6012 25842 6016
rect 25778 5956 25782 6012
rect 25782 5956 25838 6012
rect 25838 5956 25842 6012
rect 25778 5952 25842 5956
rect 25858 6012 25922 6016
rect 25858 5956 25862 6012
rect 25862 5956 25918 6012
rect 25918 5956 25922 6012
rect 25858 5952 25922 5956
rect 25938 6012 26002 6016
rect 25938 5956 25942 6012
rect 25942 5956 25998 6012
rect 25998 5956 26002 6012
rect 25938 5952 26002 5956
rect 26018 6012 26082 6016
rect 26018 5956 26022 6012
rect 26022 5956 26078 6012
rect 26078 5956 26082 6012
rect 26018 5952 26082 5956
rect 10882 5468 10946 5472
rect 10882 5412 10886 5468
rect 10886 5412 10942 5468
rect 10942 5412 10946 5468
rect 10882 5408 10946 5412
rect 10962 5468 11026 5472
rect 10962 5412 10966 5468
rect 10966 5412 11022 5468
rect 11022 5412 11026 5468
rect 10962 5408 11026 5412
rect 11042 5468 11106 5472
rect 11042 5412 11046 5468
rect 11046 5412 11102 5468
rect 11102 5412 11106 5468
rect 11042 5408 11106 5412
rect 11122 5468 11186 5472
rect 11122 5412 11126 5468
rect 11126 5412 11182 5468
rect 11182 5412 11186 5468
rect 11122 5408 11186 5412
rect 20813 5468 20877 5472
rect 20813 5412 20817 5468
rect 20817 5412 20873 5468
rect 20873 5412 20877 5468
rect 20813 5408 20877 5412
rect 20893 5468 20957 5472
rect 20893 5412 20897 5468
rect 20897 5412 20953 5468
rect 20953 5412 20957 5468
rect 20893 5408 20957 5412
rect 20973 5468 21037 5472
rect 20973 5412 20977 5468
rect 20977 5412 21033 5468
rect 21033 5412 21037 5468
rect 20973 5408 21037 5412
rect 21053 5468 21117 5472
rect 21053 5412 21057 5468
rect 21057 5412 21113 5468
rect 21113 5412 21117 5468
rect 21053 5408 21117 5412
rect 29684 5340 29748 5404
rect 5917 4924 5981 4928
rect 5917 4868 5921 4924
rect 5921 4868 5977 4924
rect 5977 4868 5981 4924
rect 5917 4864 5981 4868
rect 5997 4924 6061 4928
rect 5997 4868 6001 4924
rect 6001 4868 6057 4924
rect 6057 4868 6061 4924
rect 5997 4864 6061 4868
rect 6077 4924 6141 4928
rect 6077 4868 6081 4924
rect 6081 4868 6137 4924
rect 6137 4868 6141 4924
rect 6077 4864 6141 4868
rect 6157 4924 6221 4928
rect 6157 4868 6161 4924
rect 6161 4868 6217 4924
rect 6217 4868 6221 4924
rect 6157 4864 6221 4868
rect 15848 4924 15912 4928
rect 15848 4868 15852 4924
rect 15852 4868 15908 4924
rect 15908 4868 15912 4924
rect 15848 4864 15912 4868
rect 15928 4924 15992 4928
rect 15928 4868 15932 4924
rect 15932 4868 15988 4924
rect 15988 4868 15992 4924
rect 15928 4864 15992 4868
rect 16008 4924 16072 4928
rect 16008 4868 16012 4924
rect 16012 4868 16068 4924
rect 16068 4868 16072 4924
rect 16008 4864 16072 4868
rect 16088 4924 16152 4928
rect 16088 4868 16092 4924
rect 16092 4868 16148 4924
rect 16148 4868 16152 4924
rect 16088 4864 16152 4868
rect 25778 4924 25842 4928
rect 25778 4868 25782 4924
rect 25782 4868 25838 4924
rect 25838 4868 25842 4924
rect 25778 4864 25842 4868
rect 25858 4924 25922 4928
rect 25858 4868 25862 4924
rect 25862 4868 25918 4924
rect 25918 4868 25922 4924
rect 25858 4864 25922 4868
rect 25938 4924 26002 4928
rect 25938 4868 25942 4924
rect 25942 4868 25998 4924
rect 25998 4868 26002 4924
rect 25938 4864 26002 4868
rect 26018 4924 26082 4928
rect 26018 4868 26022 4924
rect 26022 4868 26078 4924
rect 26078 4868 26082 4924
rect 26018 4864 26082 4868
rect 28764 4720 28828 4724
rect 28764 4664 28778 4720
rect 28778 4664 28828 4720
rect 28764 4660 28828 4664
rect 10882 4380 10946 4384
rect 10882 4324 10886 4380
rect 10886 4324 10942 4380
rect 10942 4324 10946 4380
rect 10882 4320 10946 4324
rect 10962 4380 11026 4384
rect 10962 4324 10966 4380
rect 10966 4324 11022 4380
rect 11022 4324 11026 4380
rect 10962 4320 11026 4324
rect 11042 4380 11106 4384
rect 11042 4324 11046 4380
rect 11046 4324 11102 4380
rect 11102 4324 11106 4380
rect 11042 4320 11106 4324
rect 11122 4380 11186 4384
rect 11122 4324 11126 4380
rect 11126 4324 11182 4380
rect 11182 4324 11186 4380
rect 11122 4320 11186 4324
rect 20813 4380 20877 4384
rect 20813 4324 20817 4380
rect 20817 4324 20873 4380
rect 20873 4324 20877 4380
rect 20813 4320 20877 4324
rect 20893 4380 20957 4384
rect 20893 4324 20897 4380
rect 20897 4324 20953 4380
rect 20953 4324 20957 4380
rect 20893 4320 20957 4324
rect 20973 4380 21037 4384
rect 20973 4324 20977 4380
rect 20977 4324 21033 4380
rect 21033 4324 21037 4380
rect 20973 4320 21037 4324
rect 21053 4380 21117 4384
rect 21053 4324 21057 4380
rect 21057 4324 21113 4380
rect 21113 4324 21117 4380
rect 21053 4320 21117 4324
rect 29868 4040 29932 4044
rect 29868 3984 29882 4040
rect 29882 3984 29932 4040
rect 29868 3980 29932 3984
rect 5917 3836 5981 3840
rect 5917 3780 5921 3836
rect 5921 3780 5977 3836
rect 5977 3780 5981 3836
rect 5917 3776 5981 3780
rect 5997 3836 6061 3840
rect 5997 3780 6001 3836
rect 6001 3780 6057 3836
rect 6057 3780 6061 3836
rect 5997 3776 6061 3780
rect 6077 3836 6141 3840
rect 6077 3780 6081 3836
rect 6081 3780 6137 3836
rect 6137 3780 6141 3836
rect 6077 3776 6141 3780
rect 6157 3836 6221 3840
rect 6157 3780 6161 3836
rect 6161 3780 6217 3836
rect 6217 3780 6221 3836
rect 6157 3776 6221 3780
rect 15848 3836 15912 3840
rect 15848 3780 15852 3836
rect 15852 3780 15908 3836
rect 15908 3780 15912 3836
rect 15848 3776 15912 3780
rect 15928 3836 15992 3840
rect 15928 3780 15932 3836
rect 15932 3780 15988 3836
rect 15988 3780 15992 3836
rect 15928 3776 15992 3780
rect 16008 3836 16072 3840
rect 16008 3780 16012 3836
rect 16012 3780 16068 3836
rect 16068 3780 16072 3836
rect 16008 3776 16072 3780
rect 16088 3836 16152 3840
rect 16088 3780 16092 3836
rect 16092 3780 16148 3836
rect 16148 3780 16152 3836
rect 16088 3776 16152 3780
rect 25778 3836 25842 3840
rect 25778 3780 25782 3836
rect 25782 3780 25838 3836
rect 25838 3780 25842 3836
rect 25778 3776 25842 3780
rect 25858 3836 25922 3840
rect 25858 3780 25862 3836
rect 25862 3780 25918 3836
rect 25918 3780 25922 3836
rect 25858 3776 25922 3780
rect 25938 3836 26002 3840
rect 25938 3780 25942 3836
rect 25942 3780 25998 3836
rect 25998 3780 26002 3836
rect 25938 3776 26002 3780
rect 26018 3836 26082 3840
rect 26018 3780 26022 3836
rect 26022 3780 26078 3836
rect 26078 3780 26082 3836
rect 26018 3776 26082 3780
rect 10882 3292 10946 3296
rect 10882 3236 10886 3292
rect 10886 3236 10942 3292
rect 10942 3236 10946 3292
rect 10882 3232 10946 3236
rect 10962 3292 11026 3296
rect 10962 3236 10966 3292
rect 10966 3236 11022 3292
rect 11022 3236 11026 3292
rect 10962 3232 11026 3236
rect 11042 3292 11106 3296
rect 11042 3236 11046 3292
rect 11046 3236 11102 3292
rect 11102 3236 11106 3292
rect 11042 3232 11106 3236
rect 11122 3292 11186 3296
rect 11122 3236 11126 3292
rect 11126 3236 11182 3292
rect 11182 3236 11186 3292
rect 11122 3232 11186 3236
rect 20813 3292 20877 3296
rect 20813 3236 20817 3292
rect 20817 3236 20873 3292
rect 20873 3236 20877 3292
rect 20813 3232 20877 3236
rect 20893 3292 20957 3296
rect 20893 3236 20897 3292
rect 20897 3236 20953 3292
rect 20953 3236 20957 3292
rect 20893 3232 20957 3236
rect 20973 3292 21037 3296
rect 20973 3236 20977 3292
rect 20977 3236 21033 3292
rect 21033 3236 21037 3292
rect 20973 3232 21037 3236
rect 21053 3292 21117 3296
rect 21053 3236 21057 3292
rect 21057 3236 21113 3292
rect 21113 3236 21117 3292
rect 21053 3232 21117 3236
rect 5917 2748 5981 2752
rect 5917 2692 5921 2748
rect 5921 2692 5977 2748
rect 5977 2692 5981 2748
rect 5917 2688 5981 2692
rect 5997 2748 6061 2752
rect 5997 2692 6001 2748
rect 6001 2692 6057 2748
rect 6057 2692 6061 2748
rect 5997 2688 6061 2692
rect 6077 2748 6141 2752
rect 6077 2692 6081 2748
rect 6081 2692 6137 2748
rect 6137 2692 6141 2748
rect 6077 2688 6141 2692
rect 6157 2748 6221 2752
rect 6157 2692 6161 2748
rect 6161 2692 6217 2748
rect 6217 2692 6221 2748
rect 6157 2688 6221 2692
rect 15848 2748 15912 2752
rect 15848 2692 15852 2748
rect 15852 2692 15908 2748
rect 15908 2692 15912 2748
rect 15848 2688 15912 2692
rect 15928 2748 15992 2752
rect 15928 2692 15932 2748
rect 15932 2692 15988 2748
rect 15988 2692 15992 2748
rect 15928 2688 15992 2692
rect 16008 2748 16072 2752
rect 16008 2692 16012 2748
rect 16012 2692 16068 2748
rect 16068 2692 16072 2748
rect 16008 2688 16072 2692
rect 16088 2748 16152 2752
rect 16088 2692 16092 2748
rect 16092 2692 16148 2748
rect 16148 2692 16152 2748
rect 16088 2688 16152 2692
rect 25778 2748 25842 2752
rect 25778 2692 25782 2748
rect 25782 2692 25838 2748
rect 25838 2692 25842 2748
rect 25778 2688 25842 2692
rect 25858 2748 25922 2752
rect 25858 2692 25862 2748
rect 25862 2692 25918 2748
rect 25918 2692 25922 2748
rect 25858 2688 25922 2692
rect 25938 2748 26002 2752
rect 25938 2692 25942 2748
rect 25942 2692 25998 2748
rect 25998 2692 26002 2748
rect 25938 2688 26002 2692
rect 26018 2748 26082 2752
rect 26018 2692 26022 2748
rect 26022 2692 26078 2748
rect 26078 2692 26082 2748
rect 26018 2688 26082 2692
rect 10882 2204 10946 2208
rect 10882 2148 10886 2204
rect 10886 2148 10942 2204
rect 10942 2148 10946 2204
rect 10882 2144 10946 2148
rect 10962 2204 11026 2208
rect 10962 2148 10966 2204
rect 10966 2148 11022 2204
rect 11022 2148 11026 2204
rect 10962 2144 11026 2148
rect 11042 2204 11106 2208
rect 11042 2148 11046 2204
rect 11046 2148 11102 2204
rect 11102 2148 11106 2204
rect 11042 2144 11106 2148
rect 11122 2204 11186 2208
rect 11122 2148 11126 2204
rect 11126 2148 11182 2204
rect 11182 2148 11186 2204
rect 11122 2144 11186 2148
rect 20813 2204 20877 2208
rect 20813 2148 20817 2204
rect 20817 2148 20873 2204
rect 20873 2148 20877 2204
rect 20813 2144 20877 2148
rect 20893 2204 20957 2208
rect 20893 2148 20897 2204
rect 20897 2148 20953 2204
rect 20953 2148 20957 2204
rect 20893 2144 20957 2148
rect 20973 2204 21037 2208
rect 20973 2148 20977 2204
rect 20977 2148 21033 2204
rect 21033 2148 21037 2204
rect 20973 2144 21037 2148
rect 21053 2204 21117 2208
rect 21053 2148 21057 2204
rect 21057 2148 21113 2204
rect 21113 2148 21117 2204
rect 21053 2144 21117 2148
<< metal4 >>
rect 5909 77824 6230 77840
rect 5909 77760 5917 77824
rect 5981 77760 5997 77824
rect 6061 77760 6077 77824
rect 6141 77760 6157 77824
rect 6221 77760 6230 77824
rect 5909 76736 6230 77760
rect 5909 76672 5917 76736
rect 5981 76672 5997 76736
rect 6061 76672 6077 76736
rect 6141 76672 6157 76736
rect 6221 76672 6230 76736
rect 5909 75648 6230 76672
rect 5909 75584 5917 75648
rect 5981 75584 5997 75648
rect 6061 75584 6077 75648
rect 6141 75584 6157 75648
rect 6221 75584 6230 75648
rect 5909 74560 6230 75584
rect 5909 74496 5917 74560
rect 5981 74496 5997 74560
rect 6061 74496 6077 74560
rect 6141 74496 6157 74560
rect 6221 74496 6230 74560
rect 5909 73472 6230 74496
rect 5909 73408 5917 73472
rect 5981 73408 5997 73472
rect 6061 73408 6077 73472
rect 6141 73408 6157 73472
rect 6221 73408 6230 73472
rect 5909 72384 6230 73408
rect 5909 72320 5917 72384
rect 5981 72320 5997 72384
rect 6061 72320 6077 72384
rect 6141 72320 6157 72384
rect 6221 72320 6230 72384
rect 5909 71296 6230 72320
rect 5909 71232 5917 71296
rect 5981 71232 5997 71296
rect 6061 71232 6077 71296
rect 6141 71232 6157 71296
rect 6221 71232 6230 71296
rect 5909 70208 6230 71232
rect 5909 70144 5917 70208
rect 5981 70144 5997 70208
rect 6061 70144 6077 70208
rect 6141 70144 6157 70208
rect 6221 70144 6230 70208
rect 5909 69120 6230 70144
rect 5909 69056 5917 69120
rect 5981 69056 5997 69120
rect 6061 69056 6077 69120
rect 6141 69056 6157 69120
rect 6221 69056 6230 69120
rect 5909 68032 6230 69056
rect 5909 67968 5917 68032
rect 5981 67968 5997 68032
rect 6061 67968 6077 68032
rect 6141 67968 6157 68032
rect 6221 67968 6230 68032
rect 5909 66944 6230 67968
rect 5909 66880 5917 66944
rect 5981 66880 5997 66944
rect 6061 66880 6077 66944
rect 6141 66880 6157 66944
rect 6221 66880 6230 66944
rect 5909 65856 6230 66880
rect 5909 65792 5917 65856
rect 5981 65792 5997 65856
rect 6061 65792 6077 65856
rect 6141 65792 6157 65856
rect 6221 65792 6230 65856
rect 5909 64768 6230 65792
rect 5909 64704 5917 64768
rect 5981 64704 5997 64768
rect 6061 64704 6077 64768
rect 6141 64704 6157 64768
rect 6221 64704 6230 64768
rect 5909 63680 6230 64704
rect 5909 63616 5917 63680
rect 5981 63616 5997 63680
rect 6061 63616 6077 63680
rect 6141 63616 6157 63680
rect 6221 63616 6230 63680
rect 5909 62592 6230 63616
rect 5909 62528 5917 62592
rect 5981 62528 5997 62592
rect 6061 62528 6077 62592
rect 6141 62528 6157 62592
rect 6221 62528 6230 62592
rect 5909 61504 6230 62528
rect 5909 61440 5917 61504
rect 5981 61440 5997 61504
rect 6061 61440 6077 61504
rect 6141 61440 6157 61504
rect 6221 61440 6230 61504
rect 5909 60416 6230 61440
rect 5909 60352 5917 60416
rect 5981 60352 5997 60416
rect 6061 60352 6077 60416
rect 6141 60352 6157 60416
rect 6221 60352 6230 60416
rect 5909 59328 6230 60352
rect 5909 59264 5917 59328
rect 5981 59264 5997 59328
rect 6061 59264 6077 59328
rect 6141 59264 6157 59328
rect 6221 59264 6230 59328
rect 5909 58240 6230 59264
rect 5909 58176 5917 58240
rect 5981 58176 5997 58240
rect 6061 58176 6077 58240
rect 6141 58176 6157 58240
rect 6221 58176 6230 58240
rect 5909 57152 6230 58176
rect 5909 57088 5917 57152
rect 5981 57088 5997 57152
rect 6061 57088 6077 57152
rect 6141 57088 6157 57152
rect 6221 57088 6230 57152
rect 5909 56064 6230 57088
rect 5909 56000 5917 56064
rect 5981 56000 5997 56064
rect 6061 56000 6077 56064
rect 6141 56000 6157 56064
rect 6221 56000 6230 56064
rect 5909 54976 6230 56000
rect 5909 54912 5917 54976
rect 5981 54912 5997 54976
rect 6061 54912 6077 54976
rect 6141 54912 6157 54976
rect 6221 54912 6230 54976
rect 5909 53888 6230 54912
rect 5909 53824 5917 53888
rect 5981 53824 5997 53888
rect 6061 53824 6077 53888
rect 6141 53824 6157 53888
rect 6221 53824 6230 53888
rect 5909 52800 6230 53824
rect 5909 52736 5917 52800
rect 5981 52736 5997 52800
rect 6061 52736 6077 52800
rect 6141 52736 6157 52800
rect 6221 52736 6230 52800
rect 5909 51712 6230 52736
rect 5909 51648 5917 51712
rect 5981 51648 5997 51712
rect 6061 51648 6077 51712
rect 6141 51648 6157 51712
rect 6221 51648 6230 51712
rect 5909 50624 6230 51648
rect 5909 50560 5917 50624
rect 5981 50560 5997 50624
rect 6061 50560 6077 50624
rect 6141 50560 6157 50624
rect 6221 50560 6230 50624
rect 5909 49536 6230 50560
rect 5909 49472 5917 49536
rect 5981 49472 5997 49536
rect 6061 49472 6077 49536
rect 6141 49472 6157 49536
rect 6221 49472 6230 49536
rect 5909 48448 6230 49472
rect 5909 48384 5917 48448
rect 5981 48384 5997 48448
rect 6061 48384 6077 48448
rect 6141 48384 6157 48448
rect 6221 48384 6230 48448
rect 5909 47360 6230 48384
rect 5909 47296 5917 47360
rect 5981 47296 5997 47360
rect 6061 47296 6077 47360
rect 6141 47296 6157 47360
rect 6221 47296 6230 47360
rect 5909 46272 6230 47296
rect 5909 46208 5917 46272
rect 5981 46208 5997 46272
rect 6061 46208 6077 46272
rect 6141 46208 6157 46272
rect 6221 46208 6230 46272
rect 5909 45184 6230 46208
rect 5909 45120 5917 45184
rect 5981 45120 5997 45184
rect 6061 45120 6077 45184
rect 6141 45120 6157 45184
rect 6221 45120 6230 45184
rect 5909 44096 6230 45120
rect 5909 44032 5917 44096
rect 5981 44032 5997 44096
rect 6061 44032 6077 44096
rect 6141 44032 6157 44096
rect 6221 44032 6230 44096
rect 5909 43008 6230 44032
rect 5909 42944 5917 43008
rect 5981 42944 5997 43008
rect 6061 42944 6077 43008
rect 6141 42944 6157 43008
rect 6221 42944 6230 43008
rect 5909 41920 6230 42944
rect 5909 41856 5917 41920
rect 5981 41856 5997 41920
rect 6061 41856 6077 41920
rect 6141 41856 6157 41920
rect 6221 41856 6230 41920
rect 5909 40832 6230 41856
rect 5909 40768 5917 40832
rect 5981 40768 5997 40832
rect 6061 40768 6077 40832
rect 6141 40768 6157 40832
rect 6221 40768 6230 40832
rect 5909 39744 6230 40768
rect 5909 39680 5917 39744
rect 5981 39680 5997 39744
rect 6061 39680 6077 39744
rect 6141 39680 6157 39744
rect 6221 39680 6230 39744
rect 5909 38656 6230 39680
rect 5909 38592 5917 38656
rect 5981 38592 5997 38656
rect 6061 38592 6077 38656
rect 6141 38592 6157 38656
rect 6221 38592 6230 38656
rect 5909 37568 6230 38592
rect 5909 37504 5917 37568
rect 5981 37504 5997 37568
rect 6061 37504 6077 37568
rect 6141 37504 6157 37568
rect 6221 37504 6230 37568
rect 5909 36480 6230 37504
rect 5909 36416 5917 36480
rect 5981 36416 5997 36480
rect 6061 36416 6077 36480
rect 6141 36416 6157 36480
rect 6221 36416 6230 36480
rect 5909 35392 6230 36416
rect 5909 35328 5917 35392
rect 5981 35328 5997 35392
rect 6061 35328 6077 35392
rect 6141 35328 6157 35392
rect 6221 35328 6230 35392
rect 5909 34304 6230 35328
rect 5909 34240 5917 34304
rect 5981 34240 5997 34304
rect 6061 34240 6077 34304
rect 6141 34240 6157 34304
rect 6221 34240 6230 34304
rect 5909 33216 6230 34240
rect 5909 33152 5917 33216
rect 5981 33152 5997 33216
rect 6061 33152 6077 33216
rect 6141 33152 6157 33216
rect 6221 33152 6230 33216
rect 5909 32128 6230 33152
rect 5909 32064 5917 32128
rect 5981 32064 5997 32128
rect 6061 32064 6077 32128
rect 6141 32064 6157 32128
rect 6221 32064 6230 32128
rect 5909 31040 6230 32064
rect 5909 30976 5917 31040
rect 5981 30976 5997 31040
rect 6061 30976 6077 31040
rect 6141 30976 6157 31040
rect 6221 30976 6230 31040
rect 5909 29952 6230 30976
rect 5909 29888 5917 29952
rect 5981 29888 5997 29952
rect 6061 29888 6077 29952
rect 6141 29888 6157 29952
rect 6221 29888 6230 29952
rect 5909 28864 6230 29888
rect 5909 28800 5917 28864
rect 5981 28800 5997 28864
rect 6061 28800 6077 28864
rect 6141 28800 6157 28864
rect 6221 28800 6230 28864
rect 5909 27776 6230 28800
rect 5909 27712 5917 27776
rect 5981 27712 5997 27776
rect 6061 27712 6077 27776
rect 6141 27712 6157 27776
rect 6221 27712 6230 27776
rect 5909 26688 6230 27712
rect 5909 26624 5917 26688
rect 5981 26624 5997 26688
rect 6061 26624 6077 26688
rect 6141 26624 6157 26688
rect 6221 26624 6230 26688
rect 5909 25600 6230 26624
rect 5909 25536 5917 25600
rect 5981 25536 5997 25600
rect 6061 25536 6077 25600
rect 6141 25536 6157 25600
rect 6221 25536 6230 25600
rect 5909 24512 6230 25536
rect 5909 24448 5917 24512
rect 5981 24448 5997 24512
rect 6061 24448 6077 24512
rect 6141 24448 6157 24512
rect 6221 24448 6230 24512
rect 5909 23424 6230 24448
rect 5909 23360 5917 23424
rect 5981 23360 5997 23424
rect 6061 23360 6077 23424
rect 6141 23360 6157 23424
rect 6221 23360 6230 23424
rect 5909 22336 6230 23360
rect 5909 22272 5917 22336
rect 5981 22272 5997 22336
rect 6061 22272 6077 22336
rect 6141 22272 6157 22336
rect 6221 22272 6230 22336
rect 5909 21248 6230 22272
rect 5909 21184 5917 21248
rect 5981 21184 5997 21248
rect 6061 21184 6077 21248
rect 6141 21184 6157 21248
rect 6221 21184 6230 21248
rect 5909 20160 6230 21184
rect 5909 20096 5917 20160
rect 5981 20096 5997 20160
rect 6061 20096 6077 20160
rect 6141 20096 6157 20160
rect 6221 20096 6230 20160
rect 5909 19072 6230 20096
rect 5909 19008 5917 19072
rect 5981 19008 5997 19072
rect 6061 19008 6077 19072
rect 6141 19008 6157 19072
rect 6221 19008 6230 19072
rect 5909 17984 6230 19008
rect 5909 17920 5917 17984
rect 5981 17920 5997 17984
rect 6061 17920 6077 17984
rect 6141 17920 6157 17984
rect 6221 17920 6230 17984
rect 5909 16896 6230 17920
rect 5909 16832 5917 16896
rect 5981 16832 5997 16896
rect 6061 16832 6077 16896
rect 6141 16832 6157 16896
rect 6221 16832 6230 16896
rect 5909 15808 6230 16832
rect 5909 15744 5917 15808
rect 5981 15744 5997 15808
rect 6061 15744 6077 15808
rect 6141 15744 6157 15808
rect 6221 15744 6230 15808
rect 5909 14720 6230 15744
rect 5909 14656 5917 14720
rect 5981 14656 5997 14720
rect 6061 14656 6077 14720
rect 6141 14656 6157 14720
rect 6221 14656 6230 14720
rect 5909 13632 6230 14656
rect 5909 13568 5917 13632
rect 5981 13568 5997 13632
rect 6061 13568 6077 13632
rect 6141 13568 6157 13632
rect 6221 13568 6230 13632
rect 5909 12544 6230 13568
rect 5909 12480 5917 12544
rect 5981 12480 5997 12544
rect 6061 12480 6077 12544
rect 6141 12480 6157 12544
rect 6221 12480 6230 12544
rect 5909 11456 6230 12480
rect 5909 11392 5917 11456
rect 5981 11392 5997 11456
rect 6061 11392 6077 11456
rect 6141 11392 6157 11456
rect 6221 11392 6230 11456
rect 5909 10368 6230 11392
rect 5909 10304 5917 10368
rect 5981 10304 5997 10368
rect 6061 10304 6077 10368
rect 6141 10304 6157 10368
rect 6221 10304 6230 10368
rect 5909 9280 6230 10304
rect 5909 9216 5917 9280
rect 5981 9216 5997 9280
rect 6061 9216 6077 9280
rect 6141 9216 6157 9280
rect 6221 9216 6230 9280
rect 5909 8192 6230 9216
rect 5909 8128 5917 8192
rect 5981 8128 5997 8192
rect 6061 8128 6077 8192
rect 6141 8128 6157 8192
rect 6221 8128 6230 8192
rect 5909 7104 6230 8128
rect 5909 7040 5917 7104
rect 5981 7040 5997 7104
rect 6061 7040 6077 7104
rect 6141 7040 6157 7104
rect 6221 7040 6230 7104
rect 5909 6016 6230 7040
rect 5909 5952 5917 6016
rect 5981 5952 5997 6016
rect 6061 5952 6077 6016
rect 6141 5952 6157 6016
rect 6221 5952 6230 6016
rect 5909 4928 6230 5952
rect 5909 4864 5917 4928
rect 5981 4864 5997 4928
rect 6061 4864 6077 4928
rect 6141 4864 6157 4928
rect 6221 4864 6230 4928
rect 5909 3840 6230 4864
rect 5909 3776 5917 3840
rect 5981 3776 5997 3840
rect 6061 3776 6077 3840
rect 6141 3776 6157 3840
rect 6221 3776 6230 3840
rect 5909 2752 6230 3776
rect 5909 2688 5917 2752
rect 5981 2688 5997 2752
rect 6061 2688 6077 2752
rect 6141 2688 6157 2752
rect 6221 2688 6230 2752
rect 5909 2128 6230 2688
rect 10874 77280 11194 77840
rect 10874 77216 10882 77280
rect 10946 77216 10962 77280
rect 11026 77216 11042 77280
rect 11106 77216 11122 77280
rect 11186 77216 11194 77280
rect 10874 76192 11194 77216
rect 10874 76128 10882 76192
rect 10946 76128 10962 76192
rect 11026 76128 11042 76192
rect 11106 76128 11122 76192
rect 11186 76128 11194 76192
rect 10874 75104 11194 76128
rect 10874 75040 10882 75104
rect 10946 75040 10962 75104
rect 11026 75040 11042 75104
rect 11106 75040 11122 75104
rect 11186 75040 11194 75104
rect 10874 74016 11194 75040
rect 10874 73952 10882 74016
rect 10946 73952 10962 74016
rect 11026 73952 11042 74016
rect 11106 73952 11122 74016
rect 11186 73952 11194 74016
rect 10874 72928 11194 73952
rect 10874 72864 10882 72928
rect 10946 72864 10962 72928
rect 11026 72864 11042 72928
rect 11106 72864 11122 72928
rect 11186 72864 11194 72928
rect 10874 71840 11194 72864
rect 10874 71776 10882 71840
rect 10946 71776 10962 71840
rect 11026 71776 11042 71840
rect 11106 71776 11122 71840
rect 11186 71776 11194 71840
rect 10874 70752 11194 71776
rect 10874 70688 10882 70752
rect 10946 70688 10962 70752
rect 11026 70688 11042 70752
rect 11106 70688 11122 70752
rect 11186 70688 11194 70752
rect 10874 69664 11194 70688
rect 10874 69600 10882 69664
rect 10946 69600 10962 69664
rect 11026 69600 11042 69664
rect 11106 69600 11122 69664
rect 11186 69600 11194 69664
rect 10874 68576 11194 69600
rect 10874 68512 10882 68576
rect 10946 68512 10962 68576
rect 11026 68512 11042 68576
rect 11106 68512 11122 68576
rect 11186 68512 11194 68576
rect 10874 67488 11194 68512
rect 10874 67424 10882 67488
rect 10946 67424 10962 67488
rect 11026 67424 11042 67488
rect 11106 67424 11122 67488
rect 11186 67424 11194 67488
rect 10874 66400 11194 67424
rect 10874 66336 10882 66400
rect 10946 66336 10962 66400
rect 11026 66336 11042 66400
rect 11106 66336 11122 66400
rect 11186 66336 11194 66400
rect 10874 65312 11194 66336
rect 10874 65248 10882 65312
rect 10946 65248 10962 65312
rect 11026 65248 11042 65312
rect 11106 65248 11122 65312
rect 11186 65248 11194 65312
rect 10874 64224 11194 65248
rect 10874 64160 10882 64224
rect 10946 64160 10962 64224
rect 11026 64160 11042 64224
rect 11106 64160 11122 64224
rect 11186 64160 11194 64224
rect 10874 63136 11194 64160
rect 10874 63072 10882 63136
rect 10946 63072 10962 63136
rect 11026 63072 11042 63136
rect 11106 63072 11122 63136
rect 11186 63072 11194 63136
rect 10874 62048 11194 63072
rect 10874 61984 10882 62048
rect 10946 61984 10962 62048
rect 11026 61984 11042 62048
rect 11106 61984 11122 62048
rect 11186 61984 11194 62048
rect 10874 60960 11194 61984
rect 10874 60896 10882 60960
rect 10946 60896 10962 60960
rect 11026 60896 11042 60960
rect 11106 60896 11122 60960
rect 11186 60896 11194 60960
rect 10874 59872 11194 60896
rect 10874 59808 10882 59872
rect 10946 59808 10962 59872
rect 11026 59808 11042 59872
rect 11106 59808 11122 59872
rect 11186 59808 11194 59872
rect 10874 58784 11194 59808
rect 10874 58720 10882 58784
rect 10946 58720 10962 58784
rect 11026 58720 11042 58784
rect 11106 58720 11122 58784
rect 11186 58720 11194 58784
rect 10874 57696 11194 58720
rect 10874 57632 10882 57696
rect 10946 57632 10962 57696
rect 11026 57632 11042 57696
rect 11106 57632 11122 57696
rect 11186 57632 11194 57696
rect 10874 56608 11194 57632
rect 10874 56544 10882 56608
rect 10946 56544 10962 56608
rect 11026 56544 11042 56608
rect 11106 56544 11122 56608
rect 11186 56544 11194 56608
rect 10874 55520 11194 56544
rect 10874 55456 10882 55520
rect 10946 55456 10962 55520
rect 11026 55456 11042 55520
rect 11106 55456 11122 55520
rect 11186 55456 11194 55520
rect 10874 54432 11194 55456
rect 10874 54368 10882 54432
rect 10946 54368 10962 54432
rect 11026 54368 11042 54432
rect 11106 54368 11122 54432
rect 11186 54368 11194 54432
rect 10874 53344 11194 54368
rect 10874 53280 10882 53344
rect 10946 53280 10962 53344
rect 11026 53280 11042 53344
rect 11106 53280 11122 53344
rect 11186 53280 11194 53344
rect 10874 52256 11194 53280
rect 10874 52192 10882 52256
rect 10946 52192 10962 52256
rect 11026 52192 11042 52256
rect 11106 52192 11122 52256
rect 11186 52192 11194 52256
rect 10874 51168 11194 52192
rect 10874 51104 10882 51168
rect 10946 51104 10962 51168
rect 11026 51104 11042 51168
rect 11106 51104 11122 51168
rect 11186 51104 11194 51168
rect 10874 50080 11194 51104
rect 10874 50016 10882 50080
rect 10946 50016 10962 50080
rect 11026 50016 11042 50080
rect 11106 50016 11122 50080
rect 11186 50016 11194 50080
rect 10874 48992 11194 50016
rect 10874 48928 10882 48992
rect 10946 48928 10962 48992
rect 11026 48928 11042 48992
rect 11106 48928 11122 48992
rect 11186 48928 11194 48992
rect 10874 47904 11194 48928
rect 10874 47840 10882 47904
rect 10946 47840 10962 47904
rect 11026 47840 11042 47904
rect 11106 47840 11122 47904
rect 11186 47840 11194 47904
rect 10874 46816 11194 47840
rect 10874 46752 10882 46816
rect 10946 46752 10962 46816
rect 11026 46752 11042 46816
rect 11106 46752 11122 46816
rect 11186 46752 11194 46816
rect 10874 45728 11194 46752
rect 10874 45664 10882 45728
rect 10946 45664 10962 45728
rect 11026 45664 11042 45728
rect 11106 45664 11122 45728
rect 11186 45664 11194 45728
rect 10874 44640 11194 45664
rect 10874 44576 10882 44640
rect 10946 44576 10962 44640
rect 11026 44576 11042 44640
rect 11106 44576 11122 44640
rect 11186 44576 11194 44640
rect 10874 43552 11194 44576
rect 10874 43488 10882 43552
rect 10946 43488 10962 43552
rect 11026 43488 11042 43552
rect 11106 43488 11122 43552
rect 11186 43488 11194 43552
rect 10874 42464 11194 43488
rect 10874 42400 10882 42464
rect 10946 42400 10962 42464
rect 11026 42400 11042 42464
rect 11106 42400 11122 42464
rect 11186 42400 11194 42464
rect 10874 41376 11194 42400
rect 10874 41312 10882 41376
rect 10946 41312 10962 41376
rect 11026 41312 11042 41376
rect 11106 41312 11122 41376
rect 11186 41312 11194 41376
rect 10874 40288 11194 41312
rect 10874 40224 10882 40288
rect 10946 40224 10962 40288
rect 11026 40224 11042 40288
rect 11106 40224 11122 40288
rect 11186 40224 11194 40288
rect 10874 39200 11194 40224
rect 10874 39136 10882 39200
rect 10946 39136 10962 39200
rect 11026 39136 11042 39200
rect 11106 39136 11122 39200
rect 11186 39136 11194 39200
rect 10874 38112 11194 39136
rect 10874 38048 10882 38112
rect 10946 38048 10962 38112
rect 11026 38048 11042 38112
rect 11106 38048 11122 38112
rect 11186 38048 11194 38112
rect 10874 37024 11194 38048
rect 10874 36960 10882 37024
rect 10946 36960 10962 37024
rect 11026 36960 11042 37024
rect 11106 36960 11122 37024
rect 11186 36960 11194 37024
rect 10874 35936 11194 36960
rect 10874 35872 10882 35936
rect 10946 35872 10962 35936
rect 11026 35872 11042 35936
rect 11106 35872 11122 35936
rect 11186 35872 11194 35936
rect 10874 34848 11194 35872
rect 10874 34784 10882 34848
rect 10946 34784 10962 34848
rect 11026 34784 11042 34848
rect 11106 34784 11122 34848
rect 11186 34784 11194 34848
rect 10874 33760 11194 34784
rect 10874 33696 10882 33760
rect 10946 33696 10962 33760
rect 11026 33696 11042 33760
rect 11106 33696 11122 33760
rect 11186 33696 11194 33760
rect 10874 32672 11194 33696
rect 10874 32608 10882 32672
rect 10946 32608 10962 32672
rect 11026 32608 11042 32672
rect 11106 32608 11122 32672
rect 11186 32608 11194 32672
rect 10874 31584 11194 32608
rect 10874 31520 10882 31584
rect 10946 31520 10962 31584
rect 11026 31520 11042 31584
rect 11106 31520 11122 31584
rect 11186 31520 11194 31584
rect 10874 30496 11194 31520
rect 10874 30432 10882 30496
rect 10946 30432 10962 30496
rect 11026 30432 11042 30496
rect 11106 30432 11122 30496
rect 11186 30432 11194 30496
rect 10874 29408 11194 30432
rect 10874 29344 10882 29408
rect 10946 29344 10962 29408
rect 11026 29344 11042 29408
rect 11106 29344 11122 29408
rect 11186 29344 11194 29408
rect 10874 28320 11194 29344
rect 10874 28256 10882 28320
rect 10946 28256 10962 28320
rect 11026 28256 11042 28320
rect 11106 28256 11122 28320
rect 11186 28256 11194 28320
rect 10874 27232 11194 28256
rect 15840 77824 16160 77840
rect 15840 77760 15848 77824
rect 15912 77760 15928 77824
rect 15992 77760 16008 77824
rect 16072 77760 16088 77824
rect 16152 77760 16160 77824
rect 15840 76736 16160 77760
rect 15840 76672 15848 76736
rect 15912 76672 15928 76736
rect 15992 76672 16008 76736
rect 16072 76672 16088 76736
rect 16152 76672 16160 76736
rect 15840 75648 16160 76672
rect 15840 75584 15848 75648
rect 15912 75584 15928 75648
rect 15992 75584 16008 75648
rect 16072 75584 16088 75648
rect 16152 75584 16160 75648
rect 15840 74560 16160 75584
rect 15840 74496 15848 74560
rect 15912 74496 15928 74560
rect 15992 74496 16008 74560
rect 16072 74496 16088 74560
rect 16152 74496 16160 74560
rect 15840 73472 16160 74496
rect 15840 73408 15848 73472
rect 15912 73408 15928 73472
rect 15992 73408 16008 73472
rect 16072 73408 16088 73472
rect 16152 73408 16160 73472
rect 15840 72384 16160 73408
rect 15840 72320 15848 72384
rect 15912 72320 15928 72384
rect 15992 72320 16008 72384
rect 16072 72320 16088 72384
rect 16152 72320 16160 72384
rect 15840 71296 16160 72320
rect 15840 71232 15848 71296
rect 15912 71232 15928 71296
rect 15992 71232 16008 71296
rect 16072 71232 16088 71296
rect 16152 71232 16160 71296
rect 15840 70208 16160 71232
rect 15840 70144 15848 70208
rect 15912 70144 15928 70208
rect 15992 70144 16008 70208
rect 16072 70144 16088 70208
rect 16152 70144 16160 70208
rect 15840 69120 16160 70144
rect 15840 69056 15848 69120
rect 15912 69056 15928 69120
rect 15992 69056 16008 69120
rect 16072 69056 16088 69120
rect 16152 69056 16160 69120
rect 15840 68032 16160 69056
rect 15840 67968 15848 68032
rect 15912 67968 15928 68032
rect 15992 67968 16008 68032
rect 16072 67968 16088 68032
rect 16152 67968 16160 68032
rect 15840 66944 16160 67968
rect 15840 66880 15848 66944
rect 15912 66880 15928 66944
rect 15992 66880 16008 66944
rect 16072 66880 16088 66944
rect 16152 66880 16160 66944
rect 15840 65856 16160 66880
rect 15840 65792 15848 65856
rect 15912 65792 15928 65856
rect 15992 65792 16008 65856
rect 16072 65792 16088 65856
rect 16152 65792 16160 65856
rect 15840 64768 16160 65792
rect 15840 64704 15848 64768
rect 15912 64704 15928 64768
rect 15992 64704 16008 64768
rect 16072 64704 16088 64768
rect 16152 64704 16160 64768
rect 15840 63680 16160 64704
rect 15840 63616 15848 63680
rect 15912 63616 15928 63680
rect 15992 63616 16008 63680
rect 16072 63616 16088 63680
rect 16152 63616 16160 63680
rect 15840 62592 16160 63616
rect 15840 62528 15848 62592
rect 15912 62528 15928 62592
rect 15992 62528 16008 62592
rect 16072 62528 16088 62592
rect 16152 62528 16160 62592
rect 15840 61504 16160 62528
rect 15840 61440 15848 61504
rect 15912 61440 15928 61504
rect 15992 61440 16008 61504
rect 16072 61440 16088 61504
rect 16152 61440 16160 61504
rect 15840 60416 16160 61440
rect 15840 60352 15848 60416
rect 15912 60352 15928 60416
rect 15992 60352 16008 60416
rect 16072 60352 16088 60416
rect 16152 60352 16160 60416
rect 15840 59328 16160 60352
rect 15840 59264 15848 59328
rect 15912 59264 15928 59328
rect 15992 59264 16008 59328
rect 16072 59264 16088 59328
rect 16152 59264 16160 59328
rect 15840 58240 16160 59264
rect 15840 58176 15848 58240
rect 15912 58176 15928 58240
rect 15992 58176 16008 58240
rect 16072 58176 16088 58240
rect 16152 58176 16160 58240
rect 15840 57152 16160 58176
rect 15840 57088 15848 57152
rect 15912 57088 15928 57152
rect 15992 57088 16008 57152
rect 16072 57088 16088 57152
rect 16152 57088 16160 57152
rect 15840 56064 16160 57088
rect 20805 77280 21125 77840
rect 20805 77216 20813 77280
rect 20877 77216 20893 77280
rect 20957 77216 20973 77280
rect 21037 77216 21053 77280
rect 21117 77216 21125 77280
rect 20805 76192 21125 77216
rect 20805 76128 20813 76192
rect 20877 76128 20893 76192
rect 20957 76128 20973 76192
rect 21037 76128 21053 76192
rect 21117 76128 21125 76192
rect 20805 75104 21125 76128
rect 20805 75040 20813 75104
rect 20877 75040 20893 75104
rect 20957 75040 20973 75104
rect 21037 75040 21053 75104
rect 21117 75040 21125 75104
rect 20805 74016 21125 75040
rect 20805 73952 20813 74016
rect 20877 73952 20893 74016
rect 20957 73952 20973 74016
rect 21037 73952 21053 74016
rect 21117 73952 21125 74016
rect 20805 72928 21125 73952
rect 20805 72864 20813 72928
rect 20877 72864 20893 72928
rect 20957 72864 20973 72928
rect 21037 72864 21053 72928
rect 21117 72864 21125 72928
rect 20805 71840 21125 72864
rect 20805 71776 20813 71840
rect 20877 71776 20893 71840
rect 20957 71776 20973 71840
rect 21037 71776 21053 71840
rect 21117 71776 21125 71840
rect 20805 70752 21125 71776
rect 20805 70688 20813 70752
rect 20877 70688 20893 70752
rect 20957 70688 20973 70752
rect 21037 70688 21053 70752
rect 21117 70688 21125 70752
rect 20805 69664 21125 70688
rect 20805 69600 20813 69664
rect 20877 69600 20893 69664
rect 20957 69600 20973 69664
rect 21037 69600 21053 69664
rect 21117 69600 21125 69664
rect 20805 68576 21125 69600
rect 20805 68512 20813 68576
rect 20877 68512 20893 68576
rect 20957 68512 20973 68576
rect 21037 68512 21053 68576
rect 21117 68512 21125 68576
rect 20805 67488 21125 68512
rect 20805 67424 20813 67488
rect 20877 67424 20893 67488
rect 20957 67424 20973 67488
rect 21037 67424 21053 67488
rect 21117 67424 21125 67488
rect 20805 66400 21125 67424
rect 20805 66336 20813 66400
rect 20877 66336 20893 66400
rect 20957 66336 20973 66400
rect 21037 66336 21053 66400
rect 21117 66336 21125 66400
rect 20805 65312 21125 66336
rect 25770 77824 26091 77840
rect 25770 77760 25778 77824
rect 25842 77760 25858 77824
rect 25922 77760 25938 77824
rect 26002 77760 26018 77824
rect 26082 77760 26091 77824
rect 25770 76736 26091 77760
rect 25770 76672 25778 76736
rect 25842 76672 25858 76736
rect 25922 76672 25938 76736
rect 26002 76672 26018 76736
rect 26082 76672 26091 76736
rect 25770 75648 26091 76672
rect 25770 75584 25778 75648
rect 25842 75584 25858 75648
rect 25922 75584 25938 75648
rect 26002 75584 26018 75648
rect 26082 75584 26091 75648
rect 25770 74560 26091 75584
rect 25770 74496 25778 74560
rect 25842 74496 25858 74560
rect 25922 74496 25938 74560
rect 26002 74496 26018 74560
rect 26082 74496 26091 74560
rect 25770 73472 26091 74496
rect 25770 73408 25778 73472
rect 25842 73408 25858 73472
rect 25922 73408 25938 73472
rect 26002 73408 26018 73472
rect 26082 73408 26091 73472
rect 25770 72384 26091 73408
rect 25770 72320 25778 72384
rect 25842 72320 25858 72384
rect 25922 72320 25938 72384
rect 26002 72320 26018 72384
rect 26082 72320 26091 72384
rect 25770 71296 26091 72320
rect 25770 71232 25778 71296
rect 25842 71232 25858 71296
rect 25922 71232 25938 71296
rect 26002 71232 26018 71296
rect 26082 71232 26091 71296
rect 25770 70208 26091 71232
rect 25770 70144 25778 70208
rect 25842 70144 25858 70208
rect 25922 70144 25938 70208
rect 26002 70144 26018 70208
rect 26082 70144 26091 70208
rect 25770 69120 26091 70144
rect 29131 70004 29197 70005
rect 29131 69940 29132 70004
rect 29196 69940 29197 70004
rect 29131 69939 29197 69940
rect 25770 69056 25778 69120
rect 25842 69056 25858 69120
rect 25922 69056 25938 69120
rect 26002 69056 26018 69120
rect 26082 69056 26091 69120
rect 25770 68032 26091 69056
rect 25770 67968 25778 68032
rect 25842 67968 25858 68032
rect 25922 67968 25938 68032
rect 26002 67968 26018 68032
rect 26082 67968 26091 68032
rect 25770 66944 26091 67968
rect 27107 67556 27173 67557
rect 27107 67492 27108 67556
rect 27172 67492 27173 67556
rect 27107 67491 27173 67492
rect 25770 66880 25778 66944
rect 25842 66880 25858 66944
rect 25922 66880 25938 66944
rect 26002 66880 26018 66944
rect 26082 66880 26091 66944
rect 25083 66060 25149 66061
rect 25083 65996 25084 66060
rect 25148 65996 25149 66060
rect 25083 65995 25149 65996
rect 20805 65248 20813 65312
rect 20877 65248 20893 65312
rect 20957 65248 20973 65312
rect 21037 65248 21053 65312
rect 21117 65248 21125 65312
rect 20805 64224 21125 65248
rect 20805 64160 20813 64224
rect 20877 64160 20893 64224
rect 20957 64160 20973 64224
rect 21037 64160 21053 64224
rect 21117 64160 21125 64224
rect 20805 63136 21125 64160
rect 20805 63072 20813 63136
rect 20877 63072 20893 63136
rect 20957 63072 20973 63136
rect 21037 63072 21053 63136
rect 21117 63072 21125 63136
rect 20805 62048 21125 63072
rect 20805 61984 20813 62048
rect 20877 61984 20893 62048
rect 20957 61984 20973 62048
rect 21037 61984 21053 62048
rect 21117 61984 21125 62048
rect 20805 60960 21125 61984
rect 20805 60896 20813 60960
rect 20877 60896 20893 60960
rect 20957 60896 20973 60960
rect 21037 60896 21053 60960
rect 21117 60896 21125 60960
rect 20805 59872 21125 60896
rect 20805 59808 20813 59872
rect 20877 59808 20893 59872
rect 20957 59808 20973 59872
rect 21037 59808 21053 59872
rect 21117 59808 21125 59872
rect 20805 58784 21125 59808
rect 20805 58720 20813 58784
rect 20877 58720 20893 58784
rect 20957 58720 20973 58784
rect 21037 58720 21053 58784
rect 21117 58720 21125 58784
rect 20805 57696 21125 58720
rect 20805 57632 20813 57696
rect 20877 57632 20893 57696
rect 20957 57632 20973 57696
rect 21037 57632 21053 57696
rect 21117 57632 21125 57696
rect 17355 56812 17421 56813
rect 17355 56748 17356 56812
rect 17420 56748 17421 56812
rect 17355 56747 17421 56748
rect 15840 56000 15848 56064
rect 15912 56000 15928 56064
rect 15992 56000 16008 56064
rect 16072 56000 16088 56064
rect 16152 56000 16160 56064
rect 15840 54976 16160 56000
rect 15840 54912 15848 54976
rect 15912 54912 15928 54976
rect 15992 54912 16008 54976
rect 16072 54912 16088 54976
rect 16152 54912 16160 54976
rect 15840 53888 16160 54912
rect 15840 53824 15848 53888
rect 15912 53824 15928 53888
rect 15992 53824 16008 53888
rect 16072 53824 16088 53888
rect 16152 53824 16160 53888
rect 15840 52800 16160 53824
rect 15840 52736 15848 52800
rect 15912 52736 15928 52800
rect 15992 52736 16008 52800
rect 16072 52736 16088 52800
rect 16152 52736 16160 52800
rect 15840 51712 16160 52736
rect 15840 51648 15848 51712
rect 15912 51648 15928 51712
rect 15992 51648 16008 51712
rect 16072 51648 16088 51712
rect 16152 51648 16160 51712
rect 15840 50624 16160 51648
rect 15840 50560 15848 50624
rect 15912 50560 15928 50624
rect 15992 50560 16008 50624
rect 16072 50560 16088 50624
rect 16152 50560 16160 50624
rect 15840 49536 16160 50560
rect 15840 49472 15848 49536
rect 15912 49472 15928 49536
rect 15992 49472 16008 49536
rect 16072 49472 16088 49536
rect 16152 49472 16160 49536
rect 15840 48448 16160 49472
rect 15840 48384 15848 48448
rect 15912 48384 15928 48448
rect 15992 48384 16008 48448
rect 16072 48384 16088 48448
rect 16152 48384 16160 48448
rect 15840 47360 16160 48384
rect 15840 47296 15848 47360
rect 15912 47296 15928 47360
rect 15992 47296 16008 47360
rect 16072 47296 16088 47360
rect 16152 47296 16160 47360
rect 15840 46272 16160 47296
rect 15840 46208 15848 46272
rect 15912 46208 15928 46272
rect 15992 46208 16008 46272
rect 16072 46208 16088 46272
rect 16152 46208 16160 46272
rect 15840 45184 16160 46208
rect 15840 45120 15848 45184
rect 15912 45120 15928 45184
rect 15992 45120 16008 45184
rect 16072 45120 16088 45184
rect 16152 45120 16160 45184
rect 15840 44096 16160 45120
rect 15840 44032 15848 44096
rect 15912 44032 15928 44096
rect 15992 44032 16008 44096
rect 16072 44032 16088 44096
rect 16152 44032 16160 44096
rect 15840 43008 16160 44032
rect 15840 42944 15848 43008
rect 15912 42944 15928 43008
rect 15992 42944 16008 43008
rect 16072 42944 16088 43008
rect 16152 42944 16160 43008
rect 15840 41920 16160 42944
rect 15840 41856 15848 41920
rect 15912 41856 15928 41920
rect 15992 41856 16008 41920
rect 16072 41856 16088 41920
rect 16152 41856 16160 41920
rect 15840 40832 16160 41856
rect 15840 40768 15848 40832
rect 15912 40768 15928 40832
rect 15992 40768 16008 40832
rect 16072 40768 16088 40832
rect 16152 40768 16160 40832
rect 15840 39744 16160 40768
rect 15840 39680 15848 39744
rect 15912 39680 15928 39744
rect 15992 39680 16008 39744
rect 16072 39680 16088 39744
rect 16152 39680 16160 39744
rect 15840 38656 16160 39680
rect 15840 38592 15848 38656
rect 15912 38592 15928 38656
rect 15992 38592 16008 38656
rect 16072 38592 16088 38656
rect 16152 38592 16160 38656
rect 15840 37568 16160 38592
rect 15840 37504 15848 37568
rect 15912 37504 15928 37568
rect 15992 37504 16008 37568
rect 16072 37504 16088 37568
rect 16152 37504 16160 37568
rect 15840 36480 16160 37504
rect 15840 36416 15848 36480
rect 15912 36416 15928 36480
rect 15992 36416 16008 36480
rect 16072 36416 16088 36480
rect 16152 36416 16160 36480
rect 15840 35392 16160 36416
rect 15840 35328 15848 35392
rect 15912 35328 15928 35392
rect 15992 35328 16008 35392
rect 16072 35328 16088 35392
rect 16152 35328 16160 35392
rect 15840 34304 16160 35328
rect 15840 34240 15848 34304
rect 15912 34240 15928 34304
rect 15992 34240 16008 34304
rect 16072 34240 16088 34304
rect 16152 34240 16160 34304
rect 15840 33216 16160 34240
rect 17358 34101 17418 56747
rect 20805 56608 21125 57632
rect 23979 57356 24045 57357
rect 23979 57292 23980 57356
rect 24044 57292 24045 57356
rect 23979 57291 24045 57292
rect 23427 56948 23493 56949
rect 23427 56884 23428 56948
rect 23492 56884 23493 56948
rect 23427 56883 23493 56884
rect 20805 56544 20813 56608
rect 20877 56544 20893 56608
rect 20957 56544 20973 56608
rect 21037 56544 21053 56608
rect 21117 56544 21125 56608
rect 20805 55520 21125 56544
rect 20805 55456 20813 55520
rect 20877 55456 20893 55520
rect 20957 55456 20973 55520
rect 21037 55456 21053 55520
rect 21117 55456 21125 55520
rect 20805 54432 21125 55456
rect 20805 54368 20813 54432
rect 20877 54368 20893 54432
rect 20957 54368 20973 54432
rect 21037 54368 21053 54432
rect 21117 54368 21125 54432
rect 19195 53820 19261 53821
rect 19195 53756 19196 53820
rect 19260 53756 19261 53820
rect 19195 53755 19261 53756
rect 17539 53684 17605 53685
rect 17539 53620 17540 53684
rect 17604 53620 17605 53684
rect 17539 53619 17605 53620
rect 17355 34100 17421 34101
rect 17355 34036 17356 34100
rect 17420 34036 17421 34100
rect 17355 34035 17421 34036
rect 15840 33152 15848 33216
rect 15912 33152 15928 33216
rect 15992 33152 16008 33216
rect 16072 33152 16088 33216
rect 16152 33152 16160 33216
rect 15840 32128 16160 33152
rect 15840 32064 15848 32128
rect 15912 32064 15928 32128
rect 15992 32064 16008 32128
rect 16072 32064 16088 32128
rect 16152 32064 16160 32128
rect 15840 31040 16160 32064
rect 15840 30976 15848 31040
rect 15912 30976 15928 31040
rect 15992 30976 16008 31040
rect 16072 30976 16088 31040
rect 16152 30976 16160 31040
rect 15840 29952 16160 30976
rect 15840 29888 15848 29952
rect 15912 29888 15928 29952
rect 15992 29888 16008 29952
rect 16072 29888 16088 29952
rect 16152 29888 16160 29952
rect 15840 28864 16160 29888
rect 15840 28800 15848 28864
rect 15912 28800 15928 28864
rect 15992 28800 16008 28864
rect 16072 28800 16088 28864
rect 16152 28800 16160 28864
rect 15515 28252 15581 28253
rect 15515 28188 15516 28252
rect 15580 28188 15581 28252
rect 15515 28187 15581 28188
rect 15518 27845 15578 28187
rect 15515 27844 15581 27845
rect 15515 27780 15516 27844
rect 15580 27780 15581 27844
rect 15515 27779 15581 27780
rect 10874 27168 10882 27232
rect 10946 27168 10962 27232
rect 11026 27168 11042 27232
rect 11106 27168 11122 27232
rect 11186 27168 11194 27232
rect 10874 26144 11194 27168
rect 10874 26080 10882 26144
rect 10946 26080 10962 26144
rect 11026 26080 11042 26144
rect 11106 26080 11122 26144
rect 11186 26080 11194 26144
rect 10874 25056 11194 26080
rect 10874 24992 10882 25056
rect 10946 24992 10962 25056
rect 11026 24992 11042 25056
rect 11106 24992 11122 25056
rect 11186 24992 11194 25056
rect 10874 23968 11194 24992
rect 10874 23904 10882 23968
rect 10946 23904 10962 23968
rect 11026 23904 11042 23968
rect 11106 23904 11122 23968
rect 11186 23904 11194 23968
rect 10874 22880 11194 23904
rect 10874 22816 10882 22880
rect 10946 22816 10962 22880
rect 11026 22816 11042 22880
rect 11106 22816 11122 22880
rect 11186 22816 11194 22880
rect 10874 21792 11194 22816
rect 10874 21728 10882 21792
rect 10946 21728 10962 21792
rect 11026 21728 11042 21792
rect 11106 21728 11122 21792
rect 11186 21728 11194 21792
rect 10874 20704 11194 21728
rect 10874 20640 10882 20704
rect 10946 20640 10962 20704
rect 11026 20640 11042 20704
rect 11106 20640 11122 20704
rect 11186 20640 11194 20704
rect 10874 19616 11194 20640
rect 10874 19552 10882 19616
rect 10946 19552 10962 19616
rect 11026 19552 11042 19616
rect 11106 19552 11122 19616
rect 11186 19552 11194 19616
rect 10874 18528 11194 19552
rect 10874 18464 10882 18528
rect 10946 18464 10962 18528
rect 11026 18464 11042 18528
rect 11106 18464 11122 18528
rect 11186 18464 11194 18528
rect 10874 17440 11194 18464
rect 10874 17376 10882 17440
rect 10946 17376 10962 17440
rect 11026 17376 11042 17440
rect 11106 17376 11122 17440
rect 11186 17376 11194 17440
rect 10874 16352 11194 17376
rect 10874 16288 10882 16352
rect 10946 16288 10962 16352
rect 11026 16288 11042 16352
rect 11106 16288 11122 16352
rect 11186 16288 11194 16352
rect 10874 15264 11194 16288
rect 10874 15200 10882 15264
rect 10946 15200 10962 15264
rect 11026 15200 11042 15264
rect 11106 15200 11122 15264
rect 11186 15200 11194 15264
rect 10874 14176 11194 15200
rect 10874 14112 10882 14176
rect 10946 14112 10962 14176
rect 11026 14112 11042 14176
rect 11106 14112 11122 14176
rect 11186 14112 11194 14176
rect 10874 13088 11194 14112
rect 10874 13024 10882 13088
rect 10946 13024 10962 13088
rect 11026 13024 11042 13088
rect 11106 13024 11122 13088
rect 11186 13024 11194 13088
rect 10874 12000 11194 13024
rect 10874 11936 10882 12000
rect 10946 11936 10962 12000
rect 11026 11936 11042 12000
rect 11106 11936 11122 12000
rect 11186 11936 11194 12000
rect 10874 10912 11194 11936
rect 10874 10848 10882 10912
rect 10946 10848 10962 10912
rect 11026 10848 11042 10912
rect 11106 10848 11122 10912
rect 11186 10848 11194 10912
rect 10874 9824 11194 10848
rect 10874 9760 10882 9824
rect 10946 9760 10962 9824
rect 11026 9760 11042 9824
rect 11106 9760 11122 9824
rect 11186 9760 11194 9824
rect 10874 8736 11194 9760
rect 10874 8672 10882 8736
rect 10946 8672 10962 8736
rect 11026 8672 11042 8736
rect 11106 8672 11122 8736
rect 11186 8672 11194 8736
rect 10874 7648 11194 8672
rect 10874 7584 10882 7648
rect 10946 7584 10962 7648
rect 11026 7584 11042 7648
rect 11106 7584 11122 7648
rect 11186 7584 11194 7648
rect 10874 6560 11194 7584
rect 10874 6496 10882 6560
rect 10946 6496 10962 6560
rect 11026 6496 11042 6560
rect 11106 6496 11122 6560
rect 11186 6496 11194 6560
rect 10874 5472 11194 6496
rect 10874 5408 10882 5472
rect 10946 5408 10962 5472
rect 11026 5408 11042 5472
rect 11106 5408 11122 5472
rect 11186 5408 11194 5472
rect 10874 4384 11194 5408
rect 10874 4320 10882 4384
rect 10946 4320 10962 4384
rect 11026 4320 11042 4384
rect 11106 4320 11122 4384
rect 11186 4320 11194 4384
rect 10874 3296 11194 4320
rect 10874 3232 10882 3296
rect 10946 3232 10962 3296
rect 11026 3232 11042 3296
rect 11106 3232 11122 3296
rect 11186 3232 11194 3296
rect 10874 2208 11194 3232
rect 10874 2144 10882 2208
rect 10946 2144 10962 2208
rect 11026 2144 11042 2208
rect 11106 2144 11122 2208
rect 11186 2144 11194 2208
rect 10874 2128 11194 2144
rect 15840 27776 16160 28800
rect 15840 27712 15848 27776
rect 15912 27712 15928 27776
rect 15992 27712 16008 27776
rect 16072 27712 16088 27776
rect 16152 27712 16160 27776
rect 15840 26688 16160 27712
rect 17542 27573 17602 53619
rect 17723 50828 17789 50829
rect 17723 50764 17724 50828
rect 17788 50764 17789 50828
rect 17723 50763 17789 50764
rect 17539 27572 17605 27573
rect 17539 27508 17540 27572
rect 17604 27508 17605 27572
rect 17539 27507 17605 27508
rect 15840 26624 15848 26688
rect 15912 26624 15928 26688
rect 15992 26624 16008 26688
rect 16072 26624 16088 26688
rect 16152 26624 16160 26688
rect 15840 25600 16160 26624
rect 15840 25536 15848 25600
rect 15912 25536 15928 25600
rect 15992 25536 16008 25600
rect 16072 25536 16088 25600
rect 16152 25536 16160 25600
rect 15840 24512 16160 25536
rect 15840 24448 15848 24512
rect 15912 24448 15928 24512
rect 15992 24448 16008 24512
rect 16072 24448 16088 24512
rect 16152 24448 16160 24512
rect 15840 23424 16160 24448
rect 15840 23360 15848 23424
rect 15912 23360 15928 23424
rect 15992 23360 16008 23424
rect 16072 23360 16088 23424
rect 16152 23360 16160 23424
rect 15840 22336 16160 23360
rect 15840 22272 15848 22336
rect 15912 22272 15928 22336
rect 15992 22272 16008 22336
rect 16072 22272 16088 22336
rect 16152 22272 16160 22336
rect 15840 21248 16160 22272
rect 15840 21184 15848 21248
rect 15912 21184 15928 21248
rect 15992 21184 16008 21248
rect 16072 21184 16088 21248
rect 16152 21184 16160 21248
rect 15840 20160 16160 21184
rect 15840 20096 15848 20160
rect 15912 20096 15928 20160
rect 15992 20096 16008 20160
rect 16072 20096 16088 20160
rect 16152 20096 16160 20160
rect 15840 19072 16160 20096
rect 15840 19008 15848 19072
rect 15912 19008 15928 19072
rect 15992 19008 16008 19072
rect 16072 19008 16088 19072
rect 16152 19008 16160 19072
rect 15840 17984 16160 19008
rect 15840 17920 15848 17984
rect 15912 17920 15928 17984
rect 15992 17920 16008 17984
rect 16072 17920 16088 17984
rect 16152 17920 16160 17984
rect 15840 16896 16160 17920
rect 15840 16832 15848 16896
rect 15912 16832 15928 16896
rect 15992 16832 16008 16896
rect 16072 16832 16088 16896
rect 16152 16832 16160 16896
rect 15840 15808 16160 16832
rect 17726 16149 17786 50763
rect 19198 28117 19258 53755
rect 20805 53344 21125 54368
rect 20805 53280 20813 53344
rect 20877 53280 20893 53344
rect 20957 53280 20973 53344
rect 21037 53280 21053 53344
rect 21117 53280 21125 53344
rect 20805 52256 21125 53280
rect 23243 52868 23309 52869
rect 23243 52804 23244 52868
rect 23308 52804 23309 52868
rect 23243 52803 23309 52804
rect 20805 52192 20813 52256
rect 20877 52192 20893 52256
rect 20957 52192 20973 52256
rect 21037 52192 21053 52256
rect 21117 52192 21125 52256
rect 20805 51168 21125 52192
rect 20805 51104 20813 51168
rect 20877 51104 20893 51168
rect 20957 51104 20973 51168
rect 21037 51104 21053 51168
rect 21117 51104 21125 51168
rect 20805 50080 21125 51104
rect 21403 50964 21469 50965
rect 21403 50900 21404 50964
rect 21468 50900 21469 50964
rect 21403 50899 21469 50900
rect 20805 50016 20813 50080
rect 20877 50016 20893 50080
rect 20957 50016 20973 50080
rect 21037 50016 21053 50080
rect 21117 50016 21125 50080
rect 20805 48992 21125 50016
rect 20805 48928 20813 48992
rect 20877 48928 20893 48992
rect 20957 48928 20973 48992
rect 21037 48928 21053 48992
rect 21117 48928 21125 48992
rect 20805 47904 21125 48928
rect 20805 47840 20813 47904
rect 20877 47840 20893 47904
rect 20957 47840 20973 47904
rect 21037 47840 21053 47904
rect 21117 47840 21125 47904
rect 20805 46816 21125 47840
rect 20805 46752 20813 46816
rect 20877 46752 20893 46816
rect 20957 46752 20973 46816
rect 21037 46752 21053 46816
rect 21117 46752 21125 46816
rect 20805 45728 21125 46752
rect 20805 45664 20813 45728
rect 20877 45664 20893 45728
rect 20957 45664 20973 45728
rect 21037 45664 21053 45728
rect 21117 45664 21125 45728
rect 20805 44640 21125 45664
rect 20805 44576 20813 44640
rect 20877 44576 20893 44640
rect 20957 44576 20973 44640
rect 21037 44576 21053 44640
rect 21117 44576 21125 44640
rect 20805 43552 21125 44576
rect 20805 43488 20813 43552
rect 20877 43488 20893 43552
rect 20957 43488 20973 43552
rect 21037 43488 21053 43552
rect 21117 43488 21125 43552
rect 20805 42464 21125 43488
rect 21406 43349 21466 50899
rect 23246 49877 23306 52803
rect 23430 51373 23490 56883
rect 23611 56676 23677 56677
rect 23611 56612 23612 56676
rect 23676 56612 23677 56676
rect 23611 56611 23677 56612
rect 23614 53821 23674 56611
rect 23795 55860 23861 55861
rect 23795 55796 23796 55860
rect 23860 55796 23861 55860
rect 23795 55795 23861 55796
rect 23611 53820 23677 53821
rect 23611 53756 23612 53820
rect 23676 53756 23677 53820
rect 23611 53755 23677 53756
rect 23614 52461 23674 53755
rect 23611 52460 23677 52461
rect 23611 52396 23612 52460
rect 23676 52396 23677 52460
rect 23611 52395 23677 52396
rect 23427 51372 23493 51373
rect 23427 51308 23428 51372
rect 23492 51308 23493 51372
rect 23427 51307 23493 51308
rect 23611 51372 23677 51373
rect 23611 51308 23612 51372
rect 23676 51308 23677 51372
rect 23611 51307 23677 51308
rect 23614 50421 23674 51307
rect 23611 50420 23677 50421
rect 23611 50356 23612 50420
rect 23676 50356 23677 50420
rect 23611 50355 23677 50356
rect 23798 50013 23858 55795
rect 23982 51509 24042 57291
rect 25086 56677 25146 65995
rect 25770 65856 26091 66880
rect 26371 66876 26437 66877
rect 26371 66812 26372 66876
rect 26436 66812 26437 66876
rect 26371 66811 26437 66812
rect 25770 65792 25778 65856
rect 25842 65792 25858 65856
rect 25922 65792 25938 65856
rect 26002 65792 26018 65856
rect 26082 65792 26091 65856
rect 25770 64768 26091 65792
rect 25770 64704 25778 64768
rect 25842 64704 25858 64768
rect 25922 64704 25938 64768
rect 26002 64704 26018 64768
rect 26082 64704 26091 64768
rect 25770 63680 26091 64704
rect 25770 63616 25778 63680
rect 25842 63616 25858 63680
rect 25922 63616 25938 63680
rect 26002 63616 26018 63680
rect 26082 63616 26091 63680
rect 25770 62592 26091 63616
rect 25770 62528 25778 62592
rect 25842 62528 25858 62592
rect 25922 62528 25938 62592
rect 26002 62528 26018 62592
rect 26082 62528 26091 62592
rect 25267 62388 25333 62389
rect 25267 62324 25268 62388
rect 25332 62324 25333 62388
rect 25267 62323 25333 62324
rect 25270 60893 25330 62323
rect 25770 61504 26091 62528
rect 26187 62388 26253 62389
rect 26187 62324 26188 62388
rect 26252 62324 26253 62388
rect 26187 62323 26253 62324
rect 25770 61440 25778 61504
rect 25842 61440 25858 61504
rect 25922 61440 25938 61504
rect 26002 61440 26018 61504
rect 26082 61440 26091 61504
rect 25267 60892 25333 60893
rect 25267 60828 25268 60892
rect 25332 60828 25333 60892
rect 25267 60827 25333 60828
rect 25770 60416 26091 61440
rect 25770 60352 25778 60416
rect 25842 60352 25858 60416
rect 25922 60352 25938 60416
rect 26002 60352 26018 60416
rect 26082 60352 26091 60416
rect 25267 59940 25333 59941
rect 25267 59876 25268 59940
rect 25332 59876 25333 59940
rect 25267 59875 25333 59876
rect 25270 57990 25330 59875
rect 25635 59668 25701 59669
rect 25635 59604 25636 59668
rect 25700 59604 25701 59668
rect 25635 59603 25701 59604
rect 25270 57930 25514 57990
rect 25083 56676 25149 56677
rect 25083 56612 25084 56676
rect 25148 56612 25149 56676
rect 25083 56611 25149 56612
rect 24899 55860 24965 55861
rect 24899 55796 24900 55860
rect 24964 55796 24965 55860
rect 24899 55795 24965 55796
rect 24531 54908 24597 54909
rect 24531 54844 24532 54908
rect 24596 54844 24597 54908
rect 24531 54843 24597 54844
rect 24715 54908 24781 54909
rect 24715 54844 24716 54908
rect 24780 54844 24781 54908
rect 24715 54843 24781 54844
rect 24163 53004 24229 53005
rect 24163 52940 24164 53004
rect 24228 52940 24229 53004
rect 24163 52939 24229 52940
rect 23979 51508 24045 51509
rect 23979 51444 23980 51508
rect 24044 51444 24045 51508
rect 23979 51443 24045 51444
rect 24166 51370 24226 52939
rect 24347 51644 24413 51645
rect 24347 51580 24348 51644
rect 24412 51580 24413 51644
rect 24347 51579 24413 51580
rect 23982 51310 24226 51370
rect 23982 50013 24042 51310
rect 24163 50964 24229 50965
rect 24163 50900 24164 50964
rect 24228 50900 24229 50964
rect 24163 50899 24229 50900
rect 23795 50012 23861 50013
rect 23795 49948 23796 50012
rect 23860 49948 23861 50012
rect 23795 49947 23861 49948
rect 23979 50012 24045 50013
rect 23979 49948 23980 50012
rect 24044 49948 24045 50012
rect 23979 49947 24045 49948
rect 23243 49876 23309 49877
rect 23243 49812 23244 49876
rect 23308 49812 23309 49876
rect 23243 49811 23309 49812
rect 24166 48789 24226 50899
rect 24350 49741 24410 51579
rect 24534 51101 24594 54843
rect 24531 51100 24597 51101
rect 24531 51036 24532 51100
rect 24596 51036 24597 51100
rect 24531 51035 24597 51036
rect 24531 50964 24597 50965
rect 24531 50900 24532 50964
rect 24596 50900 24597 50964
rect 24531 50899 24597 50900
rect 24534 50557 24594 50899
rect 24718 50693 24778 54843
rect 24715 50692 24781 50693
rect 24715 50628 24716 50692
rect 24780 50628 24781 50692
rect 24715 50627 24781 50628
rect 24531 50556 24597 50557
rect 24531 50492 24532 50556
rect 24596 50492 24597 50556
rect 24531 50491 24597 50492
rect 24715 50012 24781 50013
rect 24715 49948 24716 50012
rect 24780 49948 24781 50012
rect 24715 49947 24781 49948
rect 24347 49740 24413 49741
rect 24347 49676 24348 49740
rect 24412 49676 24413 49740
rect 24347 49675 24413 49676
rect 24531 48924 24597 48925
rect 24531 48860 24532 48924
rect 24596 48860 24597 48924
rect 24531 48859 24597 48860
rect 24163 48788 24229 48789
rect 24163 48724 24164 48788
rect 24228 48724 24229 48788
rect 24163 48723 24229 48724
rect 23243 46476 23309 46477
rect 23243 46412 23244 46476
rect 23308 46412 23309 46476
rect 23243 46411 23309 46412
rect 21403 43348 21469 43349
rect 21403 43284 21404 43348
rect 21468 43284 21469 43348
rect 21403 43283 21469 43284
rect 20805 42400 20813 42464
rect 20877 42400 20893 42464
rect 20957 42400 20973 42464
rect 21037 42400 21053 42464
rect 21117 42400 21125 42464
rect 20805 41376 21125 42400
rect 23246 42397 23306 46411
rect 24347 45116 24413 45117
rect 24347 45052 24348 45116
rect 24412 45052 24413 45116
rect 24347 45051 24413 45052
rect 23979 43212 24045 43213
rect 23979 43148 23980 43212
rect 24044 43148 24045 43212
rect 23979 43147 24045 43148
rect 23243 42396 23309 42397
rect 23243 42332 23244 42396
rect 23308 42332 23309 42396
rect 23243 42331 23309 42332
rect 20805 41312 20813 41376
rect 20877 41312 20893 41376
rect 20957 41312 20973 41376
rect 21037 41312 21053 41376
rect 21117 41312 21125 41376
rect 20805 40288 21125 41312
rect 20805 40224 20813 40288
rect 20877 40224 20893 40288
rect 20957 40224 20973 40288
rect 21037 40224 21053 40288
rect 21117 40224 21125 40288
rect 20805 39200 21125 40224
rect 20805 39136 20813 39200
rect 20877 39136 20893 39200
rect 20957 39136 20973 39200
rect 21037 39136 21053 39200
rect 21117 39136 21125 39200
rect 20805 38112 21125 39136
rect 23611 38996 23677 38997
rect 23611 38932 23612 38996
rect 23676 38932 23677 38996
rect 23611 38931 23677 38932
rect 20805 38048 20813 38112
rect 20877 38048 20893 38112
rect 20957 38048 20973 38112
rect 21037 38048 21053 38112
rect 21117 38048 21125 38112
rect 20805 37024 21125 38048
rect 23614 38045 23674 38931
rect 23611 38044 23677 38045
rect 23611 37980 23612 38044
rect 23676 37980 23677 38044
rect 23611 37979 23677 37980
rect 23982 37773 24042 43147
rect 24163 41580 24229 41581
rect 24163 41516 24164 41580
rect 24228 41516 24229 41580
rect 24163 41515 24229 41516
rect 24166 39949 24226 41515
rect 24350 41445 24410 45051
rect 24347 41444 24413 41445
rect 24347 41380 24348 41444
rect 24412 41380 24413 41444
rect 24347 41379 24413 41380
rect 24347 41172 24413 41173
rect 24347 41108 24348 41172
rect 24412 41108 24413 41172
rect 24347 41107 24413 41108
rect 24163 39948 24229 39949
rect 24163 39884 24164 39948
rect 24228 39884 24229 39948
rect 24163 39883 24229 39884
rect 23979 37772 24045 37773
rect 23979 37708 23980 37772
rect 24044 37708 24045 37772
rect 23979 37707 24045 37708
rect 20805 36960 20813 37024
rect 20877 36960 20893 37024
rect 20957 36960 20973 37024
rect 21037 36960 21053 37024
rect 21117 36960 21125 37024
rect 20805 35936 21125 36960
rect 20805 35872 20813 35936
rect 20877 35872 20893 35936
rect 20957 35872 20973 35936
rect 21037 35872 21053 35936
rect 21117 35872 21125 35936
rect 20805 34848 21125 35872
rect 24166 35325 24226 39883
rect 24163 35324 24229 35325
rect 24163 35260 24164 35324
rect 24228 35260 24229 35324
rect 24163 35259 24229 35260
rect 20805 34784 20813 34848
rect 20877 34784 20893 34848
rect 20957 34784 20973 34848
rect 21037 34784 21053 34848
rect 21117 34784 21125 34848
rect 20805 33760 21125 34784
rect 20805 33696 20813 33760
rect 20877 33696 20893 33760
rect 20957 33696 20973 33760
rect 21037 33696 21053 33760
rect 21117 33696 21125 33760
rect 20805 32672 21125 33696
rect 20805 32608 20813 32672
rect 20877 32608 20893 32672
rect 20957 32608 20973 32672
rect 21037 32608 21053 32672
rect 21117 32608 21125 32672
rect 20805 31584 21125 32608
rect 23243 32196 23309 32197
rect 23243 32132 23244 32196
rect 23308 32132 23309 32196
rect 23243 32131 23309 32132
rect 20805 31520 20813 31584
rect 20877 31520 20893 31584
rect 20957 31520 20973 31584
rect 21037 31520 21053 31584
rect 21117 31520 21125 31584
rect 20805 30496 21125 31520
rect 23246 31517 23306 32131
rect 23243 31516 23309 31517
rect 23243 31452 23244 31516
rect 23308 31452 23309 31516
rect 23243 31451 23309 31452
rect 20805 30432 20813 30496
rect 20877 30432 20893 30496
rect 20957 30432 20973 30496
rect 21037 30432 21053 30496
rect 21117 30432 21125 30496
rect 20805 29408 21125 30432
rect 24166 30293 24226 35259
rect 24350 33829 24410 41107
rect 24534 38317 24594 48859
rect 24718 43213 24778 49947
rect 24902 48517 24962 55795
rect 25083 55044 25149 55045
rect 25083 54980 25084 55044
rect 25148 54980 25149 55044
rect 25083 54979 25149 54980
rect 24899 48516 24965 48517
rect 24899 48452 24900 48516
rect 24964 48452 24965 48516
rect 24899 48451 24965 48452
rect 25086 46610 25146 54979
rect 25267 54092 25333 54093
rect 25267 54028 25268 54092
rect 25332 54028 25333 54092
rect 25267 54027 25333 54028
rect 25270 48109 25330 54027
rect 25454 51098 25514 57930
rect 25638 51237 25698 59603
rect 25770 59328 26091 60352
rect 26190 60213 26250 62323
rect 26374 60893 26434 66811
rect 26555 63748 26621 63749
rect 26555 63684 26556 63748
rect 26620 63684 26621 63748
rect 26555 63683 26621 63684
rect 26558 61029 26618 63683
rect 26923 61436 26989 61437
rect 26923 61372 26924 61436
rect 26988 61372 26989 61436
rect 26923 61371 26989 61372
rect 26739 61300 26805 61301
rect 26739 61236 26740 61300
rect 26804 61236 26805 61300
rect 26739 61235 26805 61236
rect 26555 61028 26621 61029
rect 26555 60964 26556 61028
rect 26620 60964 26621 61028
rect 26555 60963 26621 60964
rect 26371 60892 26437 60893
rect 26371 60828 26372 60892
rect 26436 60828 26437 60892
rect 26371 60827 26437 60828
rect 26742 60750 26802 61235
rect 26558 60690 26802 60750
rect 26187 60212 26253 60213
rect 26187 60148 26188 60212
rect 26252 60148 26253 60212
rect 26187 60147 26253 60148
rect 26558 59533 26618 60690
rect 26739 60484 26805 60485
rect 26739 60420 26740 60484
rect 26804 60420 26805 60484
rect 26739 60419 26805 60420
rect 26555 59532 26621 59533
rect 26555 59468 26556 59532
rect 26620 59468 26621 59532
rect 26555 59467 26621 59468
rect 25770 59264 25778 59328
rect 25842 59264 25858 59328
rect 25922 59264 25938 59328
rect 26002 59264 26018 59328
rect 26082 59264 26091 59328
rect 25770 58240 26091 59264
rect 25770 58176 25778 58240
rect 25842 58176 25858 58240
rect 25922 58176 25938 58240
rect 26002 58176 26018 58240
rect 26082 58176 26091 58240
rect 25770 57152 26091 58176
rect 26187 57628 26253 57629
rect 26187 57564 26188 57628
rect 26252 57564 26253 57628
rect 26187 57563 26253 57564
rect 25770 57088 25778 57152
rect 25842 57088 25858 57152
rect 25922 57088 25938 57152
rect 26002 57088 26018 57152
rect 26082 57088 26091 57152
rect 25770 56064 26091 57088
rect 25770 56000 25778 56064
rect 25842 56000 25858 56064
rect 25922 56000 25938 56064
rect 26002 56000 26018 56064
rect 26082 56000 26091 56064
rect 25770 54976 26091 56000
rect 25770 54912 25778 54976
rect 25842 54912 25858 54976
rect 25922 54912 25938 54976
rect 26002 54912 26018 54976
rect 26082 54912 26091 54976
rect 25770 53888 26091 54912
rect 25770 53824 25778 53888
rect 25842 53824 25858 53888
rect 25922 53824 25938 53888
rect 26002 53824 26018 53888
rect 26082 53824 26091 53888
rect 25770 52800 26091 53824
rect 25770 52736 25778 52800
rect 25842 52736 25858 52800
rect 25922 52736 25938 52800
rect 26002 52736 26018 52800
rect 26082 52736 26091 52800
rect 25770 51712 26091 52736
rect 25770 51648 25778 51712
rect 25842 51648 25858 51712
rect 25922 51648 25938 51712
rect 26002 51648 26018 51712
rect 26082 51648 26091 51712
rect 25635 51236 25701 51237
rect 25635 51172 25636 51236
rect 25700 51172 25701 51236
rect 25635 51171 25701 51172
rect 25454 51038 25698 51098
rect 25451 50420 25517 50421
rect 25451 50356 25452 50420
rect 25516 50356 25517 50420
rect 25451 50355 25517 50356
rect 25267 48108 25333 48109
rect 25267 48044 25268 48108
rect 25332 48044 25333 48108
rect 25267 48043 25333 48044
rect 25270 46749 25330 48043
rect 25267 46748 25333 46749
rect 25267 46684 25268 46748
rect 25332 46684 25333 46748
rect 25267 46683 25333 46684
rect 25086 46550 25330 46610
rect 24899 46476 24965 46477
rect 24899 46412 24900 46476
rect 24964 46412 24965 46476
rect 24899 46411 24965 46412
rect 24715 43212 24781 43213
rect 24715 43148 24716 43212
rect 24780 43148 24781 43212
rect 24715 43147 24781 43148
rect 24715 42260 24781 42261
rect 24715 42196 24716 42260
rect 24780 42196 24781 42260
rect 24715 42195 24781 42196
rect 24531 38316 24597 38317
rect 24531 38252 24532 38316
rect 24596 38252 24597 38316
rect 24531 38251 24597 38252
rect 24718 37501 24778 42195
rect 24902 41309 24962 46411
rect 25083 46204 25149 46205
rect 25083 46140 25084 46204
rect 25148 46140 25149 46204
rect 25083 46139 25149 46140
rect 24899 41308 24965 41309
rect 24899 41244 24900 41308
rect 24964 41244 24965 41308
rect 24899 41243 24965 41244
rect 24899 38452 24965 38453
rect 24899 38388 24900 38452
rect 24964 38388 24965 38452
rect 24899 38387 24965 38388
rect 24902 37637 24962 38387
rect 25086 38181 25146 46139
rect 25270 42941 25330 46550
rect 25267 42940 25333 42941
rect 25267 42876 25268 42940
rect 25332 42876 25333 42940
rect 25267 42875 25333 42876
rect 25267 42668 25333 42669
rect 25267 42604 25268 42668
rect 25332 42604 25333 42668
rect 25267 42603 25333 42604
rect 25270 41581 25330 42603
rect 25267 41580 25333 41581
rect 25267 41516 25268 41580
rect 25332 41516 25333 41580
rect 25267 41515 25333 41516
rect 25454 41173 25514 50355
rect 25451 41172 25517 41173
rect 25451 41108 25452 41172
rect 25516 41108 25517 41172
rect 25451 41107 25517 41108
rect 25451 40900 25517 40901
rect 25451 40836 25452 40900
rect 25516 40836 25517 40900
rect 25451 40835 25517 40836
rect 25267 38588 25333 38589
rect 25267 38524 25268 38588
rect 25332 38524 25333 38588
rect 25267 38523 25333 38524
rect 25083 38180 25149 38181
rect 25083 38116 25084 38180
rect 25148 38116 25149 38180
rect 25083 38115 25149 38116
rect 24899 37636 24965 37637
rect 24899 37572 24900 37636
rect 24964 37572 24965 37636
rect 24899 37571 24965 37572
rect 24715 37500 24781 37501
rect 24715 37436 24716 37500
rect 24780 37436 24781 37500
rect 24715 37435 24781 37436
rect 25270 37229 25330 38523
rect 25454 38181 25514 40835
rect 25638 40357 25698 51038
rect 25770 50624 26091 51648
rect 25770 50560 25778 50624
rect 25842 50560 25858 50624
rect 25922 50560 25938 50624
rect 26002 50560 26018 50624
rect 26082 50560 26091 50624
rect 25770 49536 26091 50560
rect 25770 49472 25778 49536
rect 25842 49472 25858 49536
rect 25922 49472 25938 49536
rect 26002 49472 26018 49536
rect 26082 49472 26091 49536
rect 25770 48448 26091 49472
rect 25770 48384 25778 48448
rect 25842 48384 25858 48448
rect 25922 48384 25938 48448
rect 26002 48384 26018 48448
rect 26082 48384 26091 48448
rect 25770 47360 26091 48384
rect 26190 47837 26250 57563
rect 26371 57356 26437 57357
rect 26371 57292 26372 57356
rect 26436 57292 26437 57356
rect 26371 57291 26437 57292
rect 26374 54365 26434 57291
rect 26371 54364 26437 54365
rect 26371 54300 26372 54364
rect 26436 54300 26437 54364
rect 26371 54299 26437 54300
rect 26371 54228 26437 54229
rect 26371 54164 26372 54228
rect 26436 54164 26437 54228
rect 26371 54163 26437 54164
rect 26374 51373 26434 54163
rect 26558 52325 26618 59467
rect 26555 52324 26621 52325
rect 26555 52260 26556 52324
rect 26620 52260 26621 52324
rect 26555 52259 26621 52260
rect 26555 52188 26621 52189
rect 26555 52124 26556 52188
rect 26620 52124 26621 52188
rect 26555 52123 26621 52124
rect 26371 51372 26437 51373
rect 26371 51308 26372 51372
rect 26436 51308 26437 51372
rect 26371 51307 26437 51308
rect 26371 51236 26437 51237
rect 26371 51172 26372 51236
rect 26436 51172 26437 51236
rect 26371 51171 26437 51172
rect 26187 47836 26253 47837
rect 26187 47772 26188 47836
rect 26252 47772 26253 47836
rect 26187 47771 26253 47772
rect 25770 47296 25778 47360
rect 25842 47296 25858 47360
rect 25922 47296 25938 47360
rect 26002 47296 26018 47360
rect 26082 47296 26091 47360
rect 25770 46272 26091 47296
rect 26374 46885 26434 51171
rect 26371 46884 26437 46885
rect 26371 46820 26372 46884
rect 26436 46820 26437 46884
rect 26371 46819 26437 46820
rect 26187 46476 26253 46477
rect 26187 46412 26188 46476
rect 26252 46412 26253 46476
rect 26187 46411 26253 46412
rect 25770 46208 25778 46272
rect 25842 46208 25858 46272
rect 25922 46208 25938 46272
rect 26002 46208 26018 46272
rect 26082 46208 26091 46272
rect 25770 45184 26091 46208
rect 25770 45120 25778 45184
rect 25842 45120 25858 45184
rect 25922 45120 25938 45184
rect 26002 45120 26018 45184
rect 26082 45120 26091 45184
rect 25770 44096 26091 45120
rect 25770 44032 25778 44096
rect 25842 44032 25858 44096
rect 25922 44032 25938 44096
rect 26002 44032 26018 44096
rect 26082 44032 26091 44096
rect 25770 43008 26091 44032
rect 25770 42944 25778 43008
rect 25842 42944 25858 43008
rect 25922 42944 25938 43008
rect 26002 42944 26018 43008
rect 26082 42944 26091 43008
rect 25770 41920 26091 42944
rect 26190 42805 26250 46411
rect 26371 45116 26437 45117
rect 26371 45052 26372 45116
rect 26436 45052 26437 45116
rect 26371 45051 26437 45052
rect 26187 42804 26253 42805
rect 26187 42740 26188 42804
rect 26252 42740 26253 42804
rect 26187 42739 26253 42740
rect 26187 42396 26253 42397
rect 26187 42332 26188 42396
rect 26252 42332 26253 42396
rect 26187 42331 26253 42332
rect 25770 41856 25778 41920
rect 25842 41856 25858 41920
rect 25922 41856 25938 41920
rect 26002 41856 26018 41920
rect 26082 41856 26091 41920
rect 25770 40832 26091 41856
rect 25770 40768 25778 40832
rect 25842 40768 25858 40832
rect 25922 40768 25938 40832
rect 26002 40768 26018 40832
rect 26082 40768 26091 40832
rect 25635 40356 25701 40357
rect 25635 40292 25636 40356
rect 25700 40292 25701 40356
rect 25635 40291 25701 40292
rect 25770 39744 26091 40768
rect 25770 39680 25778 39744
rect 25842 39680 25858 39744
rect 25922 39680 25938 39744
rect 26002 39680 26018 39744
rect 26082 39680 26091 39744
rect 25635 38860 25701 38861
rect 25635 38796 25636 38860
rect 25700 38796 25701 38860
rect 25635 38795 25701 38796
rect 25451 38180 25517 38181
rect 25451 38116 25452 38180
rect 25516 38116 25517 38180
rect 25451 38115 25517 38116
rect 25451 37908 25517 37909
rect 25451 37844 25452 37908
rect 25516 37844 25517 37908
rect 25451 37843 25517 37844
rect 25267 37228 25333 37229
rect 25267 37164 25268 37228
rect 25332 37164 25333 37228
rect 25267 37163 25333 37164
rect 24899 36684 24965 36685
rect 24899 36620 24900 36684
rect 24964 36620 24965 36684
rect 24899 36619 24965 36620
rect 24347 33828 24413 33829
rect 24347 33764 24348 33828
rect 24412 33764 24413 33828
rect 24347 33763 24413 33764
rect 24715 32060 24781 32061
rect 24715 31996 24716 32060
rect 24780 31996 24781 32060
rect 24715 31995 24781 31996
rect 24163 30292 24229 30293
rect 24163 30228 24164 30292
rect 24228 30228 24229 30292
rect 24163 30227 24229 30228
rect 22139 29884 22205 29885
rect 22139 29820 22140 29884
rect 22204 29820 22205 29884
rect 22139 29819 22205 29820
rect 20805 29344 20813 29408
rect 20877 29344 20893 29408
rect 20957 29344 20973 29408
rect 21037 29344 21053 29408
rect 21117 29344 21125 29408
rect 20805 28320 21125 29344
rect 20805 28256 20813 28320
rect 20877 28256 20893 28320
rect 20957 28256 20973 28320
rect 21037 28256 21053 28320
rect 21117 28256 21125 28320
rect 19195 28116 19261 28117
rect 19195 28052 19196 28116
rect 19260 28052 19261 28116
rect 19195 28051 19261 28052
rect 20805 27232 21125 28256
rect 20805 27168 20813 27232
rect 20877 27168 20893 27232
rect 20957 27168 20973 27232
rect 21037 27168 21053 27232
rect 21117 27168 21125 27232
rect 20805 26144 21125 27168
rect 20805 26080 20813 26144
rect 20877 26080 20893 26144
rect 20957 26080 20973 26144
rect 21037 26080 21053 26144
rect 21117 26080 21125 26144
rect 20805 25056 21125 26080
rect 20805 24992 20813 25056
rect 20877 24992 20893 25056
rect 20957 24992 20973 25056
rect 21037 24992 21053 25056
rect 21117 24992 21125 25056
rect 20805 23968 21125 24992
rect 22142 24853 22202 29819
rect 22139 24852 22205 24853
rect 22139 24788 22140 24852
rect 22204 24788 22205 24852
rect 22139 24787 22205 24788
rect 20805 23904 20813 23968
rect 20877 23904 20893 23968
rect 20957 23904 20973 23968
rect 21037 23904 21053 23968
rect 21117 23904 21125 23968
rect 20805 22880 21125 23904
rect 20805 22816 20813 22880
rect 20877 22816 20893 22880
rect 20957 22816 20973 22880
rect 21037 22816 21053 22880
rect 21117 22816 21125 22880
rect 20805 21792 21125 22816
rect 24718 22813 24778 31995
rect 24902 29749 24962 36619
rect 25454 36141 25514 37843
rect 25451 36140 25517 36141
rect 25451 36076 25452 36140
rect 25516 36076 25517 36140
rect 25451 36075 25517 36076
rect 25451 36004 25517 36005
rect 25451 35940 25452 36004
rect 25516 35940 25517 36004
rect 25451 35939 25517 35940
rect 25083 35868 25149 35869
rect 25083 35804 25084 35868
rect 25148 35804 25149 35868
rect 25083 35803 25149 35804
rect 25086 31381 25146 35803
rect 25267 35732 25333 35733
rect 25267 35668 25268 35732
rect 25332 35668 25333 35732
rect 25267 35667 25333 35668
rect 25270 31789 25330 35667
rect 25267 31788 25333 31789
rect 25267 31724 25268 31788
rect 25332 31724 25333 31788
rect 25267 31723 25333 31724
rect 25454 31650 25514 35939
rect 25638 33013 25698 38795
rect 25770 38656 26091 39680
rect 26190 39541 26250 42331
rect 26374 41581 26434 45051
rect 26371 41580 26437 41581
rect 26371 41516 26372 41580
rect 26436 41516 26437 41580
rect 26371 41515 26437 41516
rect 26371 41444 26437 41445
rect 26371 41380 26372 41444
rect 26436 41380 26437 41444
rect 26371 41379 26437 41380
rect 26187 39540 26253 39541
rect 26187 39476 26188 39540
rect 26252 39476 26253 39540
rect 26187 39475 26253 39476
rect 26374 39405 26434 41379
rect 26371 39404 26437 39405
rect 26371 39340 26372 39404
rect 26436 39340 26437 39404
rect 26371 39339 26437 39340
rect 26371 39268 26437 39269
rect 26371 39204 26372 39268
rect 26436 39204 26437 39268
rect 26371 39203 26437 39204
rect 26187 38996 26253 38997
rect 26187 38932 26188 38996
rect 26252 38932 26253 38996
rect 26187 38931 26253 38932
rect 25770 38592 25778 38656
rect 25842 38592 25858 38656
rect 25922 38592 25938 38656
rect 26002 38592 26018 38656
rect 26082 38592 26091 38656
rect 25770 37568 26091 38592
rect 26190 37909 26250 38931
rect 26374 38589 26434 39203
rect 26371 38588 26437 38589
rect 26371 38524 26372 38588
rect 26436 38524 26437 38588
rect 26371 38523 26437 38524
rect 26187 37908 26253 37909
rect 26187 37844 26188 37908
rect 26252 37844 26253 37908
rect 26187 37843 26253 37844
rect 25770 37504 25778 37568
rect 25842 37504 25858 37568
rect 25922 37504 25938 37568
rect 26002 37504 26018 37568
rect 26082 37504 26091 37568
rect 25770 36480 26091 37504
rect 26371 37364 26437 37365
rect 26371 37300 26372 37364
rect 26436 37300 26437 37364
rect 26371 37299 26437 37300
rect 25770 36416 25778 36480
rect 25842 36416 25858 36480
rect 25922 36416 25938 36480
rect 26002 36416 26018 36480
rect 26082 36416 26091 36480
rect 25770 35392 26091 36416
rect 25770 35328 25778 35392
rect 25842 35328 25858 35392
rect 25922 35328 25938 35392
rect 26002 35328 26018 35392
rect 26082 35328 26091 35392
rect 25770 34304 26091 35328
rect 25770 34240 25778 34304
rect 25842 34240 25858 34304
rect 25922 34240 25938 34304
rect 26002 34240 26018 34304
rect 26082 34240 26091 34304
rect 25770 33216 26091 34240
rect 25770 33152 25778 33216
rect 25842 33152 25858 33216
rect 25922 33152 25938 33216
rect 26002 33152 26018 33216
rect 26082 33152 26091 33216
rect 25635 33012 25701 33013
rect 25635 32948 25636 33012
rect 25700 32948 25701 33012
rect 25635 32947 25701 32948
rect 25635 32876 25701 32877
rect 25635 32812 25636 32876
rect 25700 32812 25701 32876
rect 25635 32811 25701 32812
rect 25270 31590 25514 31650
rect 25083 31380 25149 31381
rect 25083 31316 25084 31380
rect 25148 31316 25149 31380
rect 25083 31315 25149 31316
rect 25270 30701 25330 31590
rect 25451 31244 25517 31245
rect 25451 31180 25452 31244
rect 25516 31180 25517 31244
rect 25451 31179 25517 31180
rect 25267 30700 25333 30701
rect 25267 30636 25268 30700
rect 25332 30636 25333 30700
rect 25267 30635 25333 30636
rect 25267 30156 25333 30157
rect 25267 30092 25268 30156
rect 25332 30092 25333 30156
rect 25267 30091 25333 30092
rect 24899 29748 24965 29749
rect 24899 29684 24900 29748
rect 24964 29684 24965 29748
rect 24899 29683 24965 29684
rect 25083 28660 25149 28661
rect 25083 28596 25084 28660
rect 25148 28596 25149 28660
rect 25083 28595 25149 28596
rect 24899 25396 24965 25397
rect 24899 25332 24900 25396
rect 24964 25332 24965 25396
rect 24899 25331 24965 25332
rect 24902 23085 24962 25331
rect 24899 23084 24965 23085
rect 24899 23020 24900 23084
rect 24964 23020 24965 23084
rect 24899 23019 24965 23020
rect 24715 22812 24781 22813
rect 24715 22748 24716 22812
rect 24780 22748 24781 22812
rect 24715 22747 24781 22748
rect 20805 21728 20813 21792
rect 20877 21728 20893 21792
rect 20957 21728 20973 21792
rect 21037 21728 21053 21792
rect 21117 21728 21125 21792
rect 20805 20704 21125 21728
rect 24902 21725 24962 23019
rect 24899 21724 24965 21725
rect 24899 21660 24900 21724
rect 24964 21660 24965 21724
rect 24899 21659 24965 21660
rect 25086 21453 25146 28595
rect 25270 25261 25330 30091
rect 25454 27981 25514 31179
rect 25451 27980 25517 27981
rect 25451 27916 25452 27980
rect 25516 27916 25517 27980
rect 25451 27915 25517 27916
rect 25451 27164 25517 27165
rect 25451 27100 25452 27164
rect 25516 27100 25517 27164
rect 25451 27099 25517 27100
rect 25267 25260 25333 25261
rect 25267 25196 25268 25260
rect 25332 25196 25333 25260
rect 25267 25195 25333 25196
rect 25267 24172 25333 24173
rect 25267 24108 25268 24172
rect 25332 24108 25333 24172
rect 25267 24107 25333 24108
rect 25083 21452 25149 21453
rect 25083 21388 25084 21452
rect 25148 21388 25149 21452
rect 25083 21387 25149 21388
rect 20805 20640 20813 20704
rect 20877 20640 20893 20704
rect 20957 20640 20973 20704
rect 21037 20640 21053 20704
rect 21117 20640 21125 20704
rect 20805 19616 21125 20640
rect 25270 19685 25330 24107
rect 25454 22133 25514 27099
rect 25638 26893 25698 32811
rect 25770 32128 26091 33152
rect 26187 32604 26253 32605
rect 26187 32540 26188 32604
rect 26252 32540 26253 32604
rect 26187 32539 26253 32540
rect 25770 32064 25778 32128
rect 25842 32064 25858 32128
rect 25922 32064 25938 32128
rect 26002 32064 26018 32128
rect 26082 32064 26091 32128
rect 25770 31040 26091 32064
rect 25770 30976 25778 31040
rect 25842 30976 25858 31040
rect 25922 30976 25938 31040
rect 26002 30976 26018 31040
rect 26082 30976 26091 31040
rect 25770 29952 26091 30976
rect 26190 30157 26250 32539
rect 26374 31653 26434 37299
rect 26558 36685 26618 52123
rect 26742 41445 26802 60419
rect 26926 60349 26986 61371
rect 26923 60348 26989 60349
rect 26923 60284 26924 60348
rect 26988 60284 26989 60348
rect 26923 60283 26989 60284
rect 27110 59261 27170 67491
rect 27659 65652 27725 65653
rect 27659 65588 27660 65652
rect 27724 65588 27725 65652
rect 27659 65587 27725 65588
rect 28395 65652 28461 65653
rect 28395 65588 28396 65652
rect 28460 65588 28461 65652
rect 28395 65587 28461 65588
rect 27475 62932 27541 62933
rect 27475 62868 27476 62932
rect 27540 62868 27541 62932
rect 27475 62867 27541 62868
rect 27291 60620 27357 60621
rect 27291 60556 27292 60620
rect 27356 60556 27357 60620
rect 27291 60555 27357 60556
rect 27107 59260 27173 59261
rect 27107 59196 27108 59260
rect 27172 59196 27173 59260
rect 27107 59195 27173 59196
rect 27294 58850 27354 60555
rect 27110 58790 27354 58850
rect 26923 57628 26989 57629
rect 26923 57564 26924 57628
rect 26988 57564 26989 57628
rect 26923 57563 26989 57564
rect 26926 51917 26986 57563
rect 27110 54773 27170 58790
rect 27478 57901 27538 62867
rect 27662 59805 27722 65587
rect 27843 64156 27909 64157
rect 27843 64092 27844 64156
rect 27908 64092 27909 64156
rect 27843 64091 27909 64092
rect 27846 60213 27906 64091
rect 28211 64020 28277 64021
rect 28211 63956 28212 64020
rect 28276 63956 28277 64020
rect 28211 63955 28277 63956
rect 28214 61165 28274 63955
rect 28398 63069 28458 65587
rect 28763 64972 28829 64973
rect 28763 64908 28764 64972
rect 28828 64908 28829 64972
rect 28763 64907 28829 64908
rect 28395 63068 28461 63069
rect 28395 63004 28396 63068
rect 28460 63004 28461 63068
rect 28395 63003 28461 63004
rect 28579 63068 28645 63069
rect 28579 63004 28580 63068
rect 28644 63004 28645 63068
rect 28579 63003 28645 63004
rect 28395 62116 28461 62117
rect 28395 62052 28396 62116
rect 28460 62052 28461 62116
rect 28395 62051 28461 62052
rect 28211 61164 28277 61165
rect 28211 61100 28212 61164
rect 28276 61100 28277 61164
rect 28211 61099 28277 61100
rect 28211 61028 28277 61029
rect 28211 60964 28212 61028
rect 28276 60964 28277 61028
rect 28211 60963 28277 60964
rect 28027 60348 28093 60349
rect 28027 60284 28028 60348
rect 28092 60284 28093 60348
rect 28027 60283 28093 60284
rect 27843 60212 27909 60213
rect 27843 60148 27844 60212
rect 27908 60148 27909 60212
rect 27843 60147 27909 60148
rect 27659 59804 27725 59805
rect 27659 59740 27660 59804
rect 27724 59740 27725 59804
rect 27659 59739 27725 59740
rect 27846 58581 27906 60147
rect 27843 58580 27909 58581
rect 27843 58516 27844 58580
rect 27908 58516 27909 58580
rect 27843 58515 27909 58516
rect 27475 57900 27541 57901
rect 27475 57836 27476 57900
rect 27540 57836 27541 57900
rect 27475 57835 27541 57836
rect 27475 57764 27541 57765
rect 27475 57700 27476 57764
rect 27540 57700 27541 57764
rect 27475 57699 27541 57700
rect 27291 55452 27357 55453
rect 27291 55388 27292 55452
rect 27356 55388 27357 55452
rect 27291 55387 27357 55388
rect 27107 54772 27173 54773
rect 27107 54708 27108 54772
rect 27172 54708 27173 54772
rect 27107 54707 27173 54708
rect 27107 53004 27173 53005
rect 27107 52940 27108 53004
rect 27172 52940 27173 53004
rect 27107 52939 27173 52940
rect 26923 51916 26989 51917
rect 26923 51852 26924 51916
rect 26988 51852 26989 51916
rect 26923 51851 26989 51852
rect 27110 51506 27170 52939
rect 27294 52189 27354 55387
rect 27291 52188 27357 52189
rect 27291 52124 27292 52188
rect 27356 52124 27357 52188
rect 27291 52123 27357 52124
rect 27291 52052 27357 52053
rect 27291 51988 27292 52052
rect 27356 51988 27357 52052
rect 27291 51987 27357 51988
rect 26926 51446 27170 51506
rect 26926 50013 26986 51446
rect 27107 51372 27173 51373
rect 27107 51308 27108 51372
rect 27172 51308 27173 51372
rect 27107 51307 27173 51308
rect 26923 50012 26989 50013
rect 26923 49948 26924 50012
rect 26988 49948 26989 50012
rect 26923 49947 26989 49948
rect 26923 49468 26989 49469
rect 26923 49404 26924 49468
rect 26988 49404 26989 49468
rect 26923 49403 26989 49404
rect 26926 48381 26986 49403
rect 26923 48380 26989 48381
rect 26923 48316 26924 48380
rect 26988 48316 26989 48380
rect 26923 48315 26989 48316
rect 26923 45524 26989 45525
rect 26923 45460 26924 45524
rect 26988 45460 26989 45524
rect 26923 45459 26989 45460
rect 26926 41714 26986 45459
rect 27110 42669 27170 51307
rect 27294 48109 27354 51987
rect 27478 49469 27538 57699
rect 27659 57220 27725 57221
rect 27659 57156 27660 57220
rect 27724 57156 27725 57220
rect 27659 57155 27725 57156
rect 27662 52053 27722 57155
rect 27843 53820 27909 53821
rect 27843 53756 27844 53820
rect 27908 53756 27909 53820
rect 27843 53755 27909 53756
rect 27659 52052 27725 52053
rect 27659 51988 27660 52052
rect 27724 51988 27725 52052
rect 27659 51987 27725 51988
rect 27659 51916 27725 51917
rect 27659 51852 27660 51916
rect 27724 51852 27725 51916
rect 27659 51851 27725 51852
rect 27662 51098 27722 51851
rect 27846 51237 27906 53755
rect 28030 53005 28090 60283
rect 28214 60077 28274 60963
rect 28211 60076 28277 60077
rect 28211 60012 28212 60076
rect 28276 60012 28277 60076
rect 28211 60011 28277 60012
rect 28398 59533 28458 62051
rect 28582 61709 28642 63003
rect 28579 61708 28645 61709
rect 28579 61644 28580 61708
rect 28644 61644 28645 61708
rect 28579 61643 28645 61644
rect 28766 61573 28826 64907
rect 28947 63476 29013 63477
rect 28947 63412 28948 63476
rect 29012 63412 29013 63476
rect 28947 63411 29013 63412
rect 28763 61572 28829 61573
rect 28763 61508 28764 61572
rect 28828 61508 28829 61572
rect 28763 61507 28829 61508
rect 28579 61300 28645 61301
rect 28579 61236 28580 61300
rect 28644 61236 28645 61300
rect 28579 61235 28645 61236
rect 28582 60213 28642 61235
rect 28579 60212 28645 60213
rect 28579 60148 28580 60212
rect 28644 60148 28645 60212
rect 28579 60147 28645 60148
rect 28395 59532 28461 59533
rect 28395 59468 28396 59532
rect 28460 59468 28461 59532
rect 28395 59467 28461 59468
rect 28766 58853 28826 61507
rect 28950 60077 29010 63411
rect 29134 61301 29194 69939
rect 29315 61436 29381 61437
rect 29315 61372 29316 61436
rect 29380 61372 29381 61436
rect 29315 61371 29381 61372
rect 29131 61300 29197 61301
rect 29131 61236 29132 61300
rect 29196 61236 29197 61300
rect 29131 61235 29197 61236
rect 29318 61162 29378 61371
rect 29134 61102 29378 61162
rect 29499 61164 29565 61165
rect 28947 60076 29013 60077
rect 28947 60012 28948 60076
rect 29012 60012 29013 60076
rect 28947 60011 29013 60012
rect 28763 58852 28829 58853
rect 28763 58788 28764 58852
rect 28828 58788 28829 58852
rect 28763 58787 28829 58788
rect 28763 58716 28829 58717
rect 28763 58652 28764 58716
rect 28828 58652 28829 58716
rect 28763 58651 28829 58652
rect 28211 55316 28277 55317
rect 28211 55252 28212 55316
rect 28276 55252 28277 55316
rect 28211 55251 28277 55252
rect 28027 53004 28093 53005
rect 28027 52940 28028 53004
rect 28092 52940 28093 53004
rect 28027 52939 28093 52940
rect 28027 52732 28093 52733
rect 28027 52668 28028 52732
rect 28092 52668 28093 52732
rect 28027 52667 28093 52668
rect 27843 51236 27909 51237
rect 27843 51172 27844 51236
rect 27908 51172 27909 51236
rect 27843 51171 27909 51172
rect 27662 51038 27906 51098
rect 27659 50964 27725 50965
rect 27659 50900 27660 50964
rect 27724 50900 27725 50964
rect 27659 50899 27725 50900
rect 27662 50149 27722 50899
rect 27659 50148 27725 50149
rect 27659 50084 27660 50148
rect 27724 50084 27725 50148
rect 27659 50083 27725 50084
rect 27475 49468 27541 49469
rect 27475 49404 27476 49468
rect 27540 49404 27541 49468
rect 27475 49403 27541 49404
rect 27478 48925 27538 49403
rect 27475 48924 27541 48925
rect 27475 48860 27476 48924
rect 27540 48860 27541 48924
rect 27475 48859 27541 48860
rect 27475 48788 27541 48789
rect 27475 48724 27476 48788
rect 27540 48724 27541 48788
rect 27475 48723 27541 48724
rect 27291 48108 27357 48109
rect 27291 48044 27292 48108
rect 27356 48044 27357 48108
rect 27291 48043 27357 48044
rect 27478 47973 27538 48723
rect 27475 47972 27541 47973
rect 27475 47908 27476 47972
rect 27540 47908 27541 47972
rect 27475 47907 27541 47908
rect 27475 44708 27541 44709
rect 27475 44644 27476 44708
rect 27540 44644 27541 44708
rect 27475 44643 27541 44644
rect 27291 44572 27357 44573
rect 27291 44508 27292 44572
rect 27356 44508 27357 44572
rect 27291 44507 27357 44508
rect 27107 42668 27173 42669
rect 27107 42604 27108 42668
rect 27172 42604 27173 42668
rect 27107 42603 27173 42604
rect 26926 41654 27170 41714
rect 26923 41580 26989 41581
rect 26923 41516 26924 41580
rect 26988 41516 26989 41580
rect 26923 41515 26989 41516
rect 26739 41444 26805 41445
rect 26739 41380 26740 41444
rect 26804 41380 26805 41444
rect 26739 41379 26805 41380
rect 26926 41173 26986 41515
rect 26923 41172 26989 41173
rect 26923 41108 26924 41172
rect 26988 41108 26989 41172
rect 26923 41107 26989 41108
rect 27110 39813 27170 41654
rect 27294 40901 27354 44507
rect 27291 40900 27357 40901
rect 27291 40836 27292 40900
rect 27356 40836 27357 40900
rect 27291 40835 27357 40836
rect 27478 40085 27538 44643
rect 27662 44437 27722 50083
rect 27846 48653 27906 51038
rect 27843 48652 27909 48653
rect 27843 48588 27844 48652
rect 27908 48588 27909 48652
rect 27843 48587 27909 48588
rect 28030 48517 28090 52667
rect 28027 48516 28093 48517
rect 28027 48452 28028 48516
rect 28092 48452 28093 48516
rect 28027 48451 28093 48452
rect 27843 46204 27909 46205
rect 27843 46140 27844 46204
rect 27908 46140 27909 46204
rect 27843 46139 27909 46140
rect 27659 44436 27725 44437
rect 27659 44372 27660 44436
rect 27724 44372 27725 44436
rect 27659 44371 27725 44372
rect 27659 43212 27725 43213
rect 27659 43148 27660 43212
rect 27724 43148 27725 43212
rect 27659 43147 27725 43148
rect 27662 41037 27722 43147
rect 27659 41036 27725 41037
rect 27659 40972 27660 41036
rect 27724 40972 27725 41036
rect 27659 40971 27725 40972
rect 27659 40900 27725 40901
rect 27659 40836 27660 40900
rect 27724 40836 27725 40900
rect 27659 40835 27725 40836
rect 27475 40084 27541 40085
rect 27475 40020 27476 40084
rect 27540 40020 27541 40084
rect 27475 40019 27541 40020
rect 27107 39812 27173 39813
rect 27107 39748 27108 39812
rect 27172 39748 27173 39812
rect 27107 39747 27173 39748
rect 26923 38180 26989 38181
rect 26923 38116 26924 38180
rect 26988 38116 26989 38180
rect 26923 38115 26989 38116
rect 26926 37501 26986 38115
rect 27475 37772 27541 37773
rect 27475 37708 27476 37772
rect 27540 37708 27541 37772
rect 27475 37707 27541 37708
rect 26923 37500 26989 37501
rect 26923 37436 26924 37500
rect 26988 37436 26989 37500
rect 26923 37435 26989 37436
rect 26739 37092 26805 37093
rect 26739 37028 26740 37092
rect 26804 37028 26805 37092
rect 26739 37027 26805 37028
rect 26555 36684 26621 36685
rect 26555 36620 26556 36684
rect 26620 36620 26621 36684
rect 26555 36619 26621 36620
rect 26555 32196 26621 32197
rect 26555 32132 26556 32196
rect 26620 32132 26621 32196
rect 26555 32131 26621 32132
rect 26371 31652 26437 31653
rect 26371 31588 26372 31652
rect 26436 31588 26437 31652
rect 26371 31587 26437 31588
rect 26371 30428 26437 30429
rect 26371 30364 26372 30428
rect 26436 30364 26437 30428
rect 26371 30363 26437 30364
rect 26187 30156 26253 30157
rect 26187 30092 26188 30156
rect 26252 30092 26253 30156
rect 26187 30091 26253 30092
rect 25770 29888 25778 29952
rect 25842 29888 25858 29952
rect 25922 29888 25938 29952
rect 26002 29888 26018 29952
rect 26082 29888 26091 29952
rect 25770 28864 26091 29888
rect 26187 29340 26253 29341
rect 26187 29276 26188 29340
rect 26252 29276 26253 29340
rect 26187 29275 26253 29276
rect 25770 28800 25778 28864
rect 25842 28800 25858 28864
rect 25922 28800 25938 28864
rect 26002 28800 26018 28864
rect 26082 28800 26091 28864
rect 25770 27776 26091 28800
rect 25770 27712 25778 27776
rect 25842 27712 25858 27776
rect 25922 27712 25938 27776
rect 26002 27712 26018 27776
rect 26082 27712 26091 27776
rect 25635 26892 25701 26893
rect 25635 26828 25636 26892
rect 25700 26828 25701 26892
rect 25635 26827 25701 26828
rect 25770 26688 26091 27712
rect 25770 26624 25778 26688
rect 25842 26624 25858 26688
rect 25922 26624 25938 26688
rect 26002 26624 26018 26688
rect 26082 26624 26091 26688
rect 25770 25600 26091 26624
rect 25770 25536 25778 25600
rect 25842 25536 25858 25600
rect 25922 25536 25938 25600
rect 26002 25536 26018 25600
rect 26082 25536 26091 25600
rect 25770 24512 26091 25536
rect 26190 24717 26250 29275
rect 26374 27981 26434 30363
rect 26371 27980 26437 27981
rect 26371 27916 26372 27980
rect 26436 27916 26437 27980
rect 26371 27915 26437 27916
rect 26371 27300 26437 27301
rect 26371 27236 26372 27300
rect 26436 27236 26437 27300
rect 26371 27235 26437 27236
rect 26187 24716 26253 24717
rect 26187 24652 26188 24716
rect 26252 24652 26253 24716
rect 26187 24651 26253 24652
rect 25770 24448 25778 24512
rect 25842 24448 25858 24512
rect 25922 24448 25938 24512
rect 26002 24448 26018 24512
rect 26082 24448 26091 24512
rect 25770 23424 26091 24448
rect 25770 23360 25778 23424
rect 25842 23360 25858 23424
rect 25922 23360 25938 23424
rect 26002 23360 26018 23424
rect 26082 23360 26091 23424
rect 25635 22404 25701 22405
rect 25635 22340 25636 22404
rect 25700 22340 25701 22404
rect 25635 22339 25701 22340
rect 25451 22132 25517 22133
rect 25451 22068 25452 22132
rect 25516 22068 25517 22132
rect 25451 22067 25517 22068
rect 25638 21045 25698 22339
rect 25770 22336 26091 23360
rect 26187 22812 26253 22813
rect 26187 22748 26188 22812
rect 26252 22748 26253 22812
rect 26187 22747 26253 22748
rect 25770 22272 25778 22336
rect 25842 22272 25858 22336
rect 25922 22272 25938 22336
rect 26002 22272 26018 22336
rect 26082 22272 26091 22336
rect 25770 21248 26091 22272
rect 25770 21184 25778 21248
rect 25842 21184 25858 21248
rect 25922 21184 25938 21248
rect 26002 21184 26018 21248
rect 26082 21184 26091 21248
rect 25635 21044 25701 21045
rect 25635 20980 25636 21044
rect 25700 20980 25701 21044
rect 25635 20979 25701 20980
rect 25770 20160 26091 21184
rect 25770 20096 25778 20160
rect 25842 20096 25858 20160
rect 25922 20096 25938 20160
rect 26002 20096 26018 20160
rect 26082 20096 26091 20160
rect 25267 19684 25333 19685
rect 25267 19620 25268 19684
rect 25332 19620 25333 19684
rect 25267 19619 25333 19620
rect 20805 19552 20813 19616
rect 20877 19552 20893 19616
rect 20957 19552 20973 19616
rect 21037 19552 21053 19616
rect 21117 19552 21125 19616
rect 20805 18528 21125 19552
rect 20805 18464 20813 18528
rect 20877 18464 20893 18528
rect 20957 18464 20973 18528
rect 21037 18464 21053 18528
rect 21117 18464 21125 18528
rect 20805 17440 21125 18464
rect 25770 19072 26091 20096
rect 25770 19008 25778 19072
rect 25842 19008 25858 19072
rect 25922 19008 25938 19072
rect 26002 19008 26018 19072
rect 26082 19008 26091 19072
rect 25635 18188 25701 18189
rect 25635 18124 25636 18188
rect 25700 18124 25701 18188
rect 25635 18123 25701 18124
rect 20805 17376 20813 17440
rect 20877 17376 20893 17440
rect 20957 17376 20973 17440
rect 21037 17376 21053 17440
rect 21117 17376 21125 17440
rect 20805 16352 21125 17376
rect 20805 16288 20813 16352
rect 20877 16288 20893 16352
rect 20957 16288 20973 16352
rect 21037 16288 21053 16352
rect 21117 16288 21125 16352
rect 17723 16148 17789 16149
rect 17723 16084 17724 16148
rect 17788 16084 17789 16148
rect 17723 16083 17789 16084
rect 15840 15744 15848 15808
rect 15912 15744 15928 15808
rect 15992 15744 16008 15808
rect 16072 15744 16088 15808
rect 16152 15744 16160 15808
rect 15840 14720 16160 15744
rect 15840 14656 15848 14720
rect 15912 14656 15928 14720
rect 15992 14656 16008 14720
rect 16072 14656 16088 14720
rect 16152 14656 16160 14720
rect 15840 13632 16160 14656
rect 15840 13568 15848 13632
rect 15912 13568 15928 13632
rect 15992 13568 16008 13632
rect 16072 13568 16088 13632
rect 16152 13568 16160 13632
rect 15840 12544 16160 13568
rect 15840 12480 15848 12544
rect 15912 12480 15928 12544
rect 15992 12480 16008 12544
rect 16072 12480 16088 12544
rect 16152 12480 16160 12544
rect 15840 11456 16160 12480
rect 15840 11392 15848 11456
rect 15912 11392 15928 11456
rect 15992 11392 16008 11456
rect 16072 11392 16088 11456
rect 16152 11392 16160 11456
rect 15840 10368 16160 11392
rect 15840 10304 15848 10368
rect 15912 10304 15928 10368
rect 15992 10304 16008 10368
rect 16072 10304 16088 10368
rect 16152 10304 16160 10368
rect 15840 9280 16160 10304
rect 15840 9216 15848 9280
rect 15912 9216 15928 9280
rect 15992 9216 16008 9280
rect 16072 9216 16088 9280
rect 16152 9216 16160 9280
rect 15840 8192 16160 9216
rect 15840 8128 15848 8192
rect 15912 8128 15928 8192
rect 15992 8128 16008 8192
rect 16072 8128 16088 8192
rect 16152 8128 16160 8192
rect 15840 7104 16160 8128
rect 15840 7040 15848 7104
rect 15912 7040 15928 7104
rect 15992 7040 16008 7104
rect 16072 7040 16088 7104
rect 16152 7040 16160 7104
rect 15840 6016 16160 7040
rect 15840 5952 15848 6016
rect 15912 5952 15928 6016
rect 15992 5952 16008 6016
rect 16072 5952 16088 6016
rect 16152 5952 16160 6016
rect 15840 4928 16160 5952
rect 15840 4864 15848 4928
rect 15912 4864 15928 4928
rect 15992 4864 16008 4928
rect 16072 4864 16088 4928
rect 16152 4864 16160 4928
rect 15840 3840 16160 4864
rect 15840 3776 15848 3840
rect 15912 3776 15928 3840
rect 15992 3776 16008 3840
rect 16072 3776 16088 3840
rect 16152 3776 16160 3840
rect 15840 2752 16160 3776
rect 15840 2688 15848 2752
rect 15912 2688 15928 2752
rect 15992 2688 16008 2752
rect 16072 2688 16088 2752
rect 16152 2688 16160 2752
rect 15840 2128 16160 2688
rect 20805 15264 21125 16288
rect 25638 15333 25698 18123
rect 25770 17984 26091 19008
rect 26190 18733 26250 22747
rect 26374 20773 26434 27235
rect 26558 25805 26618 32131
rect 26742 29749 26802 37027
rect 26926 32605 26986 37435
rect 27107 33556 27173 33557
rect 27107 33492 27108 33556
rect 27172 33492 27173 33556
rect 27107 33491 27173 33492
rect 26923 32604 26989 32605
rect 26923 32540 26924 32604
rect 26988 32540 26989 32604
rect 26923 32539 26989 32540
rect 26923 32468 26989 32469
rect 26923 32404 26924 32468
rect 26988 32404 26989 32468
rect 26923 32403 26989 32404
rect 26739 29748 26805 29749
rect 26739 29684 26740 29748
rect 26804 29684 26805 29748
rect 26739 29683 26805 29684
rect 26739 29612 26805 29613
rect 26739 29548 26740 29612
rect 26804 29548 26805 29612
rect 26739 29547 26805 29548
rect 26555 25804 26621 25805
rect 26555 25740 26556 25804
rect 26620 25740 26621 25804
rect 26555 25739 26621 25740
rect 26742 24037 26802 29547
rect 26926 27437 26986 32403
rect 27110 31789 27170 33491
rect 27291 32332 27357 32333
rect 27291 32268 27292 32332
rect 27356 32268 27357 32332
rect 27291 32267 27357 32268
rect 27107 31788 27173 31789
rect 27107 31724 27108 31788
rect 27172 31724 27173 31788
rect 27107 31723 27173 31724
rect 27107 29884 27173 29885
rect 27107 29820 27108 29884
rect 27172 29820 27173 29884
rect 27107 29819 27173 29820
rect 26923 27436 26989 27437
rect 26923 27372 26924 27436
rect 26988 27372 26989 27436
rect 26923 27371 26989 27372
rect 26739 24036 26805 24037
rect 26739 23972 26740 24036
rect 26804 23972 26805 24036
rect 26739 23971 26805 23972
rect 26742 22133 26802 23971
rect 27110 22133 27170 29819
rect 27294 29205 27354 32267
rect 27478 31109 27538 37707
rect 27662 32197 27722 40835
rect 27659 32196 27725 32197
rect 27659 32132 27660 32196
rect 27724 32132 27725 32196
rect 27659 32131 27725 32132
rect 27659 32060 27725 32061
rect 27659 31996 27660 32060
rect 27724 31996 27725 32060
rect 27659 31995 27725 31996
rect 27662 31517 27722 31995
rect 27659 31516 27725 31517
rect 27659 31452 27660 31516
rect 27724 31452 27725 31516
rect 27659 31451 27725 31452
rect 27659 31380 27725 31381
rect 27659 31316 27660 31380
rect 27724 31316 27725 31380
rect 27659 31315 27725 31316
rect 27475 31108 27541 31109
rect 27475 31044 27476 31108
rect 27540 31044 27541 31108
rect 27475 31043 27541 31044
rect 27475 30972 27541 30973
rect 27475 30908 27476 30972
rect 27540 30908 27541 30972
rect 27475 30907 27541 30908
rect 27291 29204 27357 29205
rect 27291 29140 27292 29204
rect 27356 29140 27357 29204
rect 27291 29139 27357 29140
rect 27291 27028 27357 27029
rect 27291 26964 27292 27028
rect 27356 26964 27357 27028
rect 27291 26963 27357 26964
rect 27294 25261 27354 26963
rect 27291 25260 27357 25261
rect 27291 25196 27292 25260
rect 27356 25196 27357 25260
rect 27291 25195 27357 25196
rect 27478 23901 27538 30907
rect 27662 26621 27722 31315
rect 27659 26620 27725 26621
rect 27659 26556 27660 26620
rect 27724 26556 27725 26620
rect 27659 26555 27725 26556
rect 27475 23900 27541 23901
rect 27475 23836 27476 23900
rect 27540 23836 27541 23900
rect 27475 23835 27541 23836
rect 26739 22132 26805 22133
rect 26739 22068 26740 22132
rect 26804 22068 26805 22132
rect 26739 22067 26805 22068
rect 27107 22132 27173 22133
rect 27107 22068 27108 22132
rect 27172 22068 27173 22132
rect 27107 22067 27173 22068
rect 27846 21997 27906 46139
rect 28214 45933 28274 55251
rect 28579 54636 28645 54637
rect 28579 54572 28580 54636
rect 28644 54572 28645 54636
rect 28579 54571 28645 54572
rect 28395 53412 28461 53413
rect 28395 53348 28396 53412
rect 28460 53348 28461 53412
rect 28395 53347 28461 53348
rect 28398 52733 28458 53347
rect 28395 52732 28461 52733
rect 28395 52668 28396 52732
rect 28460 52668 28461 52732
rect 28395 52667 28461 52668
rect 28395 51236 28461 51237
rect 28395 51172 28396 51236
rect 28460 51172 28461 51236
rect 28395 51171 28461 51172
rect 28211 45932 28277 45933
rect 28211 45868 28212 45932
rect 28276 45868 28277 45932
rect 28211 45867 28277 45868
rect 28211 41716 28277 41717
rect 28211 41652 28212 41716
rect 28276 41652 28277 41716
rect 28211 41651 28277 41652
rect 28027 41308 28093 41309
rect 28027 41244 28028 41308
rect 28092 41244 28093 41308
rect 28027 41243 28093 41244
rect 28030 38453 28090 41243
rect 28027 38452 28093 38453
rect 28027 38388 28028 38452
rect 28092 38388 28093 38452
rect 28027 38387 28093 38388
rect 28027 38180 28093 38181
rect 28027 38116 28028 38180
rect 28092 38116 28093 38180
rect 28027 38115 28093 38116
rect 28030 28933 28090 38115
rect 28214 31925 28274 41651
rect 28211 31924 28277 31925
rect 28211 31860 28212 31924
rect 28276 31860 28277 31924
rect 28211 31859 28277 31860
rect 28211 29884 28277 29885
rect 28211 29820 28212 29884
rect 28276 29820 28277 29884
rect 28211 29819 28277 29820
rect 28027 28932 28093 28933
rect 28027 28868 28028 28932
rect 28092 28868 28093 28932
rect 28027 28867 28093 28868
rect 28027 26756 28093 26757
rect 28027 26692 28028 26756
rect 28092 26692 28093 26756
rect 28027 26691 28093 26692
rect 28030 23765 28090 26691
rect 28214 25941 28274 29819
rect 28211 25940 28277 25941
rect 28211 25876 28212 25940
rect 28276 25876 28277 25940
rect 28211 25875 28277 25876
rect 28027 23764 28093 23765
rect 28027 23700 28028 23764
rect 28092 23700 28093 23764
rect 28027 23699 28093 23700
rect 27843 21996 27909 21997
rect 27843 21932 27844 21996
rect 27908 21932 27909 21996
rect 27843 21931 27909 21932
rect 26371 20772 26437 20773
rect 26371 20708 26372 20772
rect 26436 20708 26437 20772
rect 26371 20707 26437 20708
rect 26187 18732 26253 18733
rect 26187 18668 26188 18732
rect 26252 18668 26253 18732
rect 26187 18667 26253 18668
rect 25770 17920 25778 17984
rect 25842 17920 25858 17984
rect 25922 17920 25938 17984
rect 26002 17920 26018 17984
rect 26082 17920 26091 17984
rect 25770 16896 26091 17920
rect 26187 17644 26253 17645
rect 26187 17580 26188 17644
rect 26252 17580 26253 17644
rect 26187 17579 26253 17580
rect 25770 16832 25778 16896
rect 25842 16832 25858 16896
rect 25922 16832 25938 16896
rect 26002 16832 26018 16896
rect 26082 16832 26091 16896
rect 25770 15808 26091 16832
rect 25770 15744 25778 15808
rect 25842 15744 25858 15808
rect 25922 15744 25938 15808
rect 26002 15744 26018 15808
rect 26082 15744 26091 15808
rect 25635 15332 25701 15333
rect 25635 15268 25636 15332
rect 25700 15268 25701 15332
rect 25635 15267 25701 15268
rect 20805 15200 20813 15264
rect 20877 15200 20893 15264
rect 20957 15200 20973 15264
rect 21037 15200 21053 15264
rect 21117 15200 21125 15264
rect 20805 14176 21125 15200
rect 20805 14112 20813 14176
rect 20877 14112 20893 14176
rect 20957 14112 20973 14176
rect 21037 14112 21053 14176
rect 21117 14112 21125 14176
rect 20805 13088 21125 14112
rect 20805 13024 20813 13088
rect 20877 13024 20893 13088
rect 20957 13024 20973 13088
rect 21037 13024 21053 13088
rect 21117 13024 21125 13088
rect 20805 12000 21125 13024
rect 20805 11936 20813 12000
rect 20877 11936 20893 12000
rect 20957 11936 20973 12000
rect 21037 11936 21053 12000
rect 21117 11936 21125 12000
rect 20805 10912 21125 11936
rect 20805 10848 20813 10912
rect 20877 10848 20893 10912
rect 20957 10848 20973 10912
rect 21037 10848 21053 10912
rect 21117 10848 21125 10912
rect 20805 9824 21125 10848
rect 20805 9760 20813 9824
rect 20877 9760 20893 9824
rect 20957 9760 20973 9824
rect 21037 9760 21053 9824
rect 21117 9760 21125 9824
rect 20805 8736 21125 9760
rect 20805 8672 20813 8736
rect 20877 8672 20893 8736
rect 20957 8672 20973 8736
rect 21037 8672 21053 8736
rect 21117 8672 21125 8736
rect 20805 7648 21125 8672
rect 20805 7584 20813 7648
rect 20877 7584 20893 7648
rect 20957 7584 20973 7648
rect 21037 7584 21053 7648
rect 21117 7584 21125 7648
rect 20805 6560 21125 7584
rect 20805 6496 20813 6560
rect 20877 6496 20893 6560
rect 20957 6496 20973 6560
rect 21037 6496 21053 6560
rect 21117 6496 21125 6560
rect 20805 5472 21125 6496
rect 20805 5408 20813 5472
rect 20877 5408 20893 5472
rect 20957 5408 20973 5472
rect 21037 5408 21053 5472
rect 21117 5408 21125 5472
rect 20805 4384 21125 5408
rect 20805 4320 20813 4384
rect 20877 4320 20893 4384
rect 20957 4320 20973 4384
rect 21037 4320 21053 4384
rect 21117 4320 21125 4384
rect 20805 3296 21125 4320
rect 20805 3232 20813 3296
rect 20877 3232 20893 3296
rect 20957 3232 20973 3296
rect 21037 3232 21053 3296
rect 21117 3232 21125 3296
rect 20805 2208 21125 3232
rect 20805 2144 20813 2208
rect 20877 2144 20893 2208
rect 20957 2144 20973 2208
rect 21037 2144 21053 2208
rect 21117 2144 21125 2208
rect 20805 2128 21125 2144
rect 25770 14720 26091 15744
rect 25770 14656 25778 14720
rect 25842 14656 25858 14720
rect 25922 14656 25938 14720
rect 26002 14656 26018 14720
rect 26082 14656 26091 14720
rect 25770 13632 26091 14656
rect 25770 13568 25778 13632
rect 25842 13568 25858 13632
rect 25922 13568 25938 13632
rect 26002 13568 26018 13632
rect 26082 13568 26091 13632
rect 25770 12544 26091 13568
rect 25770 12480 25778 12544
rect 25842 12480 25858 12544
rect 25922 12480 25938 12544
rect 26002 12480 26018 12544
rect 26082 12480 26091 12544
rect 25770 11456 26091 12480
rect 26190 12069 26250 17579
rect 28398 15197 28458 51171
rect 28582 18733 28642 54571
rect 28766 54093 28826 58651
rect 29134 56813 29194 61102
rect 29499 61100 29500 61164
rect 29564 61100 29565 61164
rect 29499 61099 29565 61100
rect 29315 60484 29381 60485
rect 29315 60420 29316 60484
rect 29380 60420 29381 60484
rect 29315 60419 29381 60420
rect 29131 56812 29197 56813
rect 29131 56748 29132 56812
rect 29196 56748 29197 56812
rect 29131 56747 29197 56748
rect 28763 54092 28829 54093
rect 28763 54028 28764 54092
rect 28828 54028 28829 54092
rect 28763 54027 28829 54028
rect 28947 53412 29013 53413
rect 28947 53348 28948 53412
rect 29012 53348 29013 53412
rect 28947 53347 29013 53348
rect 28763 53140 28829 53141
rect 28763 53076 28764 53140
rect 28828 53076 28829 53140
rect 28763 53075 28829 53076
rect 28766 52461 28826 53075
rect 28763 52460 28829 52461
rect 28763 52396 28764 52460
rect 28828 52396 28829 52460
rect 28763 52395 28829 52396
rect 28766 48381 28826 52395
rect 28950 52189 29010 53347
rect 29318 53141 29378 60419
rect 29502 56949 29562 61099
rect 29683 59804 29749 59805
rect 29683 59740 29684 59804
rect 29748 59740 29749 59804
rect 29683 59739 29749 59740
rect 29499 56948 29565 56949
rect 29499 56884 29500 56948
rect 29564 56884 29565 56948
rect 29499 56883 29565 56884
rect 29499 53684 29565 53685
rect 29499 53620 29500 53684
rect 29564 53620 29565 53684
rect 29499 53619 29565 53620
rect 29315 53140 29381 53141
rect 29315 53076 29316 53140
rect 29380 53076 29381 53140
rect 29315 53075 29381 53076
rect 29315 52596 29381 52597
rect 29315 52532 29316 52596
rect 29380 52532 29381 52596
rect 29315 52531 29381 52532
rect 28947 52188 29013 52189
rect 28947 52124 28948 52188
rect 29012 52124 29013 52188
rect 28947 52123 29013 52124
rect 29318 51373 29378 52531
rect 29315 51372 29381 51373
rect 29315 51308 29316 51372
rect 29380 51308 29381 51372
rect 29315 51307 29381 51308
rect 29131 51100 29197 51101
rect 29131 51036 29132 51100
rect 29196 51036 29197 51100
rect 29131 51035 29197 51036
rect 28947 48516 29013 48517
rect 28947 48452 28948 48516
rect 29012 48452 29013 48516
rect 28947 48451 29013 48452
rect 28763 48380 28829 48381
rect 28763 48316 28764 48380
rect 28828 48316 28829 48380
rect 28763 48315 28829 48316
rect 28763 47972 28829 47973
rect 28763 47908 28764 47972
rect 28828 47908 28829 47972
rect 28763 47907 28829 47908
rect 28766 44573 28826 47907
rect 28950 46205 29010 48451
rect 28947 46204 29013 46205
rect 28947 46140 28948 46204
rect 29012 46140 29013 46204
rect 28947 46139 29013 46140
rect 28947 45660 29013 45661
rect 28947 45596 28948 45660
rect 29012 45596 29013 45660
rect 28947 45595 29013 45596
rect 28763 44572 28829 44573
rect 28763 44508 28764 44572
rect 28828 44508 28829 44572
rect 28763 44507 28829 44508
rect 28763 44300 28829 44301
rect 28763 44236 28764 44300
rect 28828 44236 28829 44300
rect 28763 44235 28829 44236
rect 28579 18732 28645 18733
rect 28579 18668 28580 18732
rect 28644 18668 28645 18732
rect 28579 18667 28645 18668
rect 28395 15196 28461 15197
rect 28395 15132 28396 15196
rect 28460 15132 28461 15196
rect 28395 15131 28461 15132
rect 26187 12068 26253 12069
rect 26187 12004 26188 12068
rect 26252 12004 26253 12068
rect 26187 12003 26253 12004
rect 25770 11392 25778 11456
rect 25842 11392 25858 11456
rect 25922 11392 25938 11456
rect 26002 11392 26018 11456
rect 26082 11392 26091 11456
rect 25770 10368 26091 11392
rect 25770 10304 25778 10368
rect 25842 10304 25858 10368
rect 25922 10304 25938 10368
rect 26002 10304 26018 10368
rect 26082 10304 26091 10368
rect 25770 9280 26091 10304
rect 25770 9216 25778 9280
rect 25842 9216 25858 9280
rect 25922 9216 25938 9280
rect 26002 9216 26018 9280
rect 26082 9216 26091 9280
rect 25770 8192 26091 9216
rect 25770 8128 25778 8192
rect 25842 8128 25858 8192
rect 25922 8128 25938 8192
rect 26002 8128 26018 8192
rect 26082 8128 26091 8192
rect 25770 7104 26091 8128
rect 25770 7040 25778 7104
rect 25842 7040 25858 7104
rect 25922 7040 25938 7104
rect 26002 7040 26018 7104
rect 26082 7040 26091 7104
rect 25770 6016 26091 7040
rect 25770 5952 25778 6016
rect 25842 5952 25858 6016
rect 25922 5952 25938 6016
rect 26002 5952 26018 6016
rect 26082 5952 26091 6016
rect 25770 4928 26091 5952
rect 25770 4864 25778 4928
rect 25842 4864 25858 4928
rect 25922 4864 25938 4928
rect 26002 4864 26018 4928
rect 26082 4864 26091 4928
rect 25770 3840 26091 4864
rect 28766 4725 28826 44235
rect 28950 30973 29010 45595
rect 29134 42397 29194 51035
rect 29315 48380 29381 48381
rect 29315 48316 29316 48380
rect 29380 48316 29381 48380
rect 29315 48315 29381 48316
rect 29131 42396 29197 42397
rect 29131 42332 29132 42396
rect 29196 42332 29197 42396
rect 29131 42331 29197 42332
rect 29131 42260 29197 42261
rect 29131 42196 29132 42260
rect 29196 42196 29197 42260
rect 29131 42195 29197 42196
rect 29134 41037 29194 42195
rect 29131 41036 29197 41037
rect 29131 40972 29132 41036
rect 29196 40972 29197 41036
rect 29131 40971 29197 40972
rect 29131 39404 29197 39405
rect 29131 39340 29132 39404
rect 29196 39340 29197 39404
rect 29131 39339 29197 39340
rect 29134 32877 29194 39339
rect 29131 32876 29197 32877
rect 29131 32812 29132 32876
rect 29196 32812 29197 32876
rect 29131 32811 29197 32812
rect 29131 32740 29197 32741
rect 29131 32676 29132 32740
rect 29196 32676 29197 32740
rect 29131 32675 29197 32676
rect 28947 30972 29013 30973
rect 28947 30908 28948 30972
rect 29012 30908 29013 30972
rect 28947 30907 29013 30908
rect 28947 30836 29013 30837
rect 28947 30772 28948 30836
rect 29012 30772 29013 30836
rect 28947 30771 29013 30772
rect 28950 25941 29010 30771
rect 29134 27845 29194 32675
rect 29131 27844 29197 27845
rect 29131 27780 29132 27844
rect 29196 27780 29197 27844
rect 29131 27779 29197 27780
rect 28947 25940 29013 25941
rect 28947 25876 28948 25940
rect 29012 25876 29013 25940
rect 28947 25875 29013 25876
rect 29131 21996 29197 21997
rect 29131 21932 29132 21996
rect 29196 21932 29197 21996
rect 29131 21931 29197 21932
rect 29134 18189 29194 21931
rect 29131 18188 29197 18189
rect 29131 18124 29132 18188
rect 29196 18124 29197 18188
rect 29131 18123 29197 18124
rect 29318 14109 29378 48315
rect 29502 15469 29562 53619
rect 29686 51373 29746 59739
rect 29867 57900 29933 57901
rect 29867 57836 29868 57900
rect 29932 57836 29933 57900
rect 29867 57835 29933 57836
rect 29870 51781 29930 57835
rect 30051 57220 30117 57221
rect 30051 57156 30052 57220
rect 30116 57156 30117 57220
rect 30051 57155 30117 57156
rect 30603 57220 30669 57221
rect 30603 57156 30604 57220
rect 30668 57156 30669 57220
rect 30603 57155 30669 57156
rect 30054 55045 30114 57155
rect 30051 55044 30117 55045
rect 30051 54980 30052 55044
rect 30116 54980 30117 55044
rect 30051 54979 30117 54980
rect 29867 51780 29933 51781
rect 29867 51716 29868 51780
rect 29932 51716 29933 51780
rect 29867 51715 29933 51716
rect 29867 51644 29933 51645
rect 29867 51580 29868 51644
rect 29932 51580 29933 51644
rect 29867 51579 29933 51580
rect 29683 51372 29749 51373
rect 29683 51308 29684 51372
rect 29748 51308 29749 51372
rect 29683 51307 29749 51308
rect 29870 50826 29930 51579
rect 30054 51237 30114 54979
rect 30235 53548 30301 53549
rect 30235 53484 30236 53548
rect 30300 53484 30301 53548
rect 30235 53483 30301 53484
rect 30238 52189 30298 53483
rect 30419 52732 30485 52733
rect 30419 52668 30420 52732
rect 30484 52668 30485 52732
rect 30419 52667 30485 52668
rect 30235 52188 30301 52189
rect 30235 52124 30236 52188
rect 30300 52124 30301 52188
rect 30235 52123 30301 52124
rect 30051 51236 30117 51237
rect 30051 51172 30052 51236
rect 30116 51172 30117 51236
rect 30051 51171 30117 51172
rect 30422 51090 30482 52667
rect 29686 50766 29930 50826
rect 30054 51030 30482 51090
rect 29686 48517 29746 50766
rect 29867 50692 29933 50693
rect 29867 50628 29868 50692
rect 29932 50690 29933 50692
rect 30054 50690 30114 51030
rect 30419 50964 30485 50965
rect 30419 50900 30420 50964
rect 30484 50900 30485 50964
rect 30419 50899 30485 50900
rect 29932 50630 30114 50690
rect 29932 50628 29933 50630
rect 29867 50627 29933 50628
rect 29683 48516 29749 48517
rect 29683 48452 29684 48516
rect 29748 48452 29749 48516
rect 29683 48451 29749 48452
rect 29683 44300 29749 44301
rect 29683 44236 29684 44300
rect 29748 44236 29749 44300
rect 29683 44235 29749 44236
rect 29499 15468 29565 15469
rect 29499 15404 29500 15468
rect 29564 15404 29565 15468
rect 29499 15403 29565 15404
rect 29315 14108 29381 14109
rect 29315 14044 29316 14108
rect 29380 14044 29381 14108
rect 29315 14043 29381 14044
rect 29686 5405 29746 44235
rect 29870 43077 29930 50627
rect 30051 50420 30117 50421
rect 30051 50356 30052 50420
rect 30116 50356 30117 50420
rect 30051 50355 30117 50356
rect 30054 47429 30114 50355
rect 30422 50010 30482 50899
rect 30606 50285 30666 57155
rect 30787 55724 30853 55725
rect 30787 55660 30788 55724
rect 30852 55660 30853 55724
rect 30787 55659 30853 55660
rect 30790 53141 30850 55659
rect 31523 54500 31589 54501
rect 31523 54436 31524 54500
rect 31588 54436 31589 54500
rect 31523 54435 31589 54436
rect 30787 53140 30853 53141
rect 30787 53076 30788 53140
rect 30852 53076 30853 53140
rect 30787 53075 30853 53076
rect 30787 51236 30853 51237
rect 30787 51172 30788 51236
rect 30852 51172 30853 51236
rect 30787 51171 30853 51172
rect 31155 51236 31221 51237
rect 31155 51172 31156 51236
rect 31220 51172 31221 51236
rect 31155 51171 31221 51172
rect 30790 50693 30850 51171
rect 31158 51090 31218 51171
rect 30974 51030 31218 51090
rect 30974 50965 31034 51030
rect 30971 50964 31037 50965
rect 30971 50900 30972 50964
rect 31036 50900 31037 50964
rect 30971 50899 31037 50900
rect 30787 50692 30853 50693
rect 30787 50628 30788 50692
rect 30852 50628 30853 50692
rect 30787 50627 30853 50628
rect 30603 50284 30669 50285
rect 30603 50220 30604 50284
rect 30668 50220 30669 50284
rect 30603 50219 30669 50220
rect 30238 49950 30482 50010
rect 30051 47428 30117 47429
rect 30051 47364 30052 47428
rect 30116 47364 30117 47428
rect 30051 47363 30117 47364
rect 30238 46069 30298 49950
rect 30419 49468 30485 49469
rect 30419 49404 30420 49468
rect 30484 49404 30485 49468
rect 30419 49403 30485 49404
rect 30235 46068 30301 46069
rect 30235 46004 30236 46068
rect 30300 46004 30301 46068
rect 30235 46003 30301 46004
rect 30235 44572 30301 44573
rect 30235 44508 30236 44572
rect 30300 44508 30301 44572
rect 30235 44507 30301 44508
rect 30238 43346 30298 44507
rect 30422 43349 30482 49403
rect 31155 49332 31221 49333
rect 31155 49268 31156 49332
rect 31220 49268 31221 49332
rect 31155 49267 31221 49268
rect 31158 48650 31218 49267
rect 31158 48590 31402 48650
rect 30787 47292 30853 47293
rect 30787 47228 30788 47292
rect 30852 47228 30853 47292
rect 30787 47227 30853 47228
rect 30603 46476 30669 46477
rect 30603 46412 30604 46476
rect 30668 46412 30669 46476
rect 30603 46411 30669 46412
rect 30192 43286 30298 43346
rect 30419 43348 30485 43349
rect 29867 43076 29933 43077
rect 29867 43012 29868 43076
rect 29932 43012 29933 43076
rect 29867 43011 29933 43012
rect 30051 43076 30117 43077
rect 30051 43012 30052 43076
rect 30116 43012 30117 43076
rect 30192 43074 30252 43286
rect 30419 43284 30420 43348
rect 30484 43284 30485 43348
rect 30419 43283 30485 43284
rect 30419 43076 30485 43077
rect 30192 43014 30298 43074
rect 30051 43011 30117 43012
rect 29867 42804 29933 42805
rect 29867 42740 29868 42804
rect 29932 42740 29933 42804
rect 29867 42739 29933 42740
rect 29683 5404 29749 5405
rect 29683 5340 29684 5404
rect 29748 5340 29749 5404
rect 29683 5339 29749 5340
rect 28763 4724 28829 4725
rect 28763 4660 28764 4724
rect 28828 4660 28829 4724
rect 28763 4659 28829 4660
rect 29870 4045 29930 42739
rect 30054 41717 30114 43011
rect 30051 41716 30117 41717
rect 30051 41652 30052 41716
rect 30116 41652 30117 41716
rect 30051 41651 30117 41652
rect 30051 40492 30117 40493
rect 30051 40428 30052 40492
rect 30116 40428 30117 40492
rect 30051 40427 30117 40428
rect 30054 36685 30114 40427
rect 30051 36684 30117 36685
rect 30051 36620 30052 36684
rect 30116 36620 30117 36684
rect 30051 36619 30117 36620
rect 30238 34530 30298 43014
rect 30419 43012 30420 43076
rect 30484 43012 30485 43076
rect 30419 43011 30485 43012
rect 30422 39405 30482 43011
rect 30606 42122 30666 46411
rect 30790 43213 30850 47227
rect 31342 44190 31402 48590
rect 31526 48381 31586 54435
rect 31523 48380 31589 48381
rect 31523 48316 31524 48380
rect 31588 48316 31589 48380
rect 31523 48315 31589 48316
rect 31891 47428 31957 47429
rect 31891 47364 31892 47428
rect 31956 47364 31957 47428
rect 31891 47363 31957 47364
rect 31523 46476 31589 46477
rect 31523 46412 31524 46476
rect 31588 46412 31589 46476
rect 31523 46411 31589 46412
rect 31526 45117 31586 46411
rect 31523 45116 31589 45117
rect 31523 45052 31524 45116
rect 31588 45052 31589 45116
rect 31523 45051 31589 45052
rect 31342 44130 31586 44190
rect 30971 43620 31037 43621
rect 30971 43556 30972 43620
rect 31036 43556 31037 43620
rect 30971 43555 31037 43556
rect 30787 43212 30853 43213
rect 30787 43148 30788 43212
rect 30852 43148 30853 43212
rect 30974 43210 31034 43555
rect 31339 43212 31405 43213
rect 30974 43150 31218 43210
rect 30787 43147 30853 43148
rect 30971 42668 31037 42669
rect 30971 42604 30972 42668
rect 31036 42604 31037 42668
rect 30971 42603 31037 42604
rect 30606 42062 30850 42122
rect 30790 41717 30850 42062
rect 30787 41716 30853 41717
rect 30787 41652 30788 41716
rect 30852 41652 30853 41716
rect 30787 41651 30853 41652
rect 30787 41580 30853 41581
rect 30787 41516 30788 41580
rect 30852 41516 30853 41580
rect 30787 41515 30853 41516
rect 30603 41172 30669 41173
rect 30603 41108 30604 41172
rect 30668 41108 30669 41172
rect 30603 41107 30669 41108
rect 30419 39404 30485 39405
rect 30419 39340 30420 39404
rect 30484 39340 30485 39404
rect 30419 39339 30485 39340
rect 30419 38996 30485 38997
rect 30419 38932 30420 38996
rect 30484 38932 30485 38996
rect 30419 38931 30485 38932
rect 30422 37229 30482 38931
rect 30419 37228 30485 37229
rect 30419 37164 30420 37228
rect 30484 37164 30485 37228
rect 30419 37163 30485 37164
rect 30054 34470 30298 34530
rect 30054 6493 30114 34470
rect 30235 34236 30301 34237
rect 30235 34172 30236 34236
rect 30300 34172 30301 34236
rect 30235 34171 30301 34172
rect 30238 24853 30298 34171
rect 30419 31924 30485 31925
rect 30419 31860 30420 31924
rect 30484 31860 30485 31924
rect 30419 31859 30485 31860
rect 30422 31650 30482 31859
rect 30606 31789 30666 41107
rect 30790 40765 30850 41515
rect 30787 40764 30853 40765
rect 30787 40700 30788 40764
rect 30852 40700 30853 40764
rect 30787 40699 30853 40700
rect 30787 39948 30853 39949
rect 30787 39884 30788 39948
rect 30852 39884 30853 39948
rect 30787 39883 30853 39884
rect 30603 31788 30669 31789
rect 30603 31724 30604 31788
rect 30668 31724 30669 31788
rect 30603 31723 30669 31724
rect 30422 31590 30666 31650
rect 30419 31380 30485 31381
rect 30419 31316 30420 31380
rect 30484 31316 30485 31380
rect 30419 31315 30485 31316
rect 30235 24852 30301 24853
rect 30235 24788 30236 24852
rect 30300 24788 30301 24852
rect 30235 24787 30301 24788
rect 30422 22810 30482 31315
rect 30606 31109 30666 31590
rect 30603 31108 30669 31109
rect 30603 31044 30604 31108
rect 30668 31044 30669 31108
rect 30603 31043 30669 31044
rect 30790 30429 30850 39883
rect 30974 36277 31034 42603
rect 31158 38045 31218 43150
rect 31339 43148 31340 43212
rect 31404 43148 31405 43212
rect 31339 43147 31405 43148
rect 31342 38045 31402 43147
rect 31155 38044 31221 38045
rect 31155 37980 31156 38044
rect 31220 37980 31221 38044
rect 31155 37979 31221 37980
rect 31339 38044 31405 38045
rect 31339 37980 31340 38044
rect 31404 37980 31405 38044
rect 31339 37979 31405 37980
rect 31155 37092 31221 37093
rect 31155 37028 31156 37092
rect 31220 37028 31221 37092
rect 31155 37027 31221 37028
rect 30971 36276 31037 36277
rect 30971 36212 30972 36276
rect 31036 36212 31037 36276
rect 30971 36211 31037 36212
rect 30971 32332 31037 32333
rect 30971 32268 30972 32332
rect 31036 32330 31037 32332
rect 31158 32330 31218 37027
rect 31526 36141 31586 44130
rect 31707 44164 31773 44165
rect 31707 44100 31708 44164
rect 31772 44100 31773 44164
rect 31707 44099 31773 44100
rect 31710 38997 31770 44099
rect 31894 39949 31954 47363
rect 31891 39948 31957 39949
rect 31891 39884 31892 39948
rect 31956 39884 31957 39948
rect 31891 39883 31957 39884
rect 31707 38996 31773 38997
rect 31707 38932 31708 38996
rect 31772 38932 31773 38996
rect 31707 38931 31773 38932
rect 31523 36140 31589 36141
rect 31523 36076 31524 36140
rect 31588 36076 31589 36140
rect 31523 36075 31589 36076
rect 31036 32270 31218 32330
rect 31036 32268 31037 32270
rect 30971 32267 31037 32268
rect 31155 31924 31221 31925
rect 31155 31860 31156 31924
rect 31220 31860 31221 31924
rect 31155 31859 31221 31860
rect 31158 30973 31218 31859
rect 31155 30972 31221 30973
rect 31155 30908 31156 30972
rect 31220 30908 31221 30972
rect 31155 30907 31221 30908
rect 30787 30428 30853 30429
rect 30787 30364 30788 30428
rect 30852 30364 30853 30428
rect 30787 30363 30853 30364
rect 30603 30020 30669 30021
rect 30603 29956 30604 30020
rect 30668 29956 30669 30020
rect 30603 29955 30669 29956
rect 30606 28797 30666 29955
rect 30603 28796 30669 28797
rect 30603 28732 30604 28796
rect 30668 28732 30669 28796
rect 30603 28731 30669 28732
rect 30238 22750 30482 22810
rect 30238 22133 30298 22750
rect 30419 22540 30485 22541
rect 30419 22476 30420 22540
rect 30484 22476 30485 22540
rect 30419 22475 30485 22476
rect 30235 22132 30301 22133
rect 30235 22068 30236 22132
rect 30300 22068 30301 22132
rect 30235 22067 30301 22068
rect 30422 19821 30482 22475
rect 30419 19820 30485 19821
rect 30419 19756 30420 19820
rect 30484 19756 30485 19820
rect 30419 19755 30485 19756
rect 30051 6492 30117 6493
rect 30051 6428 30052 6492
rect 30116 6428 30117 6492
rect 30051 6427 30117 6428
rect 29867 4044 29933 4045
rect 29867 3980 29868 4044
rect 29932 3980 29933 4044
rect 29867 3979 29933 3980
rect 25770 3776 25778 3840
rect 25842 3776 25858 3840
rect 25922 3776 25938 3840
rect 26002 3776 26018 3840
rect 26082 3776 26091 3840
rect 25770 2752 26091 3776
rect 25770 2688 25778 2752
rect 25842 2688 25858 2752
rect 25922 2688 25938 2752
rect 26002 2688 26018 2752
rect 26082 2688 26091 2752
rect 25770 2128 26091 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 28888 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 27968 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 28980 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 28980 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 27968 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 25300 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 28704 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform -1 0 28060 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform 1 0 28612 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1644511149
transform 1 0 28244 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1644511149
transform 1 0 27416 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1644511149
transform -1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1644511149
transform 1 0 27692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1644511149
transform 1 0 28980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1644511149
transform -1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1644511149
transform -1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1644511149
transform 1 0 1932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_296
timestamp 1644511149
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1644511149
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1644511149
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_301
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1644511149
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_316
timestamp 1644511149
transform 1 0 30176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp 1644511149
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_257
timestamp 1644511149
transform 1 0 24748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_274
timestamp 1644511149
transform 1 0 26312 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_286
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_292
timestamp 1644511149
transform 1 0 27968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_296
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_316
timestamp 1644511149
transform 1 0 30176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_23
timestamp 1644511149
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_35
timestamp 1644511149
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1644511149
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1644511149
transform 1 0 19136 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1644511149
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1644511149
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1644511149
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_287
timestamp 1644511149
transform 1 0 27508 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_291
timestamp 1644511149
transform 1 0 27876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_295
timestamp 1644511149
transform 1 0 28244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_301
timestamp 1644511149
transform 1 0 28796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_316
timestamp 1644511149
transform 1 0 30176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_7
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_241
timestamp 1644511149
transform 1 0 23276 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_259
timestamp 1644511149
transform 1 0 24932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_266
timestamp 1644511149
transform 1 0 25576 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_274
timestamp 1644511149
transform 1 0 26312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_282
timestamp 1644511149
transform 1 0 27048 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp 1644511149
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_316
timestamp 1644511149
transform 1 0 30176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1644511149
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_31
timestamp 1644511149
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1644511149
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_243
timestamp 1644511149
transform 1 0 23460 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_255
timestamp 1644511149
transform 1 0 24564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1644511149
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1644511149
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_286
timestamp 1644511149
transform 1 0 27416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_290
timestamp 1644511149
transform 1 0 27784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_295
timestamp 1644511149
transform 1 0 28244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_303
timestamp 1644511149
transform 1 0 28980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1644511149
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1644511149
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_261
timestamp 1644511149
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_270
timestamp 1644511149
transform 1 0 25944 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1644511149
transform 1 0 26496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_287
timestamp 1644511149
transform 1 0 27508 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_295
timestamp 1644511149
transform 1 0 28244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_316
timestamp 1644511149
transform 1 0 30176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_11
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_23
timestamp 1644511149
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_35
timestamp 1644511149
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1644511149
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_258
timestamp 1644511149
transform 1 0 24840 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_270
timestamp 1644511149
transform 1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1644511149
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_289
timestamp 1644511149
transform 1 0 27692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_303
timestamp 1644511149
transform 1 0 28980 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_316
timestamp 1644511149
transform 1 0 30176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_238
timestamp 1644511149
transform 1 0 23000 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1644511149
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_261
timestamp 1644511149
transform 1 0 25116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_271
timestamp 1644511149
transform 1 0 26036 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_282
timestamp 1644511149
transform 1 0 27048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1644511149
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_316
timestamp 1644511149
transform 1 0 30176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1644511149
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1644511149
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1644511149
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_256
timestamp 1644511149
transform 1 0 24656 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_268
timestamp 1644511149
transform 1 0 25760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_285
timestamp 1644511149
transform 1 0 27324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_291
timestamp 1644511149
transform 1 0 27876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_313
timestamp 1644511149
transform 1 0 29900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_319
timestamp 1644511149
transform 1 0 30452 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_14
timestamp 1644511149
transform 1 0 2392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1644511149
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_240
timestamp 1644511149
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_275
timestamp 1644511149
transform 1 0 26404 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_293
timestamp 1644511149
transform 1 0 28060 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_298
timestamp 1644511149
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1644511149
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_316
timestamp 1644511149
transform 1 0 30176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_19
timestamp 1644511149
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1644511149
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1644511149
transform 1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1644511149
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_269
timestamp 1644511149
transform 1 0 25852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_288
timestamp 1644511149
transform 1 0 27600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_313
timestamp 1644511149
transform 1 0 29900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_319
timestamp 1644511149
transform 1 0 30452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_14
timestamp 1644511149
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1644511149
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_205
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_210
timestamp 1644511149
transform 1 0 20424 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_238
timestamp 1644511149
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1644511149
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_271
timestamp 1644511149
transform 1 0 26036 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_279
timestamp 1644511149
transform 1 0 26772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_291
timestamp 1644511149
transform 1 0 27876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_316
timestamp 1644511149
transform 1 0 30176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_211
timestamp 1644511149
transform 1 0 20516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_233
timestamp 1644511149
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_240
timestamp 1644511149
transform 1 0 23184 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_248
timestamp 1644511149
transform 1 0 23920 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_253
timestamp 1644511149
transform 1 0 24380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1644511149
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_286
timestamp 1644511149
transform 1 0 27416 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_294
timestamp 1644511149
transform 1 0 28152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_316
timestamp 1644511149
transform 1 0 30176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_7
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_14
timestamp 1644511149
transform 1 0 2392 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1644511149
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_203
timestamp 1644511149
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_214
timestamp 1644511149
transform 1 0 20792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_227
timestamp 1644511149
transform 1 0 21988 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_241
timestamp 1644511149
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1644511149
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_271
timestamp 1644511149
transform 1 0 26036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1644511149
transform 1 0 26496 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_288
timestamp 1644511149
transform 1 0 27600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_294
timestamp 1644511149
transform 1 0 28152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1644511149
transform 1 0 28520 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1644511149
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_316
timestamp 1644511149
transform 1 0 30176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_19
timestamp 1644511149
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_31
timestamp 1644511149
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1644511149
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1644511149
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_202
timestamp 1644511149
transform 1 0 19688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_213
timestamp 1644511149
transform 1 0 20700 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_241
timestamp 1644511149
transform 1 0 23276 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_267
timestamp 1644511149
transform 1 0 25668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_271
timestamp 1644511149
transform 1 0 26036 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_291
timestamp 1644511149
transform 1 0 27876 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_316
timestamp 1644511149
transform 1 0 30176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_14
timestamp 1644511149
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_205
timestamp 1644511149
transform 1 0 19964 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_220
timestamp 1644511149
transform 1 0 21344 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_232
timestamp 1644511149
transform 1 0 22448 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1644511149
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_261
timestamp 1644511149
transform 1 0 25116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_269
timestamp 1644511149
transform 1 0 25852 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_275
timestamp 1644511149
transform 1 0 26404 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_280
timestamp 1644511149
transform 1 0 26864 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_296
timestamp 1644511149
transform 1 0 28336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1644511149
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1644511149
transform 1 0 30176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_19
timestamp 1644511149
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_31
timestamp 1644511149
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_43
timestamp 1644511149
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1644511149
transform 1 0 19320 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_255
timestamp 1644511149
transform 1 0 24564 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_262
timestamp 1644511149
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_266
timestamp 1644511149
transform 1 0 25576 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_302
timestamp 1644511149
transform 1 0 28888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_316
timestamp 1644511149
transform 1 0 30176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1644511149
transform 1 0 1748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_11
timestamp 1644511149
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1644511149
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_173
timestamp 1644511149
transform 1 0 17020 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1644511149
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1644511149
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1644511149
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_218
timestamp 1644511149
transform 1 0 21160 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_230
timestamp 1644511149
transform 1 0 22264 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1644511149
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1644511149
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_261
timestamp 1644511149
transform 1 0 25116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_269
timestamp 1644511149
transform 1 0 25852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_279
timestamp 1644511149
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1644511149
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_316
timestamp 1644511149
transform 1 0 30176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_233
timestamp 1644511149
transform 1 0 22540 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_241
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_253
timestamp 1644511149
transform 1 0 24380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_262
timestamp 1644511149
transform 1 0 25208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_289
timestamp 1644511149
transform 1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_302
timestamp 1644511149
transform 1 0 28888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 1644511149
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 1644511149
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_241
timestamp 1644511149
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1644511149
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_261
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_269
timestamp 1644511149
transform 1 0 25852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_278
timestamp 1644511149
transform 1 0 26680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_316
timestamp 1644511149
transform 1 0 30176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_7
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1644511149
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1644511149
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1644511149
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_242
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_254
timestamp 1644511149
transform 1 0 24472 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_289
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_302
timestamp 1644511149
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1644511149
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_7
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1644511149
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_205
timestamp 1644511149
transform 1 0 19964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1644511149
transform 1 0 20884 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_227
timestamp 1644511149
transform 1 0 21988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_231
timestamp 1644511149
transform 1 0 22356 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_238
timestamp 1644511149
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1644511149
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_281
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1644511149
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_316
timestamp 1644511149
transform 1 0 30176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1644511149
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1644511149
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1644511149
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_197
timestamp 1644511149
transform 1 0 19228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1644511149
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1644511149
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_241
timestamp 1644511149
transform 1 0 23276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_245
timestamp 1644511149
transform 1 0 23644 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_252
timestamp 1644511149
transform 1 0 24288 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_262
timestamp 1644511149
transform 1 0 25208 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_270
timestamp 1644511149
transform 1 0 25944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1644511149
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_299
timestamp 1644511149
transform 1 0 28612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1644511149
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_14
timestamp 1644511149
transform 1 0 2392 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1644511149
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1644511149
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_214
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_218
timestamp 1644511149
transform 1 0 21160 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_229
timestamp 1644511149
transform 1 0 22172 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_241
timestamp 1644511149
transform 1 0 23276 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1644511149
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_281
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_291
timestamp 1644511149
transform 1 0 27876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_299
timestamp 1644511149
transform 1 0 28612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_316
timestamp 1644511149
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1644511149
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_16
timestamp 1644511149
transform 1 0 2576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_28
timestamp 1644511149
transform 1 0 3680 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_40
timestamp 1644511149
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1644511149
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1644511149
transform 1 0 18308 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_199
timestamp 1644511149
transform 1 0 19412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1644511149
transform 1 0 20148 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1644511149
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1644511149
transform 1 0 22172 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_253
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_259
timestamp 1644511149
transform 1 0 24932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_291
timestamp 1644511149
transform 1 0 27876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_302
timestamp 1644511149
transform 1 0 28888 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_310
timestamp 1644511149
transform 1 0 29624 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1644511149
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_14
timestamp 1644511149
transform 1 0 2392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1644511149
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_161
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_176
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_205
timestamp 1644511149
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_216
timestamp 1644511149
transform 1 0 20976 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_228
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_240
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_286
timestamp 1644511149
transform 1 0 27416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1644511149
transform 1 0 27784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_316
timestamp 1644511149
transform 1 0 30176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_14
timestamp 1644511149
transform 1 0 2392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_26
timestamp 1644511149
transform 1 0 3496 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_38
timestamp 1644511149
transform 1 0 4600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1644511149
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_177
timestamp 1644511149
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_183
timestamp 1644511149
transform 1 0 17940 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_187
timestamp 1644511149
transform 1 0 18308 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_195
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_206
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1644511149
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_231
timestamp 1644511149
transform 1 0 22356 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_238
timestamp 1644511149
transform 1 0 23000 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_246
timestamp 1644511149
transform 1 0 23736 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_255
timestamp 1644511149
transform 1 0 24564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_267
timestamp 1644511149
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1644511149
transform 1 0 27784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_298
timestamp 1644511149
transform 1 0 28520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_304
timestamp 1644511149
transform 1 0 29072 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_308
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_316
timestamp 1644511149
transform 1 0 30176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1644511149
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_205
timestamp 1644511149
transform 1 0 19964 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_218
timestamp 1644511149
transform 1 0 21160 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_230
timestamp 1644511149
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_261
timestamp 1644511149
transform 1 0 25116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_273
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_293
timestamp 1644511149
transform 1 0 28060 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_297
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_316
timestamp 1644511149
transform 1 0 30176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_14
timestamp 1644511149
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1644511149
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1644511149
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_241
timestamp 1644511149
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_251
timestamp 1644511149
transform 1 0 24196 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_258
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1644511149
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_300
timestamp 1644511149
transform 1 0 28704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_304
timestamp 1644511149
transform 1 0 29072 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_314
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_9
timestamp 1644511149
transform 1 0 1932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_16
timestamp 1644511149
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_282
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_294
timestamp 1644511149
transform 1 0 28152 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_314
timestamp 1644511149
transform 1 0 29992 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_14
timestamp 1644511149
transform 1 0 2392 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_26
timestamp 1644511149
transform 1 0 3496 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_38
timestamp 1644511149
transform 1 0 4600 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1644511149
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_175
timestamp 1644511149
transform 1 0 17204 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_185
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_197
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_203
timestamp 1644511149
transform 1 0 19780 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_209
timestamp 1644511149
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1644511149
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_243
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1644511149
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_296
timestamp 1644511149
transform 1 0 28336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1644511149
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_14
timestamp 1644511149
transform 1 0 2392 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1644511149
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_172
timestamp 1644511149
transform 1 0 16928 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_212
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_224
timestamp 1644511149
transform 1 0 21712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_242
timestamp 1644511149
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1644511149
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_285
timestamp 1644511149
transform 1 0 27324 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_293
timestamp 1644511149
transform 1 0 28060 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1644511149
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_316
timestamp 1644511149
transform 1 0 30176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_7
timestamp 1644511149
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_19
timestamp 1644511149
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_31
timestamp 1644511149
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_43
timestamp 1644511149
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_185
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_209
timestamp 1644511149
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1644511149
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_298
timestamp 1644511149
transform 1 0 28520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_306
timestamp 1644511149
transform 1 0 29256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1644511149
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_7
timestamp 1644511149
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1644511149
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 1644511149
transform 1 0 16652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_174
timestamp 1644511149
transform 1 0 17112 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_183
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_213
timestamp 1644511149
transform 1 0 20700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_225
timestamp 1644511149
transform 1 0 21804 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1644511149
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1644511149
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_261
timestamp 1644511149
transform 1 0 25116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_273
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_296
timestamp 1644511149
transform 1 0 28336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_316
timestamp 1644511149
transform 1 0 30176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_14
timestamp 1644511149
transform 1 0 2392 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_26
timestamp 1644511149
transform 1 0 3496 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_38
timestamp 1644511149
transform 1 0 4600 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1644511149
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_172
timestamp 1644511149
transform 1 0 16928 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_180
timestamp 1644511149
transform 1 0 17664 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_185
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_200
timestamp 1644511149
transform 1 0 19504 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_212
timestamp 1644511149
transform 1 0 20608 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_257
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1644511149
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_300
timestamp 1644511149
transform 1 0 28704 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_307
timestamp 1644511149
transform 1 0 29348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_316
timestamp 1644511149
transform 1 0 30176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_9
timestamp 1644511149
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1644511149
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_205
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_217
timestamp 1644511149
transform 1 0 21068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_229
timestamp 1644511149
transform 1 0 22172 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_235
timestamp 1644511149
transform 1 0 22724 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_247
timestamp 1644511149
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_259
timestamp 1644511149
transform 1 0 24932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_276
timestamp 1644511149
transform 1 0 26496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_287
timestamp 1644511149
transform 1 0 27508 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_291
timestamp 1644511149
transform 1 0 27876 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1644511149
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_315
timestamp 1644511149
transform 1 0 30084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_319
timestamp 1644511149
transform 1 0 30452 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_14
timestamp 1644511149
transform 1 0 2392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_26
timestamp 1644511149
transform 1 0 3496 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_38
timestamp 1644511149
transform 1 0 4600 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_50
timestamp 1644511149
transform 1 0 5704 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_185
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_197
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_209
timestamp 1644511149
transform 1 0 20332 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_215
timestamp 1644511149
transform 1 0 20884 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_231
timestamp 1644511149
transform 1 0 22356 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_239
timestamp 1644511149
transform 1 0 23092 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_246
timestamp 1644511149
transform 1 0 23736 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_258
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_268
timestamp 1644511149
transform 1 0 25760 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_290
timestamp 1644511149
transform 1 0 27784 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_303
timestamp 1644511149
transform 1 0 28980 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_307
timestamp 1644511149
transform 1 0 29348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_313
timestamp 1644511149
transform 1 0 29900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_319
timestamp 1644511149
transform 1 0 30452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_14
timestamp 1644511149
transform 1 0 2392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1644511149
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_158
timestamp 1644511149
transform 1 0 15640 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_170
timestamp 1644511149
transform 1 0 16744 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_182
timestamp 1644511149
transform 1 0 17848 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1644511149
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_242
timestamp 1644511149
transform 1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1644511149
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_259
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_271
timestamp 1644511149
transform 1 0 26036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_283
timestamp 1644511149
transform 1 0 27140 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_291
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_296
timestamp 1644511149
transform 1 0 28336 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_314
timestamp 1644511149
transform 1 0 29992 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_14
timestamp 1644511149
transform 1 0 2392 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_26
timestamp 1644511149
transform 1 0 3496 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_38
timestamp 1644511149
transform 1 0 4600 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_50
timestamp 1644511149
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_134
timestamp 1644511149
transform 1 0 13432 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_146
timestamp 1644511149
transform 1 0 14536 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_158
timestamp 1644511149
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1644511149
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_183
timestamp 1644511149
transform 1 0 17940 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_195
timestamp 1644511149
transform 1 0 19044 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_199
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_203
timestamp 1644511149
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_215
timestamp 1644511149
transform 1 0 20884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_236
timestamp 1644511149
transform 1 0 22816 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_248
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_252
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_266
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1644511149
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_300
timestamp 1644511149
transform 1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_308
timestamp 1644511149
transform 1 0 29440 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_316
timestamp 1644511149
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_14
timestamp 1644511149
transform 1 0 2392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1644511149
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_156
timestamp 1644511149
transform 1 0 15456 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_164
timestamp 1644511149
transform 1 0 16192 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_183
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_204
timestamp 1644511149
transform 1 0 19872 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_212
timestamp 1644511149
transform 1 0 20608 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1644511149
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_226
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1644511149
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_261
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_269
timestamp 1644511149
transform 1 0 25852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_297
timestamp 1644511149
transform 1 0 28428 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_316
timestamp 1644511149
transform 1 0 30176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_7
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_14
timestamp 1644511149
transform 1 0 2392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_26
timestamp 1644511149
transform 1 0 3496 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_38
timestamp 1644511149
transform 1 0 4600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1644511149
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1644511149
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_156
timestamp 1644511149
transform 1 0 15456 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1644511149
transform 1 0 17572 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_200
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_235
timestamp 1644511149
transform 1 0 22724 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_248
timestamp 1644511149
transform 1 0 23920 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_258
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_262
timestamp 1644511149
transform 1 0 25208 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_287
timestamp 1644511149
transform 1 0 27508 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_298
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_306
timestamp 1644511149
transform 1 0 29256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_316
timestamp 1644511149
transform 1 0 30176 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_9
timestamp 1644511149
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_169
timestamp 1644511149
transform 1 0 16652 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_175
timestamp 1644511149
transform 1 0 17204 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_185
timestamp 1644511149
transform 1 0 18124 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_217
timestamp 1644511149
transform 1 0 21068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_236
timestamp 1644511149
transform 1 0 22816 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_260
timestamp 1644511149
transform 1 0 25024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_268
timestamp 1644511149
transform 1 0 25760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_280
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_288
timestamp 1644511149
transform 1 0 27600 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_297
timestamp 1644511149
transform 1 0 28428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_316
timestamp 1644511149
transform 1 0 30176 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_7
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_14
timestamp 1644511149
transform 1 0 2392 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_26
timestamp 1644511149
transform 1 0 3496 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_38
timestamp 1644511149
transform 1 0 4600 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1644511149
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_121
timestamp 1644511149
transform 1 0 12236 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_132
timestamp 1644511149
transform 1 0 13248 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_144
timestamp 1644511149
transform 1 0 14352 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_156
timestamp 1644511149
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_185
timestamp 1644511149
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_197
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_201
timestamp 1644511149
transform 1 0 19596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1644511149
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1644511149
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_229
timestamp 1644511149
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_289
timestamp 1644511149
transform 1 0 27692 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_295
timestamp 1644511149
transform 1 0 28244 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_301
timestamp 1644511149
transform 1 0 28796 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_316
timestamp 1644511149
transform 1 0 30176 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_14
timestamp 1644511149
transform 1 0 2392 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1644511149
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_129
timestamp 1644511149
transform 1 0 12972 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1644511149
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_157
timestamp 1644511149
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_175
timestamp 1644511149
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1644511149
transform 1 0 25944 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_282
timestamp 1644511149
transform 1 0 27048 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_290
timestamp 1644511149
transform 1 0 27784 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_296
timestamp 1644511149
transform 1 0 28336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_316
timestamp 1644511149
transform 1 0 30176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_7
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_14
timestamp 1644511149
transform 1 0 2392 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_26
timestamp 1644511149
transform 1 0 3496 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_38
timestamp 1644511149
transform 1 0 4600 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_50
timestamp 1644511149
transform 1 0 5704 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_133
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_138
timestamp 1644511149
transform 1 0 13800 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_144
timestamp 1644511149
transform 1 0 14352 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_148
timestamp 1644511149
transform 1 0 14720 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_213
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1644511149
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_239
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_246
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_252
timestamp 1644511149
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_260
timestamp 1644511149
transform 1 0 25024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_265
timestamp 1644511149
transform 1 0 25484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_290
timestamp 1644511149
transform 1 0 27784 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_294
timestamp 1644511149
transform 1 0 28152 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_301
timestamp 1644511149
transform 1 0 28796 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_316
timestamp 1644511149
transform 1 0 30176 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_19
timestamp 1644511149
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_117
timestamp 1644511149
transform 1 0 11868 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_147
timestamp 1644511149
transform 1 0 14628 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_168
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_181
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp 1644511149
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_226
timestamp 1644511149
transform 1 0 21896 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1644511149
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_264
timestamp 1644511149
transform 1 0 25392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_278
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1644511149
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_299
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_316
timestamp 1644511149
transform 1 0 30176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_151
timestamp 1644511149
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_187
timestamp 1644511149
transform 1 0 18308 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_204
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1644511149
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_230
timestamp 1644511149
transform 1 0 22264 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_250
timestamp 1644511149
transform 1 0 24104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_291
timestamp 1644511149
transform 1 0 27876 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_303
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_315
timestamp 1644511149
transform 1 0 30084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_319
timestamp 1644511149
transform 1 0 30452 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_7
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1644511149
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_149
timestamp 1644511149
transform 1 0 14812 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_158
timestamp 1644511149
transform 1 0 15640 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_166
timestamp 1644511149
transform 1 0 16376 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_174
timestamp 1644511149
transform 1 0 17112 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_186
timestamp 1644511149
transform 1 0 18216 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_201
timestamp 1644511149
transform 1 0 19596 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_230
timestamp 1644511149
transform 1 0 22264 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_262
timestamp 1644511149
transform 1 0 25208 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_274
timestamp 1644511149
transform 1 0 26312 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_282
timestamp 1644511149
transform 1 0 27048 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_316
timestamp 1644511149
transform 1 0 30176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_7
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_19
timestamp 1644511149
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_31
timestamp 1644511149
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_43
timestamp 1644511149
transform 1 0 5060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_121
timestamp 1644511149
transform 1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_132
timestamp 1644511149
transform 1 0 13248 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_138
timestamp 1644511149
transform 1 0 13800 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 1644511149
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_186
timestamp 1644511149
transform 1 0 18216 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_198
timestamp 1644511149
transform 1 0 19320 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1644511149
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_232
timestamp 1644511149
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_243
timestamp 1644511149
transform 1 0 23460 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_255
timestamp 1644511149
transform 1 0 24564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_267
timestamp 1644511149
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_292
timestamp 1644511149
transform 1 0 27968 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_304
timestamp 1644511149
transform 1 0 29072 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_316
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_14
timestamp 1644511149
transform 1 0 2392 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1644511149
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_125
timestamp 1644511149
transform 1 0 12604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_149
timestamp 1644511149
transform 1 0 14812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_157
timestamp 1644511149
transform 1 0 15548 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_179
timestamp 1644511149
transform 1 0 17572 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_205
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1644511149
transform 1 0 20700 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_222
timestamp 1644511149
transform 1 0 21528 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_234
timestamp 1644511149
transform 1 0 22632 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1644511149
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_274
timestamp 1644511149
transform 1 0 26312 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_284
timestamp 1644511149
transform 1 0 27232 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_294
timestamp 1644511149
transform 1 0 28152 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_316
timestamp 1644511149
transform 1 0 30176 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_7
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_14
timestamp 1644511149
transform 1 0 2392 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_26
timestamp 1644511149
transform 1 0 3496 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_38
timestamp 1644511149
transform 1 0 4600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1644511149
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_130
timestamp 1644511149
transform 1 0 13064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_134
timestamp 1644511149
transform 1 0 13432 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_143
timestamp 1644511149
transform 1 0 14260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_155
timestamp 1644511149
transform 1 0 15364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1644511149
transform 1 0 19044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_204
timestamp 1644511149
transform 1 0 19872 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_265
timestamp 1644511149
transform 1 0 25484 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_276
timestamp 1644511149
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_291
timestamp 1644511149
transform 1 0 27876 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_301
timestamp 1644511149
transform 1 0 28796 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_312
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_14
timestamp 1644511149
transform 1 0 2392 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1644511149
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_98
timestamp 1644511149
transform 1 0 10120 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_106
timestamp 1644511149
transform 1 0 10856 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_111
timestamp 1644511149
transform 1 0 11316 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_123
timestamp 1644511149
transform 1 0 12420 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1644511149
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_161
timestamp 1644511149
transform 1 0 15916 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_185
timestamp 1644511149
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_201
timestamp 1644511149
transform 1 0 19596 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_208
timestamp 1644511149
transform 1 0 20240 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_220
timestamp 1644511149
transform 1 0 21344 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_232
timestamp 1644511149
transform 1 0 22448 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_259
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_294
timestamp 1644511149
transform 1 0 28152 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_316
timestamp 1644511149
transform 1 0 30176 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_9
timestamp 1644511149
transform 1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_13
timestamp 1644511149
transform 1 0 2300 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_19
timestamp 1644511149
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_43
timestamp 1644511149
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_98
timestamp 1644511149
transform 1 0 10120 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1644511149
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_129
timestamp 1644511149
transform 1 0 12972 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_134
timestamp 1644511149
transform 1 0 13432 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_148
timestamp 1644511149
transform 1 0 14720 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_178
timestamp 1644511149
transform 1 0 17480 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_184
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_201
timestamp 1644511149
transform 1 0 19596 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_213
timestamp 1644511149
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1644511149
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_229
timestamp 1644511149
transform 1 0 22172 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1644511149
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_245
timestamp 1644511149
transform 1 0 23644 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_255
timestamp 1644511149
transform 1 0 24564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_265
timestamp 1644511149
transform 1 0 25484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_291
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_298
timestamp 1644511149
transform 1 0 28520 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_302
timestamp 1644511149
transform 1 0 28888 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_313
timestamp 1644511149
transform 1 0 29900 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_319
timestamp 1644511149
transform 1 0 30452 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_9
timestamp 1644511149
transform 1 0 1932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_13
timestamp 1644511149
transform 1 0 2300 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_94
timestamp 1644511149
transform 1 0 9752 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_122
timestamp 1644511149
transform 1 0 12328 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_130
timestamp 1644511149
transform 1 0 13064 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_135
timestamp 1644511149
transform 1 0 13524 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1644511149
transform 1 0 14352 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_156
timestamp 1644511149
transform 1 0 15456 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_162
timestamp 1644511149
transform 1 0 16008 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_167
timestamp 1644511149
transform 1 0 16468 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_179
timestamp 1644511149
transform 1 0 17572 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1644511149
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_205
timestamp 1644511149
transform 1 0 19964 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_228
timestamp 1644511149
transform 1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_259
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_275
timestamp 1644511149
transform 1 0 26404 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_288
timestamp 1644511149
transform 1 0 27600 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_316
timestamp 1644511149
transform 1 0 30176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_6
timestamp 1644511149
transform 1 0 1656 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_18
timestamp 1644511149
transform 1 0 2760 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_30
timestamp 1644511149
transform 1 0 3864 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_42
timestamp 1644511149
transform 1 0 4968 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1644511149
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_89
timestamp 1644511149
transform 1 0 9292 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_97
timestamp 1644511149
transform 1 0 10028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_109
timestamp 1644511149
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_157
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_178
timestamp 1644511149
transform 1 0 17480 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_186
timestamp 1644511149
transform 1 0 18216 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_197
timestamp 1644511149
transform 1 0 19228 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_233
timestamp 1644511149
transform 1 0 22540 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_247
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_259
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_265
timestamp 1644511149
transform 1 0 25484 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_289
timestamp 1644511149
transform 1 0 27692 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_296
timestamp 1644511149
transform 1 0 28336 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_312
timestamp 1644511149
transform 1 0 29808 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_6
timestamp 1644511149
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_18
timestamp 1644511149
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1644511149
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1644511149
transform 1 0 9476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_112
timestamp 1644511149
transform 1 0 11408 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_158
timestamp 1644511149
transform 1 0 15640 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_166
timestamp 1644511149
transform 1 0 16376 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_179
timestamp 1644511149
transform 1 0 17572 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1644511149
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_206
timestamp 1644511149
transform 1 0 20056 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_215
timestamp 1644511149
transform 1 0 20884 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_226
timestamp 1644511149
transform 1 0 21896 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_236
timestamp 1644511149
transform 1 0 22816 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_268
timestamp 1644511149
transform 1 0 25760 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_280
timestamp 1644511149
transform 1 0 26864 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_292
timestamp 1644511149
transform 1 0 27968 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_316
timestamp 1644511149
transform 1 0 30176 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_6
timestamp 1644511149
transform 1 0 1656 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_18
timestamp 1644511149
transform 1 0 2760 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1644511149
transform 1 0 3864 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1644511149
transform 1 0 4968 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1644511149
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_89
timestamp 1644511149
transform 1 0 9292 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_95
timestamp 1644511149
transform 1 0 9844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1644511149
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_117
timestamp 1644511149
transform 1 0 11868 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_123
timestamp 1644511149
transform 1 0 12420 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_133
timestamp 1644511149
transform 1 0 13340 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_146
timestamp 1644511149
transform 1 0 14536 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1644511149
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_173
timestamp 1644511149
transform 1 0 17020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_185
timestamp 1644511149
transform 1 0 18124 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_206
timestamp 1644511149
transform 1 0 20056 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_213
timestamp 1644511149
transform 1 0 20700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1644511149
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_255
timestamp 1644511149
transform 1 0 24564 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_263
timestamp 1644511149
transform 1 0 25300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_274
timestamp 1644511149
transform 1 0 26312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_301
timestamp 1644511149
transform 1 0 28796 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_308
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_316
timestamp 1644511149
transform 1 0 30176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1644511149
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_26
timestamp 1644511149
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_110
timestamp 1644511149
transform 1 0 11224 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_118
timestamp 1644511149
transform 1 0 11960 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_129
timestamp 1644511149
transform 1 0 12972 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_145
timestamp 1644511149
transform 1 0 14444 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_174
timestamp 1644511149
transform 1 0 17112 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_187
timestamp 1644511149
transform 1 0 18308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_201
timestamp 1644511149
transform 1 0 19596 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_208
timestamp 1644511149
transform 1 0 20240 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_220
timestamp 1644511149
transform 1 0 21344 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_232
timestamp 1644511149
transform 1 0 22448 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_244
timestamp 1644511149
transform 1 0 23552 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_262
timestamp 1644511149
transform 1 0 25208 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_275
timestamp 1644511149
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_287
timestamp 1644511149
transform 1 0 27508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_291
timestamp 1644511149
transform 1 0 27876 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_296
timestamp 1644511149
transform 1 0 28336 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_316
timestamp 1644511149
transform 1 0 30176 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_6
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_18
timestamp 1644511149
transform 1 0 2760 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1644511149
transform 1 0 3864 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_42
timestamp 1644511149
transform 1 0 4968 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1644511149
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_96
timestamp 1644511149
transform 1 0 9936 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_104
timestamp 1644511149
transform 1 0 10672 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_117
timestamp 1644511149
transform 1 0 11868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_133
timestamp 1644511149
transform 1 0 13340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_144
timestamp 1644511149
transform 1 0 14352 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_151
timestamp 1644511149
transform 1 0 14996 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_159
timestamp 1644511149
transform 1 0 15732 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_179
timestamp 1644511149
transform 1 0 17572 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_183
timestamp 1644511149
transform 1 0 17940 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_188
timestamp 1644511149
transform 1 0 18400 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_192
timestamp 1644511149
transform 1 0 18768 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_197
timestamp 1644511149
transform 1 0 19228 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_204
timestamp 1644511149
transform 1 0 19872 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_211
timestamp 1644511149
transform 1 0 20516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_288
timestamp 1644511149
transform 1 0 27600 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_296
timestamp 1644511149
transform 1 0 28336 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_304
timestamp 1644511149
transform 1 0 29072 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_316
timestamp 1644511149
transform 1 0 30176 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_6
timestamp 1644511149
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_18
timestamp 1644511149
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1644511149
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_103
timestamp 1644511149
transform 1 0 10580 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_107
timestamp 1644511149
transform 1 0 10948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_116
timestamp 1644511149
transform 1 0 11776 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_123
timestamp 1644511149
transform 1 0 12420 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_131
timestamp 1644511149
transform 1 0 13156 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_135
timestamp 1644511149
transform 1 0 13524 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_149
timestamp 1644511149
transform 1 0 14812 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_157
timestamp 1644511149
transform 1 0 15548 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_163
timestamp 1644511149
transform 1 0 16100 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_176
timestamp 1644511149
transform 1 0 17296 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_182
timestamp 1644511149
transform 1 0 17848 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_215
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_223
timestamp 1644511149
transform 1 0 21620 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_230
timestamp 1644511149
transform 1 0 22264 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_242
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_257
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_297
timestamp 1644511149
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1644511149
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_316
timestamp 1644511149
transform 1 0 30176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1644511149
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1644511149
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1644511149
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1644511149
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1644511149
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_89
timestamp 1644511149
transform 1 0 9292 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_101
timestamp 1644511149
transform 1 0 10396 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 1644511149
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_200
timestamp 1644511149
transform 1 0 19504 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_204
timestamp 1644511149
transform 1 0 19872 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_208
timestamp 1644511149
transform 1 0 20240 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1644511149
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_247
timestamp 1644511149
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_264
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_285
timestamp 1644511149
transform 1 0 27324 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_297
timestamp 1644511149
transform 1 0 28428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_319
timestamp 1644511149
transform 1 0 30452 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_6
timestamp 1644511149
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_18
timestamp 1644511149
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1644511149
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1644511149
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_110
timestamp 1644511149
transform 1 0 11224 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_122
timestamp 1644511149
transform 1 0 12328 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_134
timestamp 1644511149
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_149
timestamp 1644511149
transform 1 0 14812 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1644511149
transform 1 0 15272 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_166
timestamp 1644511149
transform 1 0 16376 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_200
timestamp 1644511149
transform 1 0 19504 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_204
timestamp 1644511149
transform 1 0 19872 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1644511149
transform 1 0 20424 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_223
timestamp 1644511149
transform 1 0 21620 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_232
timestamp 1644511149
transform 1 0 22448 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_240
timestamp 1644511149
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_263
timestamp 1644511149
transform 1 0 25300 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_274
timestamp 1644511149
transform 1 0 26312 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_282
timestamp 1644511149
transform 1 0 27048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_303
timestamp 1644511149
transform 1 0 28980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_315
timestamp 1644511149
transform 1 0 30084 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_319
timestamp 1644511149
transform 1 0 30452 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_6
timestamp 1644511149
transform 1 0 1656 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_18
timestamp 1644511149
transform 1 0 2760 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1644511149
transform 1 0 3864 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1644511149
transform 1 0 4968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1644511149
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_75
timestamp 1644511149
transform 1 0 8004 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_90
timestamp 1644511149
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1644511149
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1644511149
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_133
timestamp 1644511149
transform 1 0 13340 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_144
timestamp 1644511149
transform 1 0 14352 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_150
timestamp 1644511149
transform 1 0 14904 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_159
timestamp 1644511149
transform 1 0 15732 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_186
timestamp 1644511149
transform 1 0 18216 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_233
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_257
timestamp 1644511149
transform 1 0 24748 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_265
timestamp 1644511149
transform 1 0 25484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_285
timestamp 1644511149
transform 1 0 27324 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_292
timestamp 1644511149
transform 1 0 27968 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_304
timestamp 1644511149
transform 1 0 29072 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_316
timestamp 1644511149
transform 1 0 30176 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_49
timestamp 1644511149
transform 1 0 5612 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_61
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_73
timestamp 1644511149
transform 1 0 7820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_93
timestamp 1644511149
transform 1 0 9660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1644511149
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_119
timestamp 1644511149
transform 1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_131
timestamp 1644511149
transform 1 0 13156 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_149
timestamp 1644511149
transform 1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_185
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_214
timestamp 1644511149
transform 1 0 20792 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_227
timestamp 1644511149
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_235
timestamp 1644511149
transform 1 0 22724 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1644511149
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_260
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_272
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_282
timestamp 1644511149
transform 1 0 27048 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_292
timestamp 1644511149
transform 1 0 27968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1644511149
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_319
timestamp 1644511149
transform 1 0 30452 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_6
timestamp 1644511149
transform 1 0 1656 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_18
timestamp 1644511149
transform 1 0 2760 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_30
timestamp 1644511149
transform 1 0 3864 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_42
timestamp 1644511149
transform 1 0 4968 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1644511149
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_75
timestamp 1644511149
transform 1 0 8004 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_79
timestamp 1644511149
transform 1 0 8372 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_83
timestamp 1644511149
transform 1 0 8740 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_89
timestamp 1644511149
transform 1 0 9292 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_98
timestamp 1644511149
transform 1 0 10120 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_104
timestamp 1644511149
transform 1 0 10672 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_108
timestamp 1644511149
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_131
timestamp 1644511149
transform 1 0 13156 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_139
timestamp 1644511149
transform 1 0 13892 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_160
timestamp 1644511149
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_177
timestamp 1644511149
transform 1 0 17388 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_208
timestamp 1644511149
transform 1 0 20240 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_247
timestamp 1644511149
transform 1 0 23828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_253
timestamp 1644511149
transform 1 0 24380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_274
timestamp 1644511149
transform 1 0 26312 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_290
timestamp 1644511149
transform 1 0 27784 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_294
timestamp 1644511149
transform 1 0 28152 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_315
timestamp 1644511149
transform 1 0 30084 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_319
timestamp 1644511149
transform 1 0 30452 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_6
timestamp 1644511149
transform 1 0 1656 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_18
timestamp 1644511149
transform 1 0 2760 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1644511149
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_110
timestamp 1644511149
transform 1 0 11224 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_126
timestamp 1644511149
transform 1 0 12696 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1644511149
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_158
timestamp 1644511149
transform 1 0 15640 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_170
timestamp 1644511149
transform 1 0 16744 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_186
timestamp 1644511149
transform 1 0 18216 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1644511149
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_200
timestamp 1644511149
transform 1 0 19504 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_208
timestamp 1644511149
transform 1 0 20240 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_212
timestamp 1644511149
transform 1 0 20608 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_219
timestamp 1644511149
transform 1 0 21252 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_231
timestamp 1644511149
transform 1 0 22356 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_239
timestamp 1644511149
transform 1 0 23092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1644511149
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_263
timestamp 1644511149
transform 1 0 25300 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_297
timestamp 1644511149
transform 1 0 28428 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_305
timestamp 1644511149
transform 1 0 29164 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_316
timestamp 1644511149
transform 1 0 30176 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_6
timestamp 1644511149
transform 1 0 1656 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_18
timestamp 1644511149
transform 1 0 2760 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_30
timestamp 1644511149
transform 1 0 3864 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_42
timestamp 1644511149
transform 1 0 4968 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1644511149
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_77
timestamp 1644511149
transform 1 0 8188 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_84
timestamp 1644511149
transform 1 0 8832 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_96
timestamp 1644511149
transform 1 0 9936 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_108
timestamp 1644511149
transform 1 0 11040 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_121
timestamp 1644511149
transform 1 0 12236 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_135
timestamp 1644511149
transform 1 0 13524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_158
timestamp 1644511149
transform 1 0 15640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1644511149
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_178
timestamp 1644511149
transform 1 0 17480 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_186
timestamp 1644511149
transform 1 0 18216 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_201
timestamp 1644511149
transform 1 0 19596 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_207
timestamp 1644511149
transform 1 0 20148 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_229
timestamp 1644511149
transform 1 0 22172 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_234
timestamp 1644511149
transform 1 0 22632 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_248
timestamp 1644511149
transform 1 0 23920 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_254
timestamp 1644511149
transform 1 0 24472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_262
timestamp 1644511149
transform 1 0 25208 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_274
timestamp 1644511149
transform 1 0 26312 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_285
timestamp 1644511149
transform 1 0 27324 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_300
timestamp 1644511149
transform 1 0 28704 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_308
timestamp 1644511149
transform 1 0 29440 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_316
timestamp 1644511149
transform 1 0 30176 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_6
timestamp 1644511149
transform 1 0 1656 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_18
timestamp 1644511149
transform 1 0 2760 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_26
timestamp 1644511149
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_110
timestamp 1644511149
transform 1 0 11224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_131
timestamp 1644511149
transform 1 0 13156 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_145
timestamp 1644511149
transform 1 0 14444 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_155
timestamp 1644511149
transform 1 0 15364 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_172
timestamp 1644511149
transform 1 0 16928 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1644511149
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_205
timestamp 1644511149
transform 1 0 19964 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_213
timestamp 1644511149
transform 1 0 20700 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_231
timestamp 1644511149
transform 1 0 22356 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_244
timestamp 1644511149
transform 1 0 23552 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_260
timestamp 1644511149
transform 1 0 25024 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_272
timestamp 1644511149
transform 1 0 26128 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_278
timestamp 1644511149
transform 1 0 26680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_283
timestamp 1644511149
transform 1 0 27140 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_291
timestamp 1644511149
transform 1 0 27876 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_296
timestamp 1644511149
transform 1 0 28336 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_304
timestamp 1644511149
transform 1 0 29072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_316
timestamp 1644511149
transform 1 0 30176 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_6
timestamp 1644511149
transform 1 0 1656 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_18
timestamp 1644511149
transform 1 0 2760 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_30
timestamp 1644511149
transform 1 0 3864 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_42
timestamp 1644511149
transform 1 0 4968 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 1644511149
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_77
timestamp 1644511149
transform 1 0 8188 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_83
timestamp 1644511149
transform 1 0 8740 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_91
timestamp 1644511149
transform 1 0 9476 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_100
timestamp 1644511149
transform 1 0 10304 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_121
timestamp 1644511149
transform 1 0 12236 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_133
timestamp 1644511149
transform 1 0 13340 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_145
timestamp 1644511149
transform 1 0 14444 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_157
timestamp 1644511149
transform 1 0 15548 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1644511149
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_208
timestamp 1644511149
transform 1 0 20240 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1644511149
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_236
timestamp 1644511149
transform 1 0 22816 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_246
timestamp 1644511149
transform 1 0 23736 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_255
timestamp 1644511149
transform 1 0 24564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_267
timestamp 1644511149
transform 1 0 25668 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_271
timestamp 1644511149
transform 1 0 26036 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_276
timestamp 1644511149
transform 1 0 26496 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_290
timestamp 1644511149
transform 1 0 27784 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_304
timestamp 1644511149
transform 1 0 29072 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_316
timestamp 1644511149
transform 1 0 30176 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_73
timestamp 1644511149
transform 1 0 7820 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_80
timestamp 1644511149
transform 1 0 8464 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1644511149
transform 1 0 9476 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_100
timestamp 1644511149
transform 1 0 10304 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_112
timestamp 1644511149
transform 1 0 11408 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_124
timestamp 1644511149
transform 1 0 12512 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_136
timestamp 1644511149
transform 1 0 13616 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_162
timestamp 1644511149
transform 1 0 16008 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_169
timestamp 1644511149
transform 1 0 16652 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_176
timestamp 1644511149
transform 1 0 17296 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_183
timestamp 1644511149
transform 1 0 17940 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_187
timestamp 1644511149
transform 1 0 18308 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1644511149
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_200
timestamp 1644511149
transform 1 0 19504 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_226
timestamp 1644511149
transform 1 0 21896 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_234
timestamp 1644511149
transform 1 0 22632 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1644511149
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_274
timestamp 1644511149
transform 1 0 26312 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_288
timestamp 1644511149
transform 1 0 27600 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_302
timestamp 1644511149
transform 1 0 28888 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_316
timestamp 1644511149
transform 1 0 30176 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_6
timestamp 1644511149
transform 1 0 1656 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_18
timestamp 1644511149
transform 1 0 2760 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1644511149
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1644511149
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1644511149
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_156
timestamp 1644511149
transform 1 0 15456 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1644511149
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_172
timestamp 1644511149
transform 1 0 16928 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_184
timestamp 1644511149
transform 1 0 18032 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_191
timestamp 1644511149
transform 1 0 18676 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_199
timestamp 1644511149
transform 1 0 19412 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_212
timestamp 1644511149
transform 1 0 20608 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1644511149
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_235
timestamp 1644511149
transform 1 0 22724 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_242
timestamp 1644511149
transform 1 0 23368 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_254
timestamp 1644511149
transform 1 0 24472 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_260
timestamp 1644511149
transform 1 0 25024 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_264
timestamp 1644511149
transform 1 0 25392 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_274
timestamp 1644511149
transform 1 0 26312 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_291
timestamp 1644511149
transform 1 0 27876 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_303
timestamp 1644511149
transform 1 0 28980 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_307
timestamp 1644511149
transform 1 0 29348 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_316
timestamp 1644511149
transform 1 0 30176 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_6
timestamp 1644511149
transform 1 0 1656 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_18
timestamp 1644511149
transform 1 0 2760 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1644511149
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_90
timestamp 1644511149
transform 1 0 9384 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_98
timestamp 1644511149
transform 1 0 10120 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_111
timestamp 1644511149
transform 1 0 11316 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_135
timestamp 1644511149
transform 1 0 13524 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_144
timestamp 1644511149
transform 1 0 14352 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_169
timestamp 1644511149
transform 1 0 16652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_174
timestamp 1644511149
transform 1 0 17112 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_182
timestamp 1644511149
transform 1 0 17848 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_190
timestamp 1644511149
transform 1 0 18584 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_207
timestamp 1644511149
transform 1 0 20148 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_211
timestamp 1644511149
transform 1 0 20516 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_215
timestamp 1644511149
transform 1 0 20884 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_223
timestamp 1644511149
transform 1 0 21620 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_240
timestamp 1644511149
transform 1 0 23184 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_247
timestamp 1644511149
transform 1 0 23828 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_258
timestamp 1644511149
transform 1 0 24840 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_269
timestamp 1644511149
transform 1 0 25852 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_282
timestamp 1644511149
transform 1 0 27048 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_292
timestamp 1644511149
transform 1 0 27968 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1644511149
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_315
timestamp 1644511149
transform 1 0 30084 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_319
timestamp 1644511149
transform 1 0 30452 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_6
timestamp 1644511149
transform 1 0 1656 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_18
timestamp 1644511149
transform 1 0 2760 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_30
timestamp 1644511149
transform 1 0 3864 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_42
timestamp 1644511149
transform 1 0 4968 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_54
timestamp 1644511149
transform 1 0 6072 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_77
timestamp 1644511149
transform 1 0 8188 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_84
timestamp 1644511149
transform 1 0 8832 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_92
timestamp 1644511149
transform 1 0 9568 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_101
timestamp 1644511149
transform 1 0 10396 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_109
timestamp 1644511149
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_117
timestamp 1644511149
transform 1 0 11868 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_121
timestamp 1644511149
transform 1 0 12236 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_129
timestamp 1644511149
transform 1 0 12972 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_136
timestamp 1644511149
transform 1 0 13616 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_157
timestamp 1644511149
transform 1 0 15548 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1644511149
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_173
timestamp 1644511149
transform 1 0 17020 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_200
timestamp 1644511149
transform 1 0 19504 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_207
timestamp 1644511149
transform 1 0 20148 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_214
timestamp 1644511149
transform 1 0 20792 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1644511149
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_245
timestamp 1644511149
transform 1 0 23644 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_269
timestamp 1644511149
transform 1 0 25852 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_274
timestamp 1644511149
transform 1 0 26312 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_286
timestamp 1644511149
transform 1 0 27416 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_304
timestamp 1644511149
transform 1 0 29072 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_316
timestamp 1644511149
transform 1 0 30176 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_6
timestamp 1644511149
transform 1 0 1656 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_13
timestamp 1644511149
transform 1 0 2300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_25
timestamp 1644511149
transform 1 0 3404 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_94
timestamp 1644511149
transform 1 0 9752 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_117
timestamp 1644511149
transform 1 0 11868 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_125
timestamp 1644511149
transform 1 0 12604 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_151
timestamp 1644511149
transform 1 0 14996 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_163
timestamp 1644511149
transform 1 0 16100 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_171
timestamp 1644511149
transform 1 0 16836 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1644511149
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_201
timestamp 1644511149
transform 1 0 19596 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_207
timestamp 1644511149
transform 1 0 20148 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_228
timestamp 1644511149
transform 1 0 22080 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_235
timestamp 1644511149
transform 1 0 22724 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_247
timestamp 1644511149
transform 1 0 23828 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_261
timestamp 1644511149
transform 1 0 25116 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_267
timestamp 1644511149
transform 1 0 25668 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_272
timestamp 1644511149
transform 1 0 26128 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_280
timestamp 1644511149
transform 1 0 26864 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_284
timestamp 1644511149
transform 1 0 27232 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_297
timestamp 1644511149
transform 1 0 28428 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_304
timestamp 1644511149
transform 1 0 29072 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_315
timestamp 1644511149
transform 1 0 30084 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_319
timestamp 1644511149
transform 1 0 30452 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_10
timestamp 1644511149
transform 1 0 2024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_17
timestamp 1644511149
transform 1 0 2668 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_29
timestamp 1644511149
transform 1 0 3772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_41
timestamp 1644511149
transform 1 0 4876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1644511149
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_89
timestamp 1644511149
transform 1 0 9292 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_100
timestamp 1644511149
transform 1 0 10304 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_123
timestamp 1644511149
transform 1 0 12420 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_146
timestamp 1644511149
transform 1 0 14536 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_154
timestamp 1644511149
transform 1 0 15272 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_162
timestamp 1644511149
transform 1 0 16008 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_199
timestamp 1644511149
transform 1 0 19412 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_220
timestamp 1644511149
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_233
timestamp 1644511149
transform 1 0 22540 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_239
timestamp 1644511149
transform 1 0 23092 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_248
timestamp 1644511149
transform 1 0 23920 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_262
timestamp 1644511149
transform 1 0 25208 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_75_274
timestamp 1644511149
transform 1 0 26312 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_289
timestamp 1644511149
transform 1 0 27692 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_300
timestamp 1644511149
transform 1 0 28704 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_308
timestamp 1644511149
transform 1 0 29440 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_316
timestamp 1644511149
transform 1 0 30176 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_10
timestamp 1644511149
transform 1 0 2024 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_19
timestamp 1644511149
transform 1 0 2852 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_101
timestamp 1644511149
transform 1 0 10396 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_114
timestamp 1644511149
transform 1 0 11592 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_120
timestamp 1644511149
transform 1 0 12144 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_129
timestamp 1644511149
transform 1 0 12972 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_136
timestamp 1644511149
transform 1 0 13616 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_150
timestamp 1644511149
transform 1 0 14904 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_163
timestamp 1644511149
transform 1 0 16100 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_167
timestamp 1644511149
transform 1 0 16468 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_188
timestamp 1644511149
transform 1 0 18400 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_206
timestamp 1644511149
transform 1 0 20056 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_219
timestamp 1644511149
transform 1 0 21252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_228
timestamp 1644511149
transform 1 0 22080 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_235
timestamp 1644511149
transform 1 0 22724 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_248
timestamp 1644511149
transform 1 0 23920 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_261
timestamp 1644511149
transform 1 0 25116 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_273
timestamp 1644511149
transform 1 0 26220 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_279
timestamp 1644511149
transform 1 0 26772 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_286
timestamp 1644511149
transform 1 0 27416 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_76_302
timestamp 1644511149
transform 1 0 28888 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_316
timestamp 1644511149
transform 1 0 30176 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_10
timestamp 1644511149
transform 1 0 2024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_17
timestamp 1644511149
transform 1 0 2668 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_29
timestamp 1644511149
transform 1 0 3772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_41
timestamp 1644511149
transform 1 0 4876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1644511149
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_101
timestamp 1644511149
transform 1 0 10396 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_108
timestamp 1644511149
transform 1 0 11040 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_124
timestamp 1644511149
transform 1 0 12512 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_132
timestamp 1644511149
transform 1 0 13248 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_138
timestamp 1644511149
transform 1 0 13800 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_143
timestamp 1644511149
transform 1 0 14260 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_151
timestamp 1644511149
transform 1 0 14996 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_164
timestamp 1644511149
transform 1 0 16192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_178
timestamp 1644511149
transform 1 0 17480 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_190
timestamp 1644511149
transform 1 0 18584 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_198
timestamp 1644511149
transform 1 0 19320 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_220
timestamp 1644511149
transform 1 0 21344 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_229
timestamp 1644511149
transform 1 0 22172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_233
timestamp 1644511149
transform 1 0 22540 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_238
timestamp 1644511149
transform 1 0 23000 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_242
timestamp 1644511149
transform 1 0 23368 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_248
timestamp 1644511149
transform 1 0 23920 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_256
timestamp 1644511149
transform 1 0 24656 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1644511149
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_276
timestamp 1644511149
transform 1 0 26496 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_287
timestamp 1644511149
transform 1 0 27508 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_294
timestamp 1644511149
transform 1 0 28152 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_302
timestamp 1644511149
transform 1 0 28888 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_308
timestamp 1644511149
transform 1 0 29440 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_316
timestamp 1644511149
transform 1 0 30176 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_10
timestamp 1644511149
transform 1 0 2024 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_22
timestamp 1644511149
transform 1 0 3128 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_114
timestamp 1644511149
transform 1 0 11592 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_126
timestamp 1644511149
transform 1 0 12696 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_136
timestamp 1644511149
transform 1 0 13616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_171
timestamp 1644511149
transform 1 0 16836 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_192
timestamp 1644511149
transform 1 0 18768 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_206
timestamp 1644511149
transform 1 0 20056 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_219
timestamp 1644511149
transform 1 0 21252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_225
timestamp 1644511149
transform 1 0 21804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_242
timestamp 1644511149
transform 1 0 23368 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1644511149
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_257
timestamp 1644511149
transform 1 0 24748 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_266
timestamp 1644511149
transform 1 0 25576 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_278
timestamp 1644511149
transform 1 0 26680 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_282
timestamp 1644511149
transform 1 0 27048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_287
timestamp 1644511149
transform 1 0 27508 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_296
timestamp 1644511149
transform 1 0 28336 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_304
timestamp 1644511149
transform 1 0 29072 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_315
timestamp 1644511149
transform 1 0 30084 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_319
timestamp 1644511149
transform 1 0 30452 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_6
timestamp 1644511149
transform 1 0 1656 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_12
timestamp 1644511149
transform 1 0 2208 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_18
timestamp 1644511149
transform 1 0 2760 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1644511149
transform 1 0 3864 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1644511149
transform 1 0 4968 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_54
timestamp 1644511149
transform 1 0 6072 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_121
timestamp 1644511149
transform 1 0 12236 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_132
timestamp 1644511149
transform 1 0 13248 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_136
timestamp 1644511149
transform 1 0 13616 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_157
timestamp 1644511149
transform 1 0 15548 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1644511149
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_200
timestamp 1644511149
transform 1 0 19504 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_213
timestamp 1644511149
transform 1 0 20700 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 1644511149
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_229
timestamp 1644511149
transform 1 0 22172 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_241
timestamp 1644511149
transform 1 0 23276 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_255
timestamp 1644511149
transform 1 0 24564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_267
timestamp 1644511149
transform 1 0 25668 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_301
timestamp 1644511149
transform 1 0 28796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_311
timestamp 1644511149
transform 1 0 29716 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_319
timestamp 1644511149
transform 1 0 30452 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_6
timestamp 1644511149
transform 1 0 1656 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_12
timestamp 1644511149
transform 1 0 2208 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_18
timestamp 1644511149
transform 1 0 2760 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_26
timestamp 1644511149
transform 1 0 3496 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_103
timestamp 1644511149
transform 1 0 10580 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_111
timestamp 1644511149
transform 1 0 11316 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_122
timestamp 1644511149
transform 1 0 12328 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_134
timestamp 1644511149
transform 1 0 13432 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_148
timestamp 1644511149
transform 1 0 14720 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_155
timestamp 1644511149
transform 1 0 15364 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_179
timestamp 1644511149
transform 1 0 17572 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_187
timestamp 1644511149
transform 1 0 18308 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_207
timestamp 1644511149
transform 1 0 20148 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_231
timestamp 1644511149
transform 1 0 22356 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_242
timestamp 1644511149
transform 1 0 23368 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1644511149
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_261
timestamp 1644511149
transform 1 0 25116 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_275
timestamp 1644511149
transform 1 0 26404 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_287
timestamp 1644511149
transform 1 0 27508 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_299
timestamp 1644511149
transform 1 0 28612 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_315
timestamp 1644511149
transform 1 0 30084 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_319
timestamp 1644511149
transform 1 0 30452 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_6
timestamp 1644511149
transform 1 0 1656 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_18
timestamp 1644511149
transform 1 0 2760 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1644511149
transform 1 0 3864 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1644511149
transform 1 0 4968 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1644511149
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_150
timestamp 1644511149
transform 1 0 14904 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_154
timestamp 1644511149
transform 1 0 15272 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_164
timestamp 1644511149
transform 1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_178
timestamp 1644511149
transform 1 0 17480 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_186
timestamp 1644511149
transform 1 0 18216 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_192
timestamp 1644511149
transform 1 0 18768 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_196
timestamp 1644511149
transform 1 0 19136 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1644511149
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_231
timestamp 1644511149
transform 1 0 22356 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_239
timestamp 1644511149
transform 1 0 23092 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_244
timestamp 1644511149
transform 1 0 23552 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_256
timestamp 1644511149
transform 1 0 24656 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_270
timestamp 1644511149
transform 1 0 25944 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1644511149
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_301
timestamp 1644511149
transform 1 0 28796 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_306
timestamp 1644511149
transform 1 0 29256 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_316
timestamp 1644511149
transform 1 0 30176 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_6
timestamp 1644511149
transform 1 0 1656 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_17
timestamp 1644511149
transform 1 0 2668 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_25
timestamp 1644511149
transform 1 0 3404 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1644511149
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_129
timestamp 1644511149
transform 1 0 12972 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1644511149
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_164
timestamp 1644511149
transform 1 0 16192 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_172
timestamp 1644511149
transform 1 0 16928 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_192
timestamp 1644511149
transform 1 0 18768 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_200
timestamp 1644511149
transform 1 0 19504 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_207
timestamp 1644511149
transform 1 0 20148 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_215
timestamp 1644511149
transform 1 0 20884 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_227
timestamp 1644511149
transform 1 0 21988 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_233
timestamp 1644511149
transform 1 0 22540 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_244
timestamp 1644511149
transform 1 0 23552 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_261
timestamp 1644511149
transform 1 0 25116 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_273
timestamp 1644511149
transform 1 0 26220 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_282
timestamp 1644511149
transform 1 0 27048 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_296
timestamp 1644511149
transform 1 0 28336 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_304
timestamp 1644511149
transform 1 0 29072 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_316
timestamp 1644511149
transform 1 0 30176 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_6
timestamp 1644511149
transform 1 0 1656 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_13
timestamp 1644511149
transform 1 0 2300 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_25
timestamp 1644511149
transform 1 0 3404 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_37
timestamp 1644511149
transform 1 0 4508 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_49
timestamp 1644511149
transform 1 0 5612 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1644511149
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1644511149
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1644511149
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_125
timestamp 1644511149
transform 1 0 12604 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_142
timestamp 1644511149
transform 1 0 14168 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_155
timestamp 1644511149
transform 1 0 15364 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_159
timestamp 1644511149
transform 1 0 15732 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_164
timestamp 1644511149
transform 1 0 16192 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_183
timestamp 1644511149
transform 1 0 17940 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_190
timestamp 1644511149
transform 1 0 18584 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_197
timestamp 1644511149
transform 1 0 19228 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_205
timestamp 1644511149
transform 1 0 19964 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_211
timestamp 1644511149
transform 1 0 20516 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1644511149
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_237
timestamp 1644511149
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_249
timestamp 1644511149
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_261
timestamp 1644511149
transform 1 0 25116 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_269
timestamp 1644511149
transform 1 0 25852 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1644511149
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_285
timestamp 1644511149
transform 1 0 27324 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_296
timestamp 1644511149
transform 1 0 28336 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_304
timestamp 1644511149
transform 1 0 29072 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_316
timestamp 1644511149
transform 1 0 30176 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_84_3
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_9
timestamp 1644511149
transform 1 0 1932 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 1644511149
transform 1 0 2760 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_26
timestamp 1644511149
transform 1 0 3496 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1644511149
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1644511149
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_97
timestamp 1644511149
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_109
timestamp 1644511149
transform 1 0 11132 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_115
timestamp 1644511149
transform 1 0 11684 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_125
timestamp 1644511149
transform 1 0 12604 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_131
timestamp 1644511149
transform 1 0 13156 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_136
timestamp 1644511149
transform 1 0 13616 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_151
timestamp 1644511149
transform 1 0 14996 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_159
timestamp 1644511149
transform 1 0 15732 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_166
timestamp 1644511149
transform 1 0 16376 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_191
timestamp 1644511149
transform 1 0 18676 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1644511149
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_200
timestamp 1644511149
transform 1 0 19504 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_208
timestamp 1644511149
transform 1 0 20240 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_213
timestamp 1644511149
transform 1 0 20700 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_221
timestamp 1644511149
transform 1 0 21436 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_228
timestamp 1644511149
transform 1 0 22080 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_240
timestamp 1644511149
transform 1 0 23184 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_253
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_265
timestamp 1644511149
transform 1 0 25484 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_275
timestamp 1644511149
transform 1 0 26404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_281
timestamp 1644511149
transform 1 0 26956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_288
timestamp 1644511149
transform 1 0 27600 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_296
timestamp 1644511149
transform 1 0 28336 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_304
timestamp 1644511149
transform 1 0 29072 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_315
timestamp 1644511149
transform 1 0 30084 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_319
timestamp 1644511149
transform 1 0 30452 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_10
timestamp 1644511149
transform 1 0 2024 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_19
timestamp 1644511149
transform 1 0 2852 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_26
timestamp 1644511149
transform 1 0 3496 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_38
timestamp 1644511149
transform 1 0 4600 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_50
timestamp 1644511149
transform 1 0 5704 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_93
timestamp 1644511149
transform 1 0 9660 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_85_102
timestamp 1644511149
transform 1 0 10488 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_110
timestamp 1644511149
transform 1 0 11224 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_122
timestamp 1644511149
transform 1 0 12328 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_134
timestamp 1644511149
transform 1 0 13432 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_142
timestamp 1644511149
transform 1 0 14168 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_149
timestamp 1644511149
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1644511149
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1644511149
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_169
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_173
timestamp 1644511149
transform 1 0 17020 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_182
timestamp 1644511149
transform 1 0 17848 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_194
timestamp 1644511149
transform 1 0 18952 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_198
timestamp 1644511149
transform 1 0 19320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_208
timestamp 1644511149
transform 1 0 20240 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_216
timestamp 1644511149
transform 1 0 20976 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_238
timestamp 1644511149
transform 1 0 23000 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_246
timestamp 1644511149
transform 1 0 23736 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_254
timestamp 1644511149
transform 1 0 24472 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_258
timestamp 1644511149
transform 1 0 24840 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_263
timestamp 1644511149
transform 1 0 25300 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_275
timestamp 1644511149
transform 1 0 26404 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1644511149
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_289
timestamp 1644511149
transform 1 0 27692 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_293
timestamp 1644511149
transform 1 0 28060 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_303
timestamp 1644511149
transform 1 0 28980 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_316
timestamp 1644511149
transform 1 0 30176 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_10
timestamp 1644511149
transform 1 0 2024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_19
timestamp 1644511149
transform 1 0 2852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1644511149
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1644511149
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_93
timestamp 1644511149
transform 1 0 9660 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_113
timestamp 1644511149
transform 1 0 11500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_126
timestamp 1644511149
transform 1 0 12696 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_134
timestamp 1644511149
transform 1 0 13432 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_86_144
timestamp 1644511149
transform 1 0 14352 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_156
timestamp 1644511149
transform 1 0 15456 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_168
timestamp 1644511149
transform 1 0 16560 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_180
timestamp 1644511149
transform 1 0 17664 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_192
timestamp 1644511149
transform 1 0 18768 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_209
timestamp 1644511149
transform 1 0 20332 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_217
timestamp 1644511149
transform 1 0 21068 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_86_231
timestamp 1644511149
transform 1 0 22356 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_237
timestamp 1644511149
transform 1 0 22908 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_242
timestamp 1644511149
transform 1 0 23368 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_250
timestamp 1644511149
transform 1 0 24104 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_253
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_261
timestamp 1644511149
transform 1 0 25116 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_86_272
timestamp 1644511149
transform 1 0 26128 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_284
timestamp 1644511149
transform 1 0 27232 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_294
timestamp 1644511149
transform 1 0 28152 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1644511149
transform 1 0 29072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_316
timestamp 1644511149
transform 1 0 30176 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_10
timestamp 1644511149
transform 1 0 2024 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_17
timestamp 1644511149
transform 1 0 2668 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_29
timestamp 1644511149
transform 1 0 3772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_41
timestamp 1644511149
transform 1 0 4876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1644511149
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1644511149
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1644511149
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_113
timestamp 1644511149
transform 1 0 11500 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_87_118
timestamp 1644511149
transform 1 0 11960 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_126
timestamp 1644511149
transform 1 0 12696 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_87_148
timestamp 1644511149
transform 1 0 14720 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_87_159
timestamp 1644511149
transform 1 0 15732 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1644511149
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_169
timestamp 1644511149
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_181
timestamp 1644511149
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_193
timestamp 1644511149
transform 1 0 18860 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_201
timestamp 1644511149
transform 1 0 19596 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_206
timestamp 1644511149
transform 1 0 20056 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_214
timestamp 1644511149
transform 1 0 20792 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_222
timestamp 1644511149
transform 1 0 21528 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_87_225
timestamp 1644511149
transform 1 0 21804 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_239
timestamp 1644511149
transform 1 0 23092 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_245
timestamp 1644511149
transform 1 0 23644 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_254
timestamp 1644511149
transform 1 0 24472 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_266
timestamp 1644511149
transform 1 0 25576 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_278
timestamp 1644511149
transform 1 0 26680 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1644511149
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_293
timestamp 1644511149
transform 1 0 28060 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_303
timestamp 1644511149
transform 1 0 28980 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_316
timestamp 1644511149
transform 1 0 30176 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_10
timestamp 1644511149
transform 1 0 2024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_19
timestamp 1644511149
transform 1 0 2852 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1644511149
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_97
timestamp 1644511149
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_109
timestamp 1644511149
transform 1 0 11132 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_115
timestamp 1644511149
transform 1 0 11684 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1644511149
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1644511149
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_141
timestamp 1644511149
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_153
timestamp 1644511149
transform 1 0 15180 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_173
timestamp 1644511149
transform 1 0 17020 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_185
timestamp 1644511149
transform 1 0 18124 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_193
timestamp 1644511149
transform 1 0 18860 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_197
timestamp 1644511149
transform 1 0 19228 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_201
timestamp 1644511149
transform 1 0 19596 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_205
timestamp 1644511149
transform 1 0 19964 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_225
timestamp 1644511149
transform 1 0 21804 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_237
timestamp 1644511149
transform 1 0 22908 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_248
timestamp 1644511149
transform 1 0 23920 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_260
timestamp 1644511149
transform 1 0 25024 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_272
timestamp 1644511149
transform 1 0 26128 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_284
timestamp 1644511149
transform 1 0 27232 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_88_296
timestamp 1644511149
transform 1 0 28336 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_304
timestamp 1644511149
transform 1 0 29072 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_309
timestamp 1644511149
transform 1 0 29532 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_316
timestamp 1644511149
transform 1 0 30176 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_6
timestamp 1644511149
transform 1 0 1656 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_18
timestamp 1644511149
transform 1 0 2760 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_30
timestamp 1644511149
transform 1 0 3864 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_42
timestamp 1644511149
transform 1 0 4968 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_54
timestamp 1644511149
transform 1 0 6072 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1644511149
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1644511149
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_113
timestamp 1644511149
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_125
timestamp 1644511149
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_137
timestamp 1644511149
transform 1 0 13708 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_145
timestamp 1644511149
transform 1 0 14444 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_155
timestamp 1644511149
transform 1 0 15364 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1644511149
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_169
timestamp 1644511149
transform 1 0 16652 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_175
timestamp 1644511149
transform 1 0 17204 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_180
timestamp 1644511149
transform 1 0 17664 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_192
timestamp 1644511149
transform 1 0 18768 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_204
timestamp 1644511149
transform 1 0 19872 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_209
timestamp 1644511149
transform 1 0 20332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_221
timestamp 1644511149
transform 1 0 21436 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_229
timestamp 1644511149
transform 1 0 22172 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_236
timestamp 1644511149
transform 1 0 22816 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_248
timestamp 1644511149
transform 1 0 23920 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_258
timestamp 1644511149
transform 1 0 24840 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_269
timestamp 1644511149
transform 1 0 25852 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_277
timestamp 1644511149
transform 1 0 26588 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_281
timestamp 1644511149
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_293
timestamp 1644511149
transform 1 0 28060 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_301
timestamp 1644511149
transform 1 0 28796 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_306
timestamp 1644511149
transform 1 0 29256 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_316
timestamp 1644511149
transform 1 0 30176 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_6
timestamp 1644511149
transform 1 0 1656 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_13
timestamp 1644511149
transform 1 0 2300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_25
timestamp 1644511149
transform 1 0 3404 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_97
timestamp 1644511149
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_109
timestamp 1644511149
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_121
timestamp 1644511149
transform 1 0 12236 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_90_130
timestamp 1644511149
transform 1 0 13064 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1644511149
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_141
timestamp 1644511149
transform 1 0 14076 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_153
timestamp 1644511149
transform 1 0 15180 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_160
timestamp 1644511149
transform 1 0 15824 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_172
timestamp 1644511149
transform 1 0 16928 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_180
timestamp 1644511149
transform 1 0 17664 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_184
timestamp 1644511149
transform 1 0 18032 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_192
timestamp 1644511149
transform 1 0 18768 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_206
timestamp 1644511149
transform 1 0 20056 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_219
timestamp 1644511149
transform 1 0 21252 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_90_227
timestamp 1644511149
transform 1 0 21988 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_237
timestamp 1644511149
transform 1 0 22908 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_249
timestamp 1644511149
transform 1 0 24012 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_90_260
timestamp 1644511149
transform 1 0 25024 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_273
timestamp 1644511149
transform 1 0 26220 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_285
timestamp 1644511149
transform 1 0 27324 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_297
timestamp 1644511149
transform 1 0 28428 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_304
timestamp 1644511149
transform 1 0 29072 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_309
timestamp 1644511149
transform 1 0 29532 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_316
timestamp 1644511149
transform 1 0 30176 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_91_3
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_9
timestamp 1644511149
transform 1 0 1932 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_21
timestamp 1644511149
transform 1 0 3036 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_33
timestamp 1644511149
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1644511149
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1644511149
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1644511149
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1644511149
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_116
timestamp 1644511149
transform 1 0 11776 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_124
timestamp 1644511149
transform 1 0 12512 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_144
timestamp 1644511149
transform 1 0 14352 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_164
timestamp 1644511149
transform 1 0 16192 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_169
timestamp 1644511149
transform 1 0 16652 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_176
timestamp 1644511149
transform 1 0 17296 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_189
timestamp 1644511149
transform 1 0 18492 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_213
timestamp 1644511149
transform 1 0 20700 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_221
timestamp 1644511149
transform 1 0 21436 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_91_234
timestamp 1644511149
transform 1 0 22632 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_240
timestamp 1644511149
transform 1 0 23184 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_251
timestamp 1644511149
transform 1 0 24196 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_263
timestamp 1644511149
transform 1 0 25300 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1644511149
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1644511149
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_281
timestamp 1644511149
transform 1 0 26956 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_290
timestamp 1644511149
transform 1 0 27784 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_303
timestamp 1644511149
transform 1 0 28980 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_316
timestamp 1644511149
transform 1 0 30176 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_6
timestamp 1644511149
transform 1 0 1656 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_13
timestamp 1644511149
transform 1 0 2300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_25
timestamp 1644511149
transform 1 0 3404 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1644511149
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1644511149
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1644511149
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1644511149
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1644511149
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_97
timestamp 1644511149
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_109
timestamp 1644511149
transform 1 0 11132 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_115
timestamp 1644511149
transform 1 0 11684 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_135
timestamp 1644511149
transform 1 0 13524 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1644511149
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_149
timestamp 1644511149
transform 1 0 14812 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_156
timestamp 1644511149
transform 1 0 15456 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_168
timestamp 1644511149
transform 1 0 16560 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_175
timestamp 1644511149
transform 1 0 17204 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_188
timestamp 1644511149
transform 1 0 18400 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_206
timestamp 1644511149
transform 1 0 20056 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_210
timestamp 1644511149
transform 1 0 20424 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_215
timestamp 1644511149
transform 1 0 20884 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_223
timestamp 1644511149
transform 1 0 21620 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_92_242
timestamp 1644511149
transform 1 0 23368 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_250
timestamp 1644511149
transform 1 0 24104 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_253
timestamp 1644511149
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_265
timestamp 1644511149
transform 1 0 25484 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_279
timestamp 1644511149
transform 1 0 26772 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_291
timestamp 1644511149
transform 1 0 27876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_304
timestamp 1644511149
transform 1 0 29072 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_309
timestamp 1644511149
transform 1 0 29532 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_316
timestamp 1644511149
transform 1 0 30176 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_3
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_9
timestamp 1644511149
transform 1 0 1932 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_21
timestamp 1644511149
transform 1 0 3036 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_33
timestamp 1644511149
transform 1 0 4140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_45
timestamp 1644511149
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1644511149
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_93
timestamp 1644511149
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1644511149
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1644511149
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_113
timestamp 1644511149
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_125
timestamp 1644511149
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_137
timestamp 1644511149
transform 1 0 13708 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_155
timestamp 1644511149
transform 1 0 15364 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1644511149
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_169
timestamp 1644511149
transform 1 0 16652 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_177
timestamp 1644511149
transform 1 0 17388 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_183
timestamp 1644511149
transform 1 0 17940 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_190
timestamp 1644511149
transform 1 0 18584 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_198
timestamp 1644511149
transform 1 0 19320 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_205
timestamp 1644511149
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_220
timestamp 1644511149
transform 1 0 21344 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_229
timestamp 1644511149
transform 1 0 22172 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_236
timestamp 1644511149
transform 1 0 22816 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_242
timestamp 1644511149
transform 1 0 23368 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_247
timestamp 1644511149
transform 1 0 23828 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_259
timestamp 1644511149
transform 1 0 24932 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_267
timestamp 1644511149
transform 1 0 25668 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_276
timestamp 1644511149
transform 1 0 26496 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_281
timestamp 1644511149
transform 1 0 26956 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_285
timestamp 1644511149
transform 1 0 27324 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_294
timestamp 1644511149
transform 1 0 28152 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_307
timestamp 1644511149
transform 1 0 29348 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_311
timestamp 1644511149
transform 1 0 29716 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_316
timestamp 1644511149
transform 1 0 30176 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_7
timestamp 1644511149
transform 1 0 1748 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_14
timestamp 1644511149
transform 1 0 2392 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1644511149
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1644511149
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1644511149
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1644511149
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_97
timestamp 1644511149
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_109
timestamp 1644511149
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_121
timestamp 1644511149
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1644511149
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1644511149
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_141
timestamp 1644511149
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_153
timestamp 1644511149
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_165
timestamp 1644511149
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_177
timestamp 1644511149
transform 1 0 17388 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_181
timestamp 1644511149
transform 1 0 17756 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_185
timestamp 1644511149
transform 1 0 18124 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_192
timestamp 1644511149
transform 1 0 18768 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_201
timestamp 1644511149
transform 1 0 19596 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_225
timestamp 1644511149
transform 1 0 21804 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_234
timestamp 1644511149
transform 1 0 22632 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_246
timestamp 1644511149
transform 1 0 23736 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_94_253
timestamp 1644511149
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_265
timestamp 1644511149
transform 1 0 25484 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_272
timestamp 1644511149
transform 1 0 26128 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_282
timestamp 1644511149
transform 1 0 27048 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_290
timestamp 1644511149
transform 1 0 27784 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_296
timestamp 1644511149
transform 1 0 28336 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_304
timestamp 1644511149
transform 1 0 29072 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_309
timestamp 1644511149
transform 1 0 29532 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_316
timestamp 1644511149
transform 1 0 30176 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_7
timestamp 1644511149
transform 1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_14
timestamp 1644511149
transform 1 0 2392 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_26
timestamp 1644511149
transform 1 0 3496 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_38
timestamp 1644511149
transform 1 0 4600 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_50
timestamp 1644511149
transform 1 0 5704 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1644511149
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1644511149
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_93
timestamp 1644511149
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1644511149
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1644511149
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_113
timestamp 1644511149
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_125
timestamp 1644511149
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_137
timestamp 1644511149
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_149
timestamp 1644511149
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1644511149
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1644511149
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_186
timestamp 1644511149
transform 1 0 18216 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_198
timestamp 1644511149
transform 1 0 19320 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_218
timestamp 1644511149
transform 1 0 21160 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_225
timestamp 1644511149
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_237
timestamp 1644511149
transform 1 0 22908 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_245
timestamp 1644511149
transform 1 0 23644 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_257
timestamp 1644511149
transform 1 0 24748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_265
timestamp 1644511149
transform 1 0 25484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_277
timestamp 1644511149
transform 1 0 26588 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_95_281
timestamp 1644511149
transform 1 0 26956 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_292
timestamp 1644511149
transform 1 0 27968 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_300
timestamp 1644511149
transform 1 0 28704 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_306
timestamp 1644511149
transform 1 0 29256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_316
timestamp 1644511149
transform 1 0 30176 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_7
timestamp 1644511149
transform 1 0 1748 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_19
timestamp 1644511149
transform 1 0 2852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1644511149
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1644511149
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1644511149
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1644511149
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1644511149
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1644511149
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_97
timestamp 1644511149
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_109
timestamp 1644511149
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_121
timestamp 1644511149
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1644511149
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1644511149
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_141
timestamp 1644511149
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_153
timestamp 1644511149
transform 1 0 15180 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_157
timestamp 1644511149
transform 1 0 15548 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_161
timestamp 1644511149
transform 1 0 15916 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_168
timestamp 1644511149
transform 1 0 16560 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_180
timestamp 1644511149
transform 1 0 17664 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_192
timestamp 1644511149
transform 1 0 18768 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_197
timestamp 1644511149
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_209
timestamp 1644511149
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_221
timestamp 1644511149
transform 1 0 21436 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_227
timestamp 1644511149
transform 1 0 21988 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_248
timestamp 1644511149
transform 1 0 23920 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_263
timestamp 1644511149
transform 1 0 25300 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_269
timestamp 1644511149
transform 1 0 25852 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_276
timestamp 1644511149
transform 1 0 26496 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_284
timestamp 1644511149
transform 1 0 27232 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_96_292
timestamp 1644511149
transform 1 0 27968 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_304
timestamp 1644511149
transform 1 0 29072 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_309
timestamp 1644511149
transform 1 0 29532 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_316
timestamp 1644511149
transform 1 0 30176 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_7
timestamp 1644511149
transform 1 0 1748 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_14
timestamp 1644511149
transform 1 0 2392 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_26
timestamp 1644511149
transform 1 0 3496 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_38
timestamp 1644511149
transform 1 0 4600 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_50
timestamp 1644511149
transform 1 0 5704 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_93
timestamp 1644511149
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1644511149
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1644511149
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_113
timestamp 1644511149
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_125
timestamp 1644511149
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_137
timestamp 1644511149
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_149
timestamp 1644511149
transform 1 0 14812 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_157
timestamp 1644511149
transform 1 0 15548 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_164
timestamp 1644511149
transform 1 0 16192 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_169
timestamp 1644511149
transform 1 0 16652 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_173
timestamp 1644511149
transform 1 0 17020 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_178
timestamp 1644511149
transform 1 0 17480 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_185
timestamp 1644511149
transform 1 0 18124 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_197
timestamp 1644511149
transform 1 0 19228 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_208
timestamp 1644511149
transform 1 0 20240 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_216
timestamp 1644511149
transform 1 0 20976 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_97_225
timestamp 1644511149
transform 1 0 21804 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_229
timestamp 1644511149
transform 1 0 22172 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_236
timestamp 1644511149
transform 1 0 22816 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_247
timestamp 1644511149
transform 1 0 23828 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_259
timestamp 1644511149
transform 1 0 24932 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_271
timestamp 1644511149
transform 1 0 26036 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1644511149
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_287
timestamp 1644511149
transform 1 0 27508 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_293
timestamp 1644511149
transform 1 0 28060 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_303
timestamp 1644511149
transform 1 0 28980 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_316
timestamp 1644511149
transform 1 0 30176 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_98_3
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_9
timestamp 1644511149
transform 1 0 1932 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_21
timestamp 1644511149
transform 1 0 3036 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1644511149
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1644511149
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1644511149
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1644511149
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1644511149
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1644511149
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_85
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_97
timestamp 1644511149
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_109
timestamp 1644511149
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_121
timestamp 1644511149
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1644511149
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1644511149
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_141
timestamp 1644511149
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_153
timestamp 1644511149
transform 1 0 15180 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_168
timestamp 1644511149
transform 1 0 16560 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_192
timestamp 1644511149
transform 1 0 18768 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_197
timestamp 1644511149
transform 1 0 19228 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_221
timestamp 1644511149
transform 1 0 21436 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_241
timestamp 1644511149
transform 1 0 23276 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_249
timestamp 1644511149
transform 1 0 24012 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_261
timestamp 1644511149
transform 1 0 25116 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_272
timestamp 1644511149
transform 1 0 26128 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_290
timestamp 1644511149
transform 1 0 27784 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_304
timestamp 1644511149
transform 1 0 29072 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_309
timestamp 1644511149
transform 1 0 29532 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_316
timestamp 1644511149
transform 1 0 30176 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_7
timestamp 1644511149
transform 1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_14
timestamp 1644511149
transform 1 0 2392 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_26
timestamp 1644511149
transform 1 0 3496 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_38
timestamp 1644511149
transform 1 0 4600 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_50
timestamp 1644511149
transform 1 0 5704 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1644511149
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1644511149
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_93
timestamp 1644511149
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1644511149
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1644511149
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_113
timestamp 1644511149
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_125
timestamp 1644511149
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_137
timestamp 1644511149
transform 1 0 13708 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_148
timestamp 1644511149
transform 1 0 14720 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_152
timestamp 1644511149
transform 1 0 15088 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_156
timestamp 1644511149
transform 1 0 15456 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_164
timestamp 1644511149
transform 1 0 16192 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_169
timestamp 1644511149
transform 1 0 16652 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_189
timestamp 1644511149
transform 1 0 18492 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_213
timestamp 1644511149
transform 1 0 20700 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_221
timestamp 1644511149
transform 1 0 21436 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_241
timestamp 1644511149
transform 1 0 23276 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_249
timestamp 1644511149
transform 1 0 24012 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_257
timestamp 1644511149
transform 1 0 24748 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_265
timestamp 1644511149
transform 1 0 25484 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_274
timestamp 1644511149
transform 1 0 26312 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_291
timestamp 1644511149
transform 1 0 27876 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_295
timestamp 1644511149
transform 1 0 28244 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_302
timestamp 1644511149
transform 1 0 28888 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_316
timestamp 1644511149
transform 1 0 30176 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_7
timestamp 1644511149
transform 1 0 1748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_14
timestamp 1644511149
transform 1 0 2392 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 1644511149
transform 1 0 3496 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1644511149
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1644511149
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1644511149
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1644511149
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1644511149
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_97
timestamp 1644511149
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_109
timestamp 1644511149
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_121
timestamp 1644511149
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_136
timestamp 1644511149
transform 1 0 13616 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_157
timestamp 1644511149
transform 1 0 15548 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_161
timestamp 1644511149
transform 1 0 15916 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_165
timestamp 1644511149
transform 1 0 16284 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_178
timestamp 1644511149
transform 1 0 17480 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_192
timestamp 1644511149
transform 1 0 18768 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_213
timestamp 1644511149
transform 1 0 20700 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_225
timestamp 1644511149
transform 1 0 21804 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_237
timestamp 1644511149
transform 1 0 22908 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1644511149
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1644511149
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_260
timestamp 1644511149
transform 1 0 25024 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_266
timestamp 1644511149
transform 1 0 25576 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_273
timestamp 1644511149
transform 1 0 26220 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_100_290
timestamp 1644511149
transform 1 0 27784 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_304
timestamp 1644511149
transform 1 0 29072 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_313
timestamp 1644511149
transform 1 0 29900 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_319
timestamp 1644511149
transform 1 0 30452 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_7
timestamp 1644511149
transform 1 0 1748 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_14
timestamp 1644511149
transform 1 0 2392 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_26
timestamp 1644511149
transform 1 0 3496 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_38
timestamp 1644511149
transform 1 0 4600 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_50
timestamp 1644511149
transform 1 0 5704 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_93
timestamp 1644511149
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1644511149
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1644511149
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_113
timestamp 1644511149
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_125
timestamp 1644511149
transform 1 0 12604 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_133
timestamp 1644511149
transform 1 0 13340 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_143
timestamp 1644511149
transform 1 0 14260 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_164
timestamp 1644511149
transform 1 0 16192 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_169
timestamp 1644511149
transform 1 0 16652 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_193
timestamp 1644511149
transform 1 0 18860 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_205
timestamp 1644511149
transform 1 0 19964 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1644511149
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1644511149
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_225
timestamp 1644511149
transform 1 0 21804 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_233
timestamp 1644511149
transform 1 0 22540 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_242
timestamp 1644511149
transform 1 0 23368 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_249
timestamp 1644511149
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_261
timestamp 1644511149
transform 1 0 25116 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_275
timestamp 1644511149
transform 1 0 26404 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1644511149
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_285
timestamp 1644511149
transform 1 0 27324 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_293
timestamp 1644511149
transform 1 0 28060 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_306
timestamp 1644511149
transform 1 0 29256 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_316
timestamp 1644511149
transform 1 0 30176 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_7
timestamp 1644511149
transform 1 0 1748 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_19
timestamp 1644511149
transform 1 0 2852 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1644511149
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1644511149
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1644511149
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1644511149
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1644511149
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1644511149
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1644511149
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1644511149
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_97
timestamp 1644511149
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_109
timestamp 1644511149
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_121
timestamp 1644511149
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1644511149
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1644511149
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_141
timestamp 1644511149
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_157
timestamp 1644511149
transform 1 0 15548 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_170
timestamp 1644511149
transform 1 0 16744 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_183
timestamp 1644511149
transform 1 0 17940 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_191
timestamp 1644511149
transform 1 0 18676 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1644511149
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_197
timestamp 1644511149
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_209
timestamp 1644511149
transform 1 0 20332 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_217
timestamp 1644511149
transform 1 0 21068 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_229
timestamp 1644511149
transform 1 0 22172 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_241
timestamp 1644511149
transform 1 0 23276 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_102_249
timestamp 1644511149
transform 1 0 24012 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_253
timestamp 1644511149
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_265
timestamp 1644511149
transform 1 0 25484 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_102_277
timestamp 1644511149
transform 1 0 26588 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_285
timestamp 1644511149
transform 1 0 27324 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_289
timestamp 1644511149
transform 1 0 27692 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_294
timestamp 1644511149
transform 1 0 28152 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_304
timestamp 1644511149
transform 1 0 29072 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_315
timestamp 1644511149
transform 1 0 30084 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_319
timestamp 1644511149
transform 1 0 30452 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_7
timestamp 1644511149
transform 1 0 1748 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_19
timestamp 1644511149
transform 1 0 2852 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_31
timestamp 1644511149
transform 1 0 3956 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_43
timestamp 1644511149
transform 1 0 5060 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1644511149
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1644511149
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1644511149
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1644511149
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_93
timestamp 1644511149
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1644511149
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1644511149
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_113
timestamp 1644511149
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_125
timestamp 1644511149
transform 1 0 12604 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_103_136
timestamp 1644511149
transform 1 0 13616 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_148
timestamp 1644511149
transform 1 0 14720 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_164
timestamp 1644511149
transform 1 0 16192 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_178
timestamp 1644511149
transform 1 0 17480 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_190
timestamp 1644511149
transform 1 0 18584 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_196
timestamp 1644511149
transform 1 0 19136 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_103_203
timestamp 1644511149
transform 1 0 19780 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_103_215
timestamp 1644511149
transform 1 0 20884 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1644511149
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_225
timestamp 1644511149
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_237
timestamp 1644511149
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_249
timestamp 1644511149
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_261
timestamp 1644511149
transform 1 0 25116 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_269
timestamp 1644511149
transform 1 0 25852 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_103_274
timestamp 1644511149
transform 1 0 26312 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_103_281
timestamp 1644511149
transform 1 0 26956 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_285
timestamp 1644511149
transform 1 0 27324 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_294
timestamp 1644511149
transform 1 0 28152 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_298
timestamp 1644511149
transform 1 0 28520 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_303
timestamp 1644511149
transform 1 0 28980 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_316
timestamp 1644511149
transform 1 0 30176 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1644511149
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1644511149
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1644511149
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1644511149
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1644511149
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1644511149
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1644511149
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1644511149
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1644511149
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_85
timestamp 1644511149
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_97
timestamp 1644511149
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_109
timestamp 1644511149
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_121
timestamp 1644511149
transform 1 0 12236 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_104_129
timestamp 1644511149
transform 1 0 12972 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_104_136
timestamp 1644511149
transform 1 0 13616 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_141
timestamp 1644511149
transform 1 0 14076 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_145
timestamp 1644511149
transform 1 0 14444 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_150
timestamp 1644511149
transform 1 0 14904 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_162
timestamp 1644511149
transform 1 0 16008 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_174
timestamp 1644511149
transform 1 0 17112 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_180
timestamp 1644511149
transform 1 0 17664 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_185
timestamp 1644511149
transform 1 0 18124 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_193
timestamp 1644511149
transform 1 0 18860 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_197
timestamp 1644511149
transform 1 0 19228 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_104_205
timestamp 1644511149
transform 1 0 19964 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_211
timestamp 1644511149
transform 1 0 20516 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_216
timestamp 1644511149
transform 1 0 20976 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_228
timestamp 1644511149
transform 1 0 22080 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_240
timestamp 1644511149
transform 1 0 23184 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_253
timestamp 1644511149
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_265
timestamp 1644511149
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_104_277
timestamp 1644511149
transform 1 0 26588 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_104_290
timestamp 1644511149
transform 1 0 27784 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_104_304
timestamp 1644511149
transform 1 0 29072 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_309
timestamp 1644511149
transform 1 0 29532 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_316
timestamp 1644511149
transform 1 0 30176 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_6
timestamp 1644511149
transform 1 0 1656 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_18
timestamp 1644511149
transform 1 0 2760 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_30
timestamp 1644511149
transform 1 0 3864 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_42
timestamp 1644511149
transform 1 0 4968 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_54
timestamp 1644511149
transform 1 0 6072 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1644511149
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1644511149
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1644511149
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_93
timestamp 1644511149
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1644511149
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1644511149
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_113
timestamp 1644511149
transform 1 0 11500 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_105_121
timestamp 1644511149
transform 1 0 12236 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_129
timestamp 1644511149
transform 1 0 12972 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_137
timestamp 1644511149
transform 1 0 13708 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_144
timestamp 1644511149
transform 1 0 14352 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_156
timestamp 1644511149
transform 1 0 15456 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_172
timestamp 1644511149
transform 1 0 16928 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_184
timestamp 1644511149
transform 1 0 18032 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_196
timestamp 1644511149
transform 1 0 19136 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_214
timestamp 1644511149
transform 1 0 20792 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_222
timestamp 1644511149
transform 1 0 21528 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_225
timestamp 1644511149
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_243
timestamp 1644511149
transform 1 0 23460 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_250
timestamp 1644511149
transform 1 0 24104 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_262
timestamp 1644511149
transform 1 0 25208 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_105_270
timestamp 1644511149
transform 1 0 25944 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_278
timestamp 1644511149
transform 1 0 26680 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_281
timestamp 1644511149
transform 1 0 26956 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_285
timestamp 1644511149
transform 1 0 27324 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_294
timestamp 1644511149
transform 1 0 28152 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_105_306
timestamp 1644511149
transform 1 0 29256 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_316
timestamp 1644511149
transform 1 0 30176 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_6
timestamp 1644511149
transform 1 0 1656 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_18
timestamp 1644511149
transform 1 0 2760 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_26
timestamp 1644511149
transform 1 0 3496 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1644511149
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1644511149
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1644511149
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1644511149
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1644511149
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1644511149
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1644511149
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_97
timestamp 1644511149
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_109
timestamp 1644511149
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_121
timestamp 1644511149
transform 1 0 12236 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_129
timestamp 1644511149
transform 1 0 12972 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_137
timestamp 1644511149
transform 1 0 13708 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_106_150
timestamp 1644511149
transform 1 0 14904 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_106_176
timestamp 1644511149
transform 1 0 17296 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_183
timestamp 1644511149
transform 1 0 17940 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1644511149
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_205
timestamp 1644511149
transform 1 0 19964 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_213
timestamp 1644511149
transform 1 0 20700 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_106_232
timestamp 1644511149
transform 1 0 22448 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_236
timestamp 1644511149
transform 1 0 22816 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_243
timestamp 1644511149
transform 1 0 23460 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_251
timestamp 1644511149
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_253
timestamp 1644511149
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_265
timestamp 1644511149
transform 1 0 25484 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_272
timestamp 1644511149
transform 1 0 26128 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_284
timestamp 1644511149
transform 1 0 27232 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_288
timestamp 1644511149
transform 1 0 27600 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_106_299
timestamp 1644511149
transform 1 0 28612 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_307
timestamp 1644511149
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_106_309
timestamp 1644511149
transform 1 0 29532 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_106_316
timestamp 1644511149
transform 1 0 30176 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_6
timestamp 1644511149
transform 1 0 1656 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_18
timestamp 1644511149
transform 1 0 2760 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_30
timestamp 1644511149
transform 1 0 3864 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_42
timestamp 1644511149
transform 1 0 4968 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_54
timestamp 1644511149
transform 1 0 6072 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1644511149
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1644511149
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1644511149
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_93
timestamp 1644511149
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1644511149
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1644511149
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_113
timestamp 1644511149
transform 1 0 11500 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_121
timestamp 1644511149
transform 1 0 12236 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_129
timestamp 1644511149
transform 1 0 12972 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_141
timestamp 1644511149
transform 1 0 14076 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_107_162
timestamp 1644511149
transform 1 0 16008 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_107_169
timestamp 1644511149
transform 1 0 16652 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_189
timestamp 1644511149
transform 1 0 18492 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_201
timestamp 1644511149
transform 1 0 19596 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_209
timestamp 1644511149
transform 1 0 20332 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_220
timestamp 1644511149
transform 1 0 21344 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_225
timestamp 1644511149
transform 1 0 21804 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_233
timestamp 1644511149
transform 1 0 22540 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_242
timestamp 1644511149
transform 1 0 23368 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_252
timestamp 1644511149
transform 1 0 24288 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_262
timestamp 1644511149
transform 1 0 25208 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_107_276
timestamp 1644511149
transform 1 0 26496 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_287
timestamp 1644511149
transform 1 0 27508 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_291
timestamp 1644511149
transform 1 0 27876 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_296
timestamp 1644511149
transform 1 0 28336 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_107_306
timestamp 1644511149
transform 1 0 29256 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_316
timestamp 1644511149
transform 1 0 30176 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_6
timestamp 1644511149
transform 1 0 1656 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_18
timestamp 1644511149
transform 1 0 2760 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_26
timestamp 1644511149
transform 1 0 3496 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1644511149
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1644511149
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1644511149
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1644511149
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1644511149
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1644511149
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_85
timestamp 1644511149
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_97
timestamp 1644511149
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_109
timestamp 1644511149
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_121
timestamp 1644511149
transform 1 0 12236 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_125
timestamp 1644511149
transform 1 0 12604 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_129
timestamp 1644511149
transform 1 0 12972 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_108_137
timestamp 1644511149
transform 1 0 13708 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_108_146
timestamp 1644511149
transform 1 0 14536 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_108_172
timestamp 1644511149
transform 1 0 16928 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_184
timestamp 1644511149
transform 1 0 18032 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_188
timestamp 1644511149
transform 1 0 18400 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_192
timestamp 1644511149
transform 1 0 18768 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_197
timestamp 1644511149
transform 1 0 19228 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_205
timestamp 1644511149
transform 1 0 19964 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_217
timestamp 1644511149
transform 1 0 21068 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_229
timestamp 1644511149
transform 1 0 22172 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_247
timestamp 1644511149
transform 1 0 23828 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_251
timestamp 1644511149
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_263
timestamp 1644511149
transform 1 0 25300 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_108_275
timestamp 1644511149
transform 1 0 26404 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_283
timestamp 1644511149
transform 1 0 27140 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_292
timestamp 1644511149
transform 1 0 27968 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_108_304
timestamp 1644511149
transform 1 0 29072 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_315
timestamp 1644511149
transform 1 0 30084 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_319
timestamp 1644511149
transform 1 0 30452 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_6
timestamp 1644511149
transform 1 0 1656 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_18
timestamp 1644511149
transform 1 0 2760 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_30
timestamp 1644511149
transform 1 0 3864 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_42
timestamp 1644511149
transform 1 0 4968 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_54
timestamp 1644511149
transform 1 0 6072 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1644511149
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1644511149
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1644511149
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_93
timestamp 1644511149
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1644511149
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1644511149
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_113
timestamp 1644511149
transform 1 0 11500 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_109_121
timestamp 1644511149
transform 1 0 12236 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_129
timestamp 1644511149
transform 1 0 12972 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_141
timestamp 1644511149
transform 1 0 14076 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_149
timestamp 1644511149
transform 1 0 14812 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_158
timestamp 1644511149
transform 1 0 15640 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_166
timestamp 1644511149
transform 1 0 16376 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_109_179
timestamp 1644511149
transform 1 0 17572 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_187
timestamp 1644511149
transform 1 0 18308 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_205
timestamp 1644511149
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_217
timestamp 1644511149
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_223
timestamp 1644511149
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_109_233
timestamp 1644511149
transform 1 0 22540 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_109_242
timestamp 1644511149
transform 1 0 23368 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_252
timestamp 1644511149
transform 1 0 24288 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_262
timestamp 1644511149
transform 1 0 25208 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_266
timestamp 1644511149
transform 1 0 25576 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_109_273
timestamp 1644511149
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_279
timestamp 1644511149
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_109_289
timestamp 1644511149
transform 1 0 27692 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_293
timestamp 1644511149
transform 1 0 28060 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_109_298
timestamp 1644511149
transform 1 0 28520 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_109_312
timestamp 1644511149
transform 1 0 29808 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1644511149
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1644511149
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1644511149
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1644511149
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1644511149
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1644511149
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1644511149
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1644511149
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1644511149
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_85
timestamp 1644511149
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_97
timestamp 1644511149
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_109
timestamp 1644511149
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_121
timestamp 1644511149
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1644511149
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1644511149
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_110_141
timestamp 1644511149
transform 1 0 14076 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_147
timestamp 1644511149
transform 1 0 14628 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_152
timestamp 1644511149
transform 1 0 15088 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_110_168
timestamp 1644511149
transform 1 0 16560 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_110_192
timestamp 1644511149
transform 1 0 18768 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_110_197
timestamp 1644511149
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_209
timestamp 1644511149
transform 1 0 20332 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_110_233
timestamp 1644511149
transform 1 0 22540 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_110_247
timestamp 1644511149
transform 1 0 23828 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_251
timestamp 1644511149
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_110_253
timestamp 1644511149
transform 1 0 24380 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_260
timestamp 1644511149
transform 1 0 25024 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_272
timestamp 1644511149
transform 1 0 26128 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_110_288
timestamp 1644511149
transform 1 0 27600 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_110_296
timestamp 1644511149
transform 1 0 28336 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_110_304
timestamp 1644511149
transform 1 0 29072 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_315
timestamp 1644511149
transform 1 0 30084 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_319
timestamp 1644511149
transform 1 0 30452 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_6
timestamp 1644511149
transform 1 0 1656 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_18
timestamp 1644511149
transform 1 0 2760 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_30
timestamp 1644511149
transform 1 0 3864 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_42
timestamp 1644511149
transform 1 0 4968 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_54
timestamp 1644511149
transform 1 0 6072 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1644511149
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1644511149
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1644511149
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_93
timestamp 1644511149
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1644511149
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1644511149
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_113
timestamp 1644511149
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_130
timestamp 1644511149
transform 1 0 13064 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_142
timestamp 1644511149
transform 1 0 14168 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_154
timestamp 1644511149
transform 1 0 15272 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_166
timestamp 1644511149
transform 1 0 16376 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_111_169
timestamp 1644511149
transform 1 0 16652 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_111_183
timestamp 1644511149
transform 1 0 17940 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_195
timestamp 1644511149
transform 1 0 19044 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_111_201
timestamp 1644511149
transform 1 0 19596 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_212
timestamp 1644511149
transform 1 0 20608 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_225
timestamp 1644511149
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_237
timestamp 1644511149
transform 1 0 22908 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_243
timestamp 1644511149
transform 1 0 23460 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_248
timestamp 1644511149
transform 1 0 23920 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_260
timestamp 1644511149
transform 1 0 25024 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_272
timestamp 1644511149
transform 1 0 26128 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_111_285
timestamp 1644511149
transform 1 0 27324 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_111_297
timestamp 1644511149
transform 1 0 28428 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_111_305
timestamp 1644511149
transform 1 0 29164 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_111_316
timestamp 1644511149
transform 1 0 30176 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_6
timestamp 1644511149
transform 1 0 1656 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_18
timestamp 1644511149
transform 1 0 2760 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_112_26
timestamp 1644511149
transform 1 0 3496 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_112_29
timestamp 1644511149
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_41
timestamp 1644511149
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_53
timestamp 1644511149
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_65
timestamp 1644511149
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1644511149
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1644511149
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_85
timestamp 1644511149
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_97
timestamp 1644511149
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_109
timestamp 1644511149
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_121
timestamp 1644511149
transform 1 0 12236 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_112_132
timestamp 1644511149
transform 1 0 13248 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_112_150
timestamp 1644511149
transform 1 0 14904 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_112_158
timestamp 1644511149
transform 1 0 15640 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_166
timestamp 1644511149
transform 1 0 16376 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_171
timestamp 1644511149
transform 1 0 16836 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_183
timestamp 1644511149
transform 1 0 17940 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1644511149
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_112_197
timestamp 1644511149
transform 1 0 19228 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_112_212
timestamp 1644511149
transform 1 0 20608 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_224
timestamp 1644511149
transform 1 0 21712 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_112_236
timestamp 1644511149
transform 1 0 22816 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_240
timestamp 1644511149
transform 1 0 23184 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_244
timestamp 1644511149
transform 1 0 23552 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_112_253
timestamp 1644511149
transform 1 0 24380 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_112_265
timestamp 1644511149
transform 1 0 25484 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_112_273
timestamp 1644511149
transform 1 0 26220 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_112_283
timestamp 1644511149
transform 1 0 27140 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_112_289
timestamp 1644511149
transform 1 0 27692 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_112_293
timestamp 1644511149
transform 1 0 28060 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_112_304
timestamp 1644511149
transform 1 0 29072 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_112_309
timestamp 1644511149
transform 1 0 29532 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_316
timestamp 1644511149
transform 1 0 30176 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_6
timestamp 1644511149
transform 1 0 1656 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_18
timestamp 1644511149
transform 1 0 2760 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_30
timestamp 1644511149
transform 1 0 3864 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_42
timestamp 1644511149
transform 1 0 4968 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_54
timestamp 1644511149
transform 1 0 6072 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1644511149
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1644511149
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1644511149
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_93
timestamp 1644511149
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1644511149
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1644511149
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_113
timestamp 1644511149
transform 1 0 11500 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_117
timestamp 1644511149
transform 1 0 11868 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_123
timestamp 1644511149
transform 1 0 12420 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_113_132
timestamp 1644511149
transform 1 0 13248 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_138
timestamp 1644511149
transform 1 0 13800 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_148
timestamp 1644511149
transform 1 0 14720 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_160
timestamp 1644511149
transform 1 0 15824 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_113_169
timestamp 1644511149
transform 1 0 16652 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_177
timestamp 1644511149
transform 1 0 17388 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_189
timestamp 1644511149
transform 1 0 18492 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_113_201
timestamp 1644511149
transform 1 0 19596 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_206
timestamp 1644511149
transform 1 0 20056 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_113_214
timestamp 1644511149
transform 1 0 20792 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_222
timestamp 1644511149
transform 1 0 21528 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_225
timestamp 1644511149
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_237
timestamp 1644511149
transform 1 0 22908 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_241
timestamp 1644511149
transform 1 0 23276 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_113_248
timestamp 1644511149
transform 1 0 23920 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_256
timestamp 1644511149
transform 1 0 24656 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_113_269
timestamp 1644511149
transform 1 0 25852 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_277
timestamp 1644511149
transform 1 0 26588 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_113_289
timestamp 1644511149
transform 1 0 27692 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_293
timestamp 1644511149
transform 1 0 28060 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_303
timestamp 1644511149
transform 1 0 28980 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_316
timestamp 1644511149
transform 1 0 30176 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_114_6
timestamp 1644511149
transform 1 0 1656 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_18
timestamp 1644511149
transform 1 0 2760 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_114_26
timestamp 1644511149
transform 1 0 3496 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1644511149
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1644511149
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1644511149
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1644511149
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1644511149
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1644511149
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_85
timestamp 1644511149
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_97
timestamp 1644511149
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_109
timestamp 1644511149
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_121
timestamp 1644511149
transform 1 0 12236 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_114_125
timestamp 1644511149
transform 1 0 12604 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_131
timestamp 1644511149
transform 1 0 13156 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1644511149
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_141
timestamp 1644511149
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_153
timestamp 1644511149
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_165
timestamp 1644511149
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_177
timestamp 1644511149
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1644511149
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1644511149
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_114_200
timestamp 1644511149
transform 1 0 19504 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_114_208
timestamp 1644511149
transform 1 0 20240 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_114_216
timestamp 1644511149
transform 1 0 20976 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_226
timestamp 1644511149
transform 1 0 21896 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_238
timestamp 1644511149
transform 1 0 23000 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_248
timestamp 1644511149
transform 1 0 23920 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_114_253
timestamp 1644511149
transform 1 0 24380 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_262
timestamp 1644511149
transform 1 0 25208 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_114_266
timestamp 1644511149
transform 1 0 25576 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_114_273
timestamp 1644511149
transform 1 0 26220 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_286
timestamp 1644511149
transform 1 0 27416 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_114_300
timestamp 1644511149
transform 1 0 28704 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_114_309
timestamp 1644511149
transform 1 0 29532 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_316
timestamp 1644511149
transform 1 0 30176 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_3
timestamp 1644511149
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_15
timestamp 1644511149
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_27
timestamp 1644511149
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_39
timestamp 1644511149
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1644511149
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1644511149
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1644511149
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1644511149
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1644511149
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_93
timestamp 1644511149
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_105
timestamp 1644511149
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1644511149
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_113
timestamp 1644511149
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_115_125
timestamp 1644511149
transform 1 0 12604 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_129
timestamp 1644511149
transform 1 0 12972 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_140
timestamp 1644511149
transform 1 0 13984 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_152
timestamp 1644511149
transform 1 0 15088 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_164
timestamp 1644511149
transform 1 0 16192 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_115_169
timestamp 1644511149
transform 1 0 16652 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_115_179
timestamp 1644511149
transform 1 0 17572 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_115_187
timestamp 1644511149
transform 1 0 18308 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_115_192
timestamp 1644511149
transform 1 0 18768 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_200
timestamp 1644511149
transform 1 0 19504 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_213
timestamp 1644511149
transform 1 0 20700 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_220
timestamp 1644511149
transform 1 0 21344 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_241
timestamp 1644511149
transform 1 0 23276 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_253
timestamp 1644511149
transform 1 0 24380 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_265
timestamp 1644511149
transform 1 0 25484 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_269
timestamp 1644511149
transform 1 0 25852 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_115_276
timestamp 1644511149
transform 1 0 26496 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_115_281
timestamp 1644511149
transform 1 0 26956 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_289
timestamp 1644511149
transform 1 0 27692 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_302
timestamp 1644511149
transform 1 0 28888 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_316
timestamp 1644511149
transform 1 0 30176 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_6
timestamp 1644511149
transform 1 0 1656 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_18
timestamp 1644511149
transform 1 0 2760 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_116_26
timestamp 1644511149
transform 1 0 3496 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_116_29
timestamp 1644511149
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_41
timestamp 1644511149
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_53
timestamp 1644511149
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_65
timestamp 1644511149
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1644511149
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1644511149
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1644511149
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_97
timestamp 1644511149
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_109
timestamp 1644511149
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_121
timestamp 1644511149
transform 1 0 12236 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_125
timestamp 1644511149
transform 1 0 12604 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_129
timestamp 1644511149
transform 1 0 12972 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_116_137
timestamp 1644511149
transform 1 0 13708 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_141
timestamp 1644511149
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_153
timestamp 1644511149
transform 1 0 15180 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_157
timestamp 1644511149
transform 1 0 15548 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_169
timestamp 1644511149
transform 1 0 16652 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_179
timestamp 1644511149
transform 1 0 17572 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_116_186
timestamp 1644511149
transform 1 0 18216 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_116_194
timestamp 1644511149
transform 1 0 18952 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_116_200
timestamp 1644511149
transform 1 0 19504 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_116_213
timestamp 1644511149
transform 1 0 20700 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_219
timestamp 1644511149
transform 1 0 21252 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_236
timestamp 1644511149
transform 1 0 22816 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_248
timestamp 1644511149
transform 1 0 23920 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_116_253
timestamp 1644511149
transform 1 0 24380 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_116_269
timestamp 1644511149
transform 1 0 25852 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_281
timestamp 1644511149
transform 1 0 26956 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_285
timestamp 1644511149
transform 1 0 27324 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_294
timestamp 1644511149
transform 1 0 28152 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_116_302
timestamp 1644511149
transform 1 0 28888 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_116_309
timestamp 1644511149
transform 1 0 29532 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_316
timestamp 1644511149
transform 1 0 30176 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_117_6
timestamp 1644511149
transform 1 0 1656 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_18
timestamp 1644511149
transform 1 0 2760 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_30
timestamp 1644511149
transform 1 0 3864 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_42
timestamp 1644511149
transform 1 0 4968 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_54
timestamp 1644511149
transform 1 0 6072 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1644511149
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1644511149
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1644511149
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_93
timestamp 1644511149
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1644511149
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1644511149
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_113
timestamp 1644511149
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_130
timestamp 1644511149
transform 1 0 13064 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_136
timestamp 1644511149
transform 1 0 13616 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_153
timestamp 1644511149
transform 1 0 15180 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_117_164
timestamp 1644511149
transform 1 0 16192 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_169
timestamp 1644511149
transform 1 0 16652 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_117_190
timestamp 1644511149
transform 1 0 18584 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_198
timestamp 1644511149
transform 1 0 19320 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_117_220
timestamp 1644511149
transform 1 0 21344 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_117_233
timestamp 1644511149
transform 1 0 22540 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_247
timestamp 1644511149
transform 1 0 23828 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_259
timestamp 1644511149
transform 1 0 24932 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_266
timestamp 1644511149
transform 1 0 25576 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_278
timestamp 1644511149
transform 1 0 26680 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_117_281
timestamp 1644511149
transform 1 0 26956 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_289
timestamp 1644511149
transform 1 0 27692 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_117_295
timestamp 1644511149
transform 1 0 28244 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_303
timestamp 1644511149
transform 1 0 28980 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_316
timestamp 1644511149
transform 1 0 30176 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_6
timestamp 1644511149
transform 1 0 1656 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_18
timestamp 1644511149
transform 1 0 2760 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_118_26
timestamp 1644511149
transform 1 0 3496 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1644511149
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1644511149
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1644511149
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1644511149
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1644511149
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1644511149
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_85
timestamp 1644511149
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_97
timestamp 1644511149
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_109
timestamp 1644511149
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_121
timestamp 1644511149
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1644511149
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1644511149
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_149
timestamp 1644511149
transform 1 0 14812 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_153
timestamp 1644511149
transform 1 0 15180 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_170
timestamp 1644511149
transform 1 0 16744 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_182
timestamp 1644511149
transform 1 0 17848 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1644511149
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1644511149
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_200
timestamp 1644511149
transform 1 0 19504 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_208
timestamp 1644511149
transform 1 0 20240 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_214
timestamp 1644511149
transform 1 0 20792 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_226
timestamp 1644511149
transform 1 0 21896 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_230
timestamp 1644511149
transform 1 0 22264 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_237
timestamp 1644511149
transform 1 0 22908 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_247
timestamp 1644511149
transform 1 0 23828 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1644511149
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_259
timestamp 1644511149
transform 1 0 24932 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_118_269
timestamp 1644511149
transform 1 0 25852 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_118_283
timestamp 1644511149
transform 1 0 27140 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_297
timestamp 1644511149
transform 1 0 28428 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_305
timestamp 1644511149
transform 1 0 29164 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_118_309
timestamp 1644511149
transform 1 0 29532 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_316
timestamp 1644511149
transform 1 0 30176 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_6
timestamp 1644511149
transform 1 0 1656 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_18
timestamp 1644511149
transform 1 0 2760 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_30
timestamp 1644511149
transform 1 0 3864 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_42
timestamp 1644511149
transform 1 0 4968 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_54
timestamp 1644511149
transform 1 0 6072 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1644511149
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1644511149
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1644511149
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_93
timestamp 1644511149
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1644511149
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1644511149
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_113
timestamp 1644511149
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_130
timestamp 1644511149
transform 1 0 13064 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_142
timestamp 1644511149
transform 1 0 14168 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_148
timestamp 1644511149
transform 1 0 14720 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_157
timestamp 1644511149
transform 1 0 15548 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_165
timestamp 1644511149
transform 1 0 16284 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_169
timestamp 1644511149
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_181
timestamp 1644511149
transform 1 0 17756 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_189
timestamp 1644511149
transform 1 0 18492 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_199
timestamp 1644511149
transform 1 0 19412 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_211
timestamp 1644511149
transform 1 0 20516 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1644511149
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_225
timestamp 1644511149
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_237
timestamp 1644511149
transform 1 0 22908 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_119_247
timestamp 1644511149
transform 1 0 23828 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_255
timestamp 1644511149
transform 1 0 24564 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_264
timestamp 1644511149
transform 1 0 25392 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_119_274
timestamp 1644511149
transform 1 0 26312 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_289
timestamp 1644511149
transform 1 0 27692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_301
timestamp 1644511149
transform 1 0 28796 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_308
timestamp 1644511149
transform 1 0 29440 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_316
timestamp 1644511149
transform 1 0 30176 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_120_6
timestamp 1644511149
transform 1 0 1656 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_18
timestamp 1644511149
transform 1 0 2760 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_26
timestamp 1644511149
transform 1 0 3496 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1644511149
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1644511149
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1644511149
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1644511149
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1644511149
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1644511149
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_85
timestamp 1644511149
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_97
timestamp 1644511149
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_109
timestamp 1644511149
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_121
timestamp 1644511149
transform 1 0 12236 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_125
timestamp 1644511149
transform 1 0 12604 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_131
timestamp 1644511149
transform 1 0 13156 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1644511149
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_141
timestamp 1644511149
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_153
timestamp 1644511149
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_165
timestamp 1644511149
transform 1 0 16284 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_172
timestamp 1644511149
transform 1 0 16928 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_120_180
timestamp 1644511149
transform 1 0 17664 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_186
timestamp 1644511149
transform 1 0 18216 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_190
timestamp 1644511149
transform 1 0 18584 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_120_197
timestamp 1644511149
transform 1 0 19228 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_225
timestamp 1644511149
transform 1 0 21804 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_237
timestamp 1644511149
transform 1 0 22908 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_249
timestamp 1644511149
transform 1 0 24012 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_253
timestamp 1644511149
transform 1 0 24380 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_257
timestamp 1644511149
transform 1 0 24748 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_264
timestamp 1644511149
transform 1 0 25392 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_272
timestamp 1644511149
transform 1 0 26128 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_281
timestamp 1644511149
transform 1 0 26956 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_120_293
timestamp 1644511149
transform 1 0 28060 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_299
timestamp 1644511149
transform 1 0 28612 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_304
timestamp 1644511149
transform 1 0 29072 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_120_309
timestamp 1644511149
transform 1 0 29532 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_316
timestamp 1644511149
transform 1 0 30176 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_3
timestamp 1644511149
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_15
timestamp 1644511149
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_27
timestamp 1644511149
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_39
timestamp 1644511149
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1644511149
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1644511149
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1644511149
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1644511149
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1644511149
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_93
timestamp 1644511149
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1644511149
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1644511149
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_113
timestamp 1644511149
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_125
timestamp 1644511149
transform 1 0 12604 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_121_134
timestamp 1644511149
transform 1 0 13432 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_146
timestamp 1644511149
transform 1 0 14536 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_158
timestamp 1644511149
transform 1 0 15640 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_166
timestamp 1644511149
transform 1 0 16376 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_121_169
timestamp 1644511149
transform 1 0 16652 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_121_179
timestamp 1644511149
transform 1 0 17572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_191
timestamp 1644511149
transform 1 0 18676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_121_201
timestamp 1644511149
transform 1 0 19596 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_121_214
timestamp 1644511149
transform 1 0 20792 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_222
timestamp 1644511149
transform 1 0 21528 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_225
timestamp 1644511149
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_237
timestamp 1644511149
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_249
timestamp 1644511149
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_261
timestamp 1644511149
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1644511149
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1644511149
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_289
timestamp 1644511149
transform 1 0 27692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_301
timestamp 1644511149
transform 1 0 28796 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_121_309
timestamp 1644511149
transform 1 0 29532 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_316
timestamp 1644511149
transform 1 0 30176 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_6
timestamp 1644511149
transform 1 0 1656 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_18
timestamp 1644511149
transform 1 0 2760 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_26
timestamp 1644511149
transform 1 0 3496 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1644511149
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1644511149
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_53
timestamp 1644511149
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_65
timestamp 1644511149
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1644511149
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1644511149
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_85
timestamp 1644511149
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_97
timestamp 1644511149
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_109
timestamp 1644511149
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_121
timestamp 1644511149
transform 1 0 12236 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_122_130
timestamp 1644511149
transform 1 0 13064 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_138
timestamp 1644511149
transform 1 0 13800 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_122_141
timestamp 1644511149
transform 1 0 14076 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_122_155
timestamp 1644511149
transform 1 0 15364 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_167
timestamp 1644511149
transform 1 0 16468 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_171
timestamp 1644511149
transform 1 0 16836 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_181
timestamp 1644511149
transform 1 0 17756 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_122_191
timestamp 1644511149
transform 1 0 18676 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1644511149
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_197
timestamp 1644511149
transform 1 0 19228 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_203
timestamp 1644511149
transform 1 0 19780 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_213
timestamp 1644511149
transform 1 0 20700 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_221
timestamp 1644511149
transform 1 0 21436 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_228
timestamp 1644511149
transform 1 0 22080 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_240
timestamp 1644511149
transform 1 0 23184 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_253
timestamp 1644511149
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_265
timestamp 1644511149
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_277
timestamp 1644511149
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_289
timestamp 1644511149
transform 1 0 27692 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_297
timestamp 1644511149
transform 1 0 28428 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_304
timestamp 1644511149
transform 1 0 29072 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_122_309
timestamp 1644511149
transform 1 0 29532 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_316
timestamp 1644511149
transform 1 0 30176 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_6
timestamp 1644511149
transform 1 0 1656 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_18
timestamp 1644511149
transform 1 0 2760 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_30
timestamp 1644511149
transform 1 0 3864 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_42
timestamp 1644511149
transform 1 0 4968 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_54
timestamp 1644511149
transform 1 0 6072 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1644511149
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1644511149
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1644511149
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_93
timestamp 1644511149
transform 1 0 9660 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1644511149
transform 1 0 10764 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1644511149
transform 1 0 11316 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_113
timestamp 1644511149
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_125
timestamp 1644511149
transform 1 0 12604 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_123_132
timestamp 1644511149
transform 1 0 13248 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_138
timestamp 1644511149
transform 1 0 13800 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_155
timestamp 1644511149
transform 1 0 15364 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1644511149
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_123_169
timestamp 1644511149
transform 1 0 16652 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_123_181
timestamp 1644511149
transform 1 0 17756 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_201
timestamp 1644511149
transform 1 0 19596 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_123_209
timestamp 1644511149
transform 1 0 20332 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_215
timestamp 1644511149
transform 1 0 20884 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_220
timestamp 1644511149
transform 1 0 21344 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_233
timestamp 1644511149
transform 1 0 22540 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_245
timestamp 1644511149
transform 1 0 23644 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_257
timestamp 1644511149
transform 1 0 24748 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_269
timestamp 1644511149
transform 1 0 25852 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_277
timestamp 1644511149
transform 1 0 26588 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_281
timestamp 1644511149
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_293
timestamp 1644511149
transform 1 0 28060 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_301
timestamp 1644511149
transform 1 0 28796 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_123_308
timestamp 1644511149
transform 1 0 29440 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_316
timestamp 1644511149
transform 1 0 30176 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_6
timestamp 1644511149
transform 1 0 1656 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_18
timestamp 1644511149
transform 1 0 2760 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_124_26
timestamp 1644511149
transform 1 0 3496 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_124_29
timestamp 1644511149
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_41
timestamp 1644511149
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_53
timestamp 1644511149
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_65
timestamp 1644511149
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1644511149
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1644511149
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_85
timestamp 1644511149
transform 1 0 8924 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_97
timestamp 1644511149
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_109
timestamp 1644511149
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_121
timestamp 1644511149
transform 1 0 12236 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_124_132
timestamp 1644511149
transform 1 0 13248 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_124_141
timestamp 1644511149
transform 1 0 14076 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_147
timestamp 1644511149
transform 1 0 14628 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_124_165
timestamp 1644511149
transform 1 0 16284 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1644511149
transform 1 0 18492 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1644511149
transform 1 0 19044 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_124_206
timestamp 1644511149
transform 1 0 20056 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_226
timestamp 1644511149
transform 1 0 21896 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_124_246
timestamp 1644511149
transform 1 0 23736 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_124_253
timestamp 1644511149
transform 1 0 24380 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_265
timestamp 1644511149
transform 1 0 25484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_277
timestamp 1644511149
transform 1 0 26588 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_289
timestamp 1644511149
transform 1 0 27692 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1644511149
transform 1 0 28796 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1644511149
transform 1 0 29348 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_124_309
timestamp 1644511149
transform 1 0 29532 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_316
timestamp 1644511149
transform 1 0 30176 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_125_6
timestamp 1644511149
transform 1 0 1656 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_18
timestamp 1644511149
transform 1 0 2760 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_30
timestamp 1644511149
transform 1 0 3864 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_42
timestamp 1644511149
transform 1 0 4968 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_125_54
timestamp 1644511149
transform 1 0 6072 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1644511149
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1644511149
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1644511149
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_93
timestamp 1644511149
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1644511149
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1644511149
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_125_113
timestamp 1644511149
transform 1 0 11500 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_119
timestamp 1644511149
transform 1 0 12052 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_125_123
timestamp 1644511149
transform 1 0 12420 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_125_132
timestamp 1644511149
transform 1 0 13248 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_125_141
timestamp 1644511149
transform 1 0 14076 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_125_149
timestamp 1644511149
transform 1 0 14812 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_125_153
timestamp 1644511149
transform 1 0 15180 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_125_160
timestamp 1644511149
transform 1 0 15824 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_125_169
timestamp 1644511149
transform 1 0 16652 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_125_187
timestamp 1644511149
transform 1 0 18308 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_125_211
timestamp 1644511149
transform 1 0 20516 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_125_218
timestamp 1644511149
transform 1 0 21160 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_125_233
timestamp 1644511149
transform 1 0 22540 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_245
timestamp 1644511149
transform 1 0 23644 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_257
timestamp 1644511149
transform 1 0 24748 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_269
timestamp 1644511149
transform 1 0 25852 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_277
timestamp 1644511149
transform 1 0 26588 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_281
timestamp 1644511149
transform 1 0 26956 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_293
timestamp 1644511149
transform 1 0 28060 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_305
timestamp 1644511149
transform 1 0 29164 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_311
timestamp 1644511149
transform 1 0 29716 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_125_316
timestamp 1644511149
transform 1 0 30176 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_13
timestamp 1644511149
transform 1 0 2300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_126_25
timestamp 1644511149
transform 1 0 3404 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_126_29
timestamp 1644511149
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_41
timestamp 1644511149
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_53
timestamp 1644511149
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_65
timestamp 1644511149
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1644511149
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1644511149
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_85
timestamp 1644511149
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_97
timestamp 1644511149
transform 1 0 10028 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_109
timestamp 1644511149
transform 1 0 11132 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_121
timestamp 1644511149
transform 1 0 12236 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_126_132
timestamp 1644511149
transform 1 0 13248 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_126_141
timestamp 1644511149
transform 1 0 14076 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_126_152
timestamp 1644511149
transform 1 0 15088 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_158
timestamp 1644511149
transform 1 0 15640 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_126_168
timestamp 1644511149
transform 1 0 16560 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_126_192
timestamp 1644511149
transform 1 0 18768 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_126_197
timestamp 1644511149
transform 1 0 19228 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_221
timestamp 1644511149
transform 1 0 21436 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_233
timestamp 1644511149
transform 1 0 22540 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1644511149
transform 1 0 23644 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1644511149
transform 1 0 24196 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_253
timestamp 1644511149
transform 1 0 24380 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_265
timestamp 1644511149
transform 1 0 25484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_277
timestamp 1644511149
transform 1 0 26588 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_289
timestamp 1644511149
transform 1 0 27692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1644511149
transform 1 0 28796 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1644511149
transform 1 0 29348 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_126_309
timestamp 1644511149
transform 1 0 29532 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_126_316
timestamp 1644511149
transform 1 0 30176 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_127_3
timestamp 1644511149
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_15
timestamp 1644511149
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_27
timestamp 1644511149
transform 1 0 3588 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_39
timestamp 1644511149
transform 1 0 4692 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_51
timestamp 1644511149
transform 1 0 5796 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1644511149
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1644511149
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1644511149
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1644511149
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_93
timestamp 1644511149
transform 1 0 9660 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1644511149
transform 1 0 10764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1644511149
transform 1 0 11316 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_113
timestamp 1644511149
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_125
timestamp 1644511149
transform 1 0 12604 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_127_132
timestamp 1644511149
transform 1 0 13248 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_144
timestamp 1644511149
transform 1 0 14352 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_156
timestamp 1644511149
transform 1 0 15456 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_169
timestamp 1644511149
transform 1 0 16652 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_175
timestamp 1644511149
transform 1 0 17204 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_184
timestamp 1644511149
transform 1 0 18032 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_196
timestamp 1644511149
transform 1 0 19136 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_127_204
timestamp 1644511149
transform 1 0 19872 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_127_210
timestamp 1644511149
transform 1 0 20424 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_214
timestamp 1644511149
transform 1 0 20792 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_219
timestamp 1644511149
transform 1 0 21252 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_223
timestamp 1644511149
transform 1 0 21620 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_225
timestamp 1644511149
transform 1 0 21804 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_237
timestamp 1644511149
transform 1 0 22908 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_249
timestamp 1644511149
transform 1 0 24012 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_261
timestamp 1644511149
transform 1 0 25116 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_273
timestamp 1644511149
transform 1 0 26220 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_279
timestamp 1644511149
transform 1 0 26772 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_281
timestamp 1644511149
transform 1 0 26956 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_293
timestamp 1644511149
transform 1 0 28060 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_305
timestamp 1644511149
transform 1 0 29164 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_311
timestamp 1644511149
transform 1 0 29716 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_316
timestamp 1644511149
transform 1 0 30176 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_128_6
timestamp 1644511149
transform 1 0 1656 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_18
timestamp 1644511149
transform 1 0 2760 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_128_26
timestamp 1644511149
transform 1 0 3496 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_128_29
timestamp 1644511149
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1644511149
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_53
timestamp 1644511149
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_65
timestamp 1644511149
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1644511149
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1644511149
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_85
timestamp 1644511149
transform 1 0 8924 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_97
timestamp 1644511149
transform 1 0 10028 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_109
timestamp 1644511149
transform 1 0 11132 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_121
timestamp 1644511149
transform 1 0 12236 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_128_136
timestamp 1644511149
transform 1 0 13616 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_128_141
timestamp 1644511149
transform 1 0 14076 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_128_152
timestamp 1644511149
transform 1 0 15088 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_164
timestamp 1644511149
transform 1 0 16192 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_170
timestamp 1644511149
transform 1 0 16744 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_179
timestamp 1644511149
transform 1 0 17572 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_128_191
timestamp 1644511149
transform 1 0 18676 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_128_195
timestamp 1644511149
transform 1 0 19044 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_197
timestamp 1644511149
transform 1 0 19228 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_209
timestamp 1644511149
transform 1 0 20332 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_221
timestamp 1644511149
transform 1 0 21436 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_233
timestamp 1644511149
transform 1 0 22540 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_245
timestamp 1644511149
transform 1 0 23644 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_251
timestamp 1644511149
transform 1 0 24196 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_253
timestamp 1644511149
transform 1 0 24380 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_265
timestamp 1644511149
transform 1 0 25484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_277
timestamp 1644511149
transform 1 0 26588 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_289
timestamp 1644511149
transform 1 0 27692 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_301
timestamp 1644511149
transform 1 0 28796 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_307
timestamp 1644511149
transform 1 0 29348 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_128_309
timestamp 1644511149
transform 1 0 29532 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_316
timestamp 1644511149
transform 1 0 30176 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_6
timestamp 1644511149
transform 1 0 1656 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_18
timestamp 1644511149
transform 1 0 2760 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_30
timestamp 1644511149
transform 1 0 3864 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_42
timestamp 1644511149
transform 1 0 4968 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_54
timestamp 1644511149
transform 1 0 6072 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1644511149
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1644511149
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1644511149
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_93
timestamp 1644511149
transform 1 0 9660 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1644511149
transform 1 0 10764 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1644511149
transform 1 0 11316 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_113
timestamp 1644511149
transform 1 0 11500 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_125
timestamp 1644511149
transform 1 0 12604 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_137
timestamp 1644511149
transform 1 0 13708 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_129_145
timestamp 1644511149
transform 1 0 14444 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_129_152
timestamp 1644511149
transform 1 0 15088 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_129_164
timestamp 1644511149
transform 1 0 16192 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_169
timestamp 1644511149
transform 1 0 16652 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_177
timestamp 1644511149
transform 1 0 17388 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_189
timestamp 1644511149
transform 1 0 18492 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_201
timestamp 1644511149
transform 1 0 19596 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_213
timestamp 1644511149
transform 1 0 20700 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_129_221
timestamp 1644511149
transform 1 0 21436 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_225
timestamp 1644511149
transform 1 0 21804 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_237
timestamp 1644511149
transform 1 0 22908 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_249
timestamp 1644511149
transform 1 0 24012 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_261
timestamp 1644511149
transform 1 0 25116 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_273
timestamp 1644511149
transform 1 0 26220 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_279
timestamp 1644511149
transform 1 0 26772 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_281
timestamp 1644511149
transform 1 0 26956 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_293
timestamp 1644511149
transform 1 0 28060 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_305
timestamp 1644511149
transform 1 0 29164 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_311
timestamp 1644511149
transform 1 0 29716 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_129_316
timestamp 1644511149
transform 1 0 30176 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_130_6
timestamp 1644511149
transform 1 0 1656 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_18
timestamp 1644511149
transform 1 0 2760 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_130_26
timestamp 1644511149
transform 1 0 3496 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1644511149
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1644511149
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1644511149
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1644511149
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1644511149
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1644511149
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_85
timestamp 1644511149
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_97
timestamp 1644511149
transform 1 0 10028 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_109
timestamp 1644511149
transform 1 0 11132 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_121
timestamp 1644511149
transform 1 0 12236 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_133
timestamp 1644511149
transform 1 0 13340 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_139
timestamp 1644511149
transform 1 0 13892 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_130_141
timestamp 1644511149
transform 1 0 14076 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_130_152
timestamp 1644511149
transform 1 0 15088 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_130_161
timestamp 1644511149
transform 1 0 15916 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_169
timestamp 1644511149
transform 1 0 16652 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_178
timestamp 1644511149
transform 1 0 17480 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_130_186
timestamp 1644511149
transform 1 0 18216 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_130_192
timestamp 1644511149
transform 1 0 18768 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_130_197
timestamp 1644511149
transform 1 0 19228 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_130_205
timestamp 1644511149
transform 1 0 19964 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_130_214
timestamp 1644511149
transform 1 0 20792 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_226
timestamp 1644511149
transform 1 0 21896 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_238
timestamp 1644511149
transform 1 0 23000 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_130_250
timestamp 1644511149
transform 1 0 24104 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_130_253
timestamp 1644511149
transform 1 0 24380 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_265
timestamp 1644511149
transform 1 0 25484 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_277
timestamp 1644511149
transform 1 0 26588 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_289
timestamp 1644511149
transform 1 0 27692 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_301
timestamp 1644511149
transform 1 0 28796 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_307
timestamp 1644511149
transform 1 0 29348 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_130_309
timestamp 1644511149
transform 1 0 29532 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_130_316
timestamp 1644511149
transform 1 0 30176 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_131_6
timestamp 1644511149
transform 1 0 1656 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_18
timestamp 1644511149
transform 1 0 2760 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_30
timestamp 1644511149
transform 1 0 3864 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_42
timestamp 1644511149
transform 1 0 4968 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_54
timestamp 1644511149
transform 1 0 6072 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1644511149
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1644511149
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1644511149
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_93
timestamp 1644511149
transform 1 0 9660 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_105
timestamp 1644511149
transform 1 0 10764 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_111
timestamp 1644511149
transform 1 0 11316 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_113
timestamp 1644511149
transform 1 0 11500 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_125
timestamp 1644511149
transform 1 0 12604 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_140
timestamp 1644511149
transform 1 0 13984 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_152
timestamp 1644511149
transform 1 0 15088 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_164
timestamp 1644511149
transform 1 0 16192 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_131_177
timestamp 1644511149
transform 1 0 17388 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_131_191
timestamp 1644511149
transform 1 0 18676 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_195
timestamp 1644511149
transform 1 0 19044 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_131_205
timestamp 1644511149
transform 1 0 19964 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_211
timestamp 1644511149
transform 1 0 20516 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_131_220
timestamp 1644511149
transform 1 0 21344 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_131_225
timestamp 1644511149
transform 1 0 21804 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_237
timestamp 1644511149
transform 1 0 22908 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_249
timestamp 1644511149
transform 1 0 24012 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_261
timestamp 1644511149
transform 1 0 25116 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_273
timestamp 1644511149
transform 1 0 26220 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_279
timestamp 1644511149
transform 1 0 26772 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_281
timestamp 1644511149
transform 1 0 26956 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_293
timestamp 1644511149
transform 1 0 28060 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_305
timestamp 1644511149
transform 1 0 29164 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_311
timestamp 1644511149
transform 1 0 29716 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_131_316
timestamp 1644511149
transform 1 0 30176 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_132_3
timestamp 1644511149
transform 1 0 1380 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_15
timestamp 1644511149
transform 1 0 2484 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1644511149
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_29
timestamp 1644511149
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_41
timestamp 1644511149
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_53
timestamp 1644511149
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_65
timestamp 1644511149
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1644511149
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1644511149
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_85
timestamp 1644511149
transform 1 0 8924 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_97
timestamp 1644511149
transform 1 0 10028 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_109
timestamp 1644511149
transform 1 0 11132 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_121
timestamp 1644511149
transform 1 0 12236 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_133
timestamp 1644511149
transform 1 0 13340 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_139
timestamp 1644511149
transform 1 0 13892 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_132_141
timestamp 1644511149
transform 1 0 14076 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_132_145
timestamp 1644511149
transform 1 0 14444 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_151
timestamp 1644511149
transform 1 0 14996 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_132_159
timestamp 1644511149
transform 1 0 15732 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_132_170
timestamp 1644511149
transform 1 0 16744 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_132_179
timestamp 1644511149
transform 1 0 17572 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_132_192
timestamp 1644511149
transform 1 0 18768 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_132_206
timestamp 1644511149
transform 1 0 20056 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_132_213
timestamp 1644511149
transform 1 0 20700 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_132_217
timestamp 1644511149
transform 1 0 21068 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_235
timestamp 1644511149
transform 1 0 22724 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_247
timestamp 1644511149
transform 1 0 23828 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_132_251
timestamp 1644511149
transform 1 0 24196 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_253
timestamp 1644511149
transform 1 0 24380 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_265
timestamp 1644511149
transform 1 0 25484 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_277
timestamp 1644511149
transform 1 0 26588 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_289
timestamp 1644511149
transform 1 0 27692 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_301
timestamp 1644511149
transform 1 0 28796 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_307
timestamp 1644511149
transform 1 0 29348 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_132_309
timestamp 1644511149
transform 1 0 29532 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_316
timestamp 1644511149
transform 1 0 30176 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_133_6
timestamp 1644511149
transform 1 0 1656 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_18
timestamp 1644511149
transform 1 0 2760 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_30
timestamp 1644511149
transform 1 0 3864 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_42
timestamp 1644511149
transform 1 0 4968 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_54
timestamp 1644511149
transform 1 0 6072 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1644511149
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1644511149
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1644511149
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_93
timestamp 1644511149
transform 1 0 9660 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_105
timestamp 1644511149
transform 1 0 10764 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1644511149
transform 1 0 11316 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_113
timestamp 1644511149
transform 1 0 11500 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_125
timestamp 1644511149
transform 1 0 12604 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_137
timestamp 1644511149
transform 1 0 13708 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_133_150
timestamp 1644511149
transform 1 0 14904 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_133_159
timestamp 1644511149
transform 1 0 15732 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_133_167
timestamp 1644511149
transform 1 0 16468 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_133_178
timestamp 1644511149
transform 1 0 17480 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_133_202
timestamp 1644511149
transform 1 0 19688 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_210
timestamp 1644511149
transform 1 0 20424 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_133_220
timestamp 1644511149
transform 1 0 21344 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_133_241
timestamp 1644511149
transform 1 0 23276 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_253
timestamp 1644511149
transform 1 0 24380 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_265
timestamp 1644511149
transform 1 0 25484 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_277
timestamp 1644511149
transform 1 0 26588 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_133_281
timestamp 1644511149
transform 1 0 26956 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_293
timestamp 1644511149
transform 1 0 28060 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_305
timestamp 1644511149
transform 1 0 29164 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_311
timestamp 1644511149
transform 1 0 29716 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_133_316
timestamp 1644511149
transform 1 0 30176 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_134_6
timestamp 1644511149
transform 1 0 1656 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_18
timestamp 1644511149
transform 1 0 2760 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_134_26
timestamp 1644511149
transform 1 0 3496 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1644511149
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1644511149
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1644511149
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1644511149
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1644511149
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1644511149
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_85
timestamp 1644511149
transform 1 0 8924 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_97
timestamp 1644511149
transform 1 0 10028 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_109
timestamp 1644511149
transform 1 0 11132 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_121
timestamp 1644511149
transform 1 0 12236 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_133
timestamp 1644511149
transform 1 0 13340 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_139
timestamp 1644511149
transform 1 0 13892 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_134_141
timestamp 1644511149
transform 1 0 14076 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_149
timestamp 1644511149
transform 1 0 14812 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_134_170
timestamp 1644511149
transform 1 0 16744 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_134_191
timestamp 1644511149
transform 1 0 18676 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_134_195
timestamp 1644511149
transform 1 0 19044 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_134_197
timestamp 1644511149
transform 1 0 19228 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_134_220
timestamp 1644511149
transform 1 0 21344 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_232
timestamp 1644511149
transform 1 0 22448 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_244
timestamp 1644511149
transform 1 0 23552 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_134_253
timestamp 1644511149
transform 1 0 24380 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_265
timestamp 1644511149
transform 1 0 25484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_277
timestamp 1644511149
transform 1 0 26588 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_289
timestamp 1644511149
transform 1 0 27692 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_301
timestamp 1644511149
transform 1 0 28796 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_307
timestamp 1644511149
transform 1 0 29348 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_134_309
timestamp 1644511149
transform 1 0 29532 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_316
timestamp 1644511149
transform 1 0 30176 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_6
timestamp 1644511149
transform 1 0 1656 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_18
timestamp 1644511149
transform 1 0 2760 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_30
timestamp 1644511149
transform 1 0 3864 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_42
timestamp 1644511149
transform 1 0 4968 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_135_54
timestamp 1644511149
transform 1 0 6072 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1644511149
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1644511149
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1644511149
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_93
timestamp 1644511149
transform 1 0 9660 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_105
timestamp 1644511149
transform 1 0 10764 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_111
timestamp 1644511149
transform 1 0 11316 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_113
timestamp 1644511149
transform 1 0 11500 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_125
timestamp 1644511149
transform 1 0 12604 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_137
timestamp 1644511149
transform 1 0 13708 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_135_150
timestamp 1644511149
transform 1 0 14904 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_158
timestamp 1644511149
transform 1 0 15640 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_135_163
timestamp 1644511149
transform 1 0 16100 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_167
timestamp 1644511149
transform 1 0 16468 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_135_169
timestamp 1644511149
transform 1 0 16652 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_174
timestamp 1644511149
transform 1 0 17112 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_186
timestamp 1644511149
transform 1 0 18216 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_135_194
timestamp 1644511149
transform 1 0 18952 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_135_198
timestamp 1644511149
transform 1 0 19320 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_210
timestamp 1644511149
transform 1 0 20424 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_135_222
timestamp 1644511149
transform 1 0 21528 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_225
timestamp 1644511149
transform 1 0 21804 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_237
timestamp 1644511149
transform 1 0 22908 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_249
timestamp 1644511149
transform 1 0 24012 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_261
timestamp 1644511149
transform 1 0 25116 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_273
timestamp 1644511149
transform 1 0 26220 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_279
timestamp 1644511149
transform 1 0 26772 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_281
timestamp 1644511149
transform 1 0 26956 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_293
timestamp 1644511149
transform 1 0 28060 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_301
timestamp 1644511149
transform 1 0 28796 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_308
timestamp 1644511149
transform 1 0 29440 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_135_316
timestamp 1644511149
transform 1 0 30176 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_136_13
timestamp 1644511149
transform 1 0 2300 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_136_20
timestamp 1644511149
transform 1 0 2944 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_29
timestamp 1644511149
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_41
timestamp 1644511149
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_53
timestamp 1644511149
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_65
timestamp 1644511149
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1644511149
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1644511149
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_85
timestamp 1644511149
transform 1 0 8924 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_97
timestamp 1644511149
transform 1 0 10028 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_109
timestamp 1644511149
transform 1 0 11132 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_121
timestamp 1644511149
transform 1 0 12236 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_133
timestamp 1644511149
transform 1 0 13340 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_139
timestamp 1644511149
transform 1 0 13892 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_141
timestamp 1644511149
transform 1 0 14076 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_153
timestamp 1644511149
transform 1 0 15180 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_165
timestamp 1644511149
transform 1 0 16284 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_177
timestamp 1644511149
transform 1 0 17388 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_189
timestamp 1644511149
transform 1 0 18492 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_195
timestamp 1644511149
transform 1 0 19044 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_197
timestamp 1644511149
transform 1 0 19228 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_209
timestamp 1644511149
transform 1 0 20332 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_221
timestamp 1644511149
transform 1 0 21436 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_233
timestamp 1644511149
transform 1 0 22540 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_245
timestamp 1644511149
transform 1 0 23644 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_251
timestamp 1644511149
transform 1 0 24196 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_253
timestamp 1644511149
transform 1 0 24380 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_265
timestamp 1644511149
transform 1 0 25484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_277
timestamp 1644511149
transform 1 0 26588 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_289
timestamp 1644511149
transform 1 0 27692 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_136_297
timestamp 1644511149
transform 1 0 28428 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_304
timestamp 1644511149
transform 1 0 29072 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_136_309
timestamp 1644511149
transform 1 0 29532 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_316
timestamp 1644511149
transform 1 0 30176 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_13
timestamp 1644511149
transform 1 0 2300 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_27
timestamp 1644511149
transform 1 0 3588 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_39
timestamp 1644511149
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1644511149
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1644511149
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1644511149
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1644511149
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_81
timestamp 1644511149
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_93
timestamp 1644511149
transform 1 0 9660 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1644511149
transform 1 0 10764 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1644511149
transform 1 0 11316 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_113
timestamp 1644511149
transform 1 0 11500 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_125
timestamp 1644511149
transform 1 0 12604 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_137
timestamp 1644511149
transform 1 0 13708 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_149
timestamp 1644511149
transform 1 0 14812 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_161
timestamp 1644511149
transform 1 0 15916 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_167
timestamp 1644511149
transform 1 0 16468 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_169
timestamp 1644511149
transform 1 0 16652 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_181
timestamp 1644511149
transform 1 0 17756 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_193
timestamp 1644511149
transform 1 0 18860 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_205
timestamp 1644511149
transform 1 0 19964 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_217
timestamp 1644511149
transform 1 0 21068 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_223
timestamp 1644511149
transform 1 0 21620 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_225
timestamp 1644511149
transform 1 0 21804 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_237
timestamp 1644511149
transform 1 0 22908 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_249
timestamp 1644511149
transform 1 0 24012 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_261
timestamp 1644511149
transform 1 0 25116 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_273
timestamp 1644511149
transform 1 0 26220 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_279
timestamp 1644511149
transform 1 0 26772 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_281
timestamp 1644511149
transform 1 0 26956 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_293
timestamp 1644511149
transform 1 0 28060 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_300
timestamp 1644511149
transform 1 0 28704 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_308
timestamp 1644511149
transform 1 0 29440 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_316
timestamp 1644511149
transform 1 0 30176 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_13
timestamp 1644511149
transform 1 0 2300 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_25
timestamp 1644511149
transform 1 0 3404 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_39
timestamp 1644511149
transform 1 0 4692 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_51
timestamp 1644511149
transform 1 0 5796 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_55
timestamp 1644511149
transform 1 0 6164 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_57
timestamp 1644511149
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_69
timestamp 1644511149
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1644511149
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_85
timestamp 1644511149
transform 1 0 8924 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_97
timestamp 1644511149
transform 1 0 10028 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_109
timestamp 1644511149
transform 1 0 11132 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_113
timestamp 1644511149
transform 1 0 11500 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_125
timestamp 1644511149
transform 1 0 12604 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_137
timestamp 1644511149
transform 1 0 13708 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_141
timestamp 1644511149
transform 1 0 14076 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_153
timestamp 1644511149
transform 1 0 15180 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_165
timestamp 1644511149
transform 1 0 16284 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_169
timestamp 1644511149
transform 1 0 16652 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_181
timestamp 1644511149
transform 1 0 17756 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_193
timestamp 1644511149
transform 1 0 18860 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_197
timestamp 1644511149
transform 1 0 19228 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_209
timestamp 1644511149
transform 1 0 20332 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_221
timestamp 1644511149
transform 1 0 21436 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_225
timestamp 1644511149
transform 1 0 21804 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_237
timestamp 1644511149
transform 1 0 22908 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_249
timestamp 1644511149
transform 1 0 24012 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_253
timestamp 1644511149
transform 1 0 24380 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_265
timestamp 1644511149
transform 1 0 25484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_277
timestamp 1644511149
transform 1 0 26588 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_138_281
timestamp 1644511149
transform 1 0 26956 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_288
timestamp 1644511149
transform 1 0 27600 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_296
timestamp 1644511149
transform 1 0 28336 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_304
timestamp 1644511149
transform 1 0 29072 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_138_309
timestamp 1644511149
transform 1 0 29532 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_316
timestamp 1644511149
transform 1 0 30176 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 30820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 30820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 30820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 30820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 30820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 30820 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 30820 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 30820 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 30820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 30820 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 30820 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 30820 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 30820 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 30820 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 30820 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 30820 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 30820 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 30820 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 30820 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 30820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 30820 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 30820 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 30820 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 30820 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 30820 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 30820 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 30820 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 30820 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 30820 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 30820 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 30820 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 30820 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 30820 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 30820 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 30820 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 30820 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 30820 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 30820 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 30820 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 30820 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 30820 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 30820 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 30820 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 30820 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 30820 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 30820 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 30820 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 30820 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 30820 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 30820 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 30820 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 30820 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 30820 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 30820 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 30820 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 30820 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 30820 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1644511149
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1644511149
transform -1 0 30820 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1644511149
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1644511149
transform -1 0 30820 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1644511149
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1644511149
transform -1 0 30820 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1644511149
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1644511149
transform -1 0 30820 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1644511149
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1644511149
transform -1 0 30820 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1644511149
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1644511149
transform -1 0 30820 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1644511149
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1644511149
transform -1 0 30820 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1644511149
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1644511149
transform -1 0 30820 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1644511149
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1644511149
transform -1 0 30820 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1644511149
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1644511149
transform -1 0 30820 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1644511149
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1644511149
transform -1 0 30820 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1644511149
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1644511149
transform -1 0 30820 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1644511149
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1644511149
transform -1 0 30820 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1644511149
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1644511149
transform -1 0 30820 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1644511149
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1644511149
transform -1 0 30820 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1644511149
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1644511149
transform -1 0 30820 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1644511149
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1644511149
transform -1 0 30820 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1644511149
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1644511149
transform -1 0 30820 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1644511149
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1644511149
transform -1 0 30820 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1644511149
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1644511149
transform -1 0 30820 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1644511149
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1644511149
transform -1 0 30820 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1644511149
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1644511149
transform -1 0 30820 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1644511149
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1644511149
transform -1 0 30820 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1644511149
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1644511149
transform -1 0 30820 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1644511149
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1644511149
transform -1 0 30820 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1644511149
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1644511149
transform -1 0 30820 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1644511149
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1644511149
transform -1 0 30820 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1644511149
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1644511149
transform -1 0 30820 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1644511149
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1644511149
transform -1 0 30820 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1644511149
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1644511149
transform -1 0 30820 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1644511149
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1644511149
transform -1 0 30820 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1644511149
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1644511149
transform -1 0 30820 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1644511149
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1644511149
transform -1 0 30820 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1644511149
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1644511149
transform -1 0 30820 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1644511149
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1644511149
transform -1 0 30820 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1644511149
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1644511149
transform -1 0 30820 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1644511149
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1644511149
transform -1 0 30820 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 19136 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 24288 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 29440 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 21712 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 26864 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 19136 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 24288 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 29440 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 21712 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 26864 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 13984 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 19136 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 24288 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 29440 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 11408 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 16560 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 21712 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 26864 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 13984 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 19136 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 24288 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 29440 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 11408 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 16560 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 21712 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 26864 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 13984 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 19136 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 24288 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 29440 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 11408 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 16560 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 21712 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 26864 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 13984 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 19136 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 24288 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 29440 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 11408 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 16560 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 21712 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 26864 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 13984 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 19136 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 24288 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 29440 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 11408 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 16560 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 21712 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 26864 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 11408 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 13984 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 16560 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 19136 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 21712 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 24288 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 26864 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 29440 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0878_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _0880_
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0882_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18400 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0883_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19320 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _0884_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0885_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19872 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0890_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0892_
timestamp 1644511149
transform 1 0 24932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24196 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _0896_
timestamp 1644511149
transform 1 0 16100 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0898_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0899_
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0900_
timestamp 1644511149
transform 1 0 17848 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19412 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0903_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0904_
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0905_
timestamp 1644511149
transform 1 0 19872 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _0906_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0909_
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1644511149
transform 1 0 20884 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0912_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0913_
timestamp 1644511149
transform 1 0 21160 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0914_
timestamp 1644511149
transform 1 0 20516 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0915_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0916_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0917_
timestamp 1644511149
transform 1 0 20516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20700 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0919_
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0920_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0921_
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0922_
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0923_
timestamp 1644511149
transform 1 0 16836 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0924_
timestamp 1644511149
transform 1 0 17480 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0925_
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0926_
timestamp 1644511149
transform 1 0 17020 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0928_
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 1644511149
transform 1 0 1656 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0930_
timestamp 1644511149
transform 1 0 1564 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0931_
timestamp 1644511149
transform 1 0 17296 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0932_
timestamp 1644511149
transform 1 0 2392 0 1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0933_
timestamp 1644511149
transform 1 0 17848 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1644511149
transform 1 0 1564 0 -1 50048
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0935_
timestamp 1644511149
transform 1 0 17204 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0936_
timestamp 1644511149
transform 1 0 1564 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0937_
timestamp 1644511149
transform 1 0 17112 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0938_
timestamp 1644511149
transform 1 0 14996 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0939_
timestamp 1644511149
transform 1 0 14904 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0940_
timestamp 1644511149
transform 1 0 15180 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1644511149
transform 1 0 1564 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0942_
timestamp 1644511149
transform 1 0 14260 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1644511149
transform 1 0 2392 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 1644511149
transform 1 0 2392 0 1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1644511149
transform 1 0 14444 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0946_
timestamp 1644511149
transform 1 0 2392 0 -1 48960
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0947_
timestamp 1644511149
transform 1 0 14628 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1644511149
transform 1 0 2300 0 1 47872
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0949_
timestamp 1644511149
transform 1 0 14076 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1644511149
transform 1 0 2300 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1644511149
transform 1 0 15364 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0952_
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0953_
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0954_
timestamp 1644511149
transform 1 0 2300 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0955_
timestamp 1644511149
transform 1 0 12696 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1644511149
transform 1 0 2392 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1644511149
transform 1 0 1564 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1644511149
transform 1 0 12512 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0959_
timestamp 1644511149
transform 1 0 1564 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0960_
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0961_
timestamp 1644511149
transform 1 0 1564 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0962_
timestamp 1644511149
transform 1 0 11960 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 1644511149
transform 1 0 2392 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0964_
timestamp 1644511149
transform 1 0 11776 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0965_
timestamp 1644511149
transform 1 0 10304 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0966_
timestamp 1644511149
transform 1 0 10396 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1644511149
transform 1 0 1564 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0968_
timestamp 1644511149
transform 1 0 9660 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0969_
timestamp 1644511149
transform 1 0 8096 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0970_
timestamp 1644511149
transform 1 0 8372 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0971_
timestamp 1644511149
transform 1 0 9568 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0972_
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0973_
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0974_
timestamp 1644511149
transform 1 0 8004 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0975_
timestamp 1644511149
transform 1 0 9568 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0976_
timestamp 1644511149
transform 1 0 8280 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0977_
timestamp 1644511149
transform 1 0 9568 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0978_
timestamp 1644511149
transform 1 0 11776 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0979_
timestamp 1644511149
transform 1 0 13432 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1644511149
transform 1 0 8372 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0981_
timestamp 1644511149
transform 1 0 11316 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0982_
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0983_
timestamp 1644511149
transform 1 0 8832 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0984_
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0985_
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0986_
timestamp 1644511149
transform 1 0 12420 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1644511149
transform 1 0 8924 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0988_
timestamp 1644511149
transform 1 0 12788 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0989_
timestamp 1644511149
transform 1 0 8096 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0990_
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0991_
timestamp 1644511149
transform 1 0 12696 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0992_
timestamp 1644511149
transform 1 0 13800 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 1644511149
transform 1 0 8832 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0994_
timestamp 1644511149
transform 1 0 12512 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1644511149
transform 1 0 9476 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0996_
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0997_
timestamp 1644511149
transform 1 0 13524 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0998_
timestamp 1644511149
transform 1 0 10488 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0999_
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1000_
timestamp 1644511149
transform 1 0 9568 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1001_
timestamp 1644511149
transform 1 0 14076 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1002_
timestamp 1644511149
transform 1 0 9660 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1003_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1644511149
transform 1 0 9568 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1005_
timestamp 1644511149
transform 1 0 14996 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1006_
timestamp 1644511149
transform 1 0 2392 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1007_
timestamp 1644511149
transform 1 0 15456 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1010_
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1011_
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26496 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1013_
timestamp 1644511149
transform 1 0 23092 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _1014_
timestamp 1644511149
transform 1 0 20700 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1015_
timestamp 1644511149
transform 1 0 22632 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1016_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1017_
timestamp 1644511149
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1018_
timestamp 1644511149
transform 1 0 21804 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1019_
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1020_
timestamp 1644511149
transform 1 0 22816 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _1021_
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1022_
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1023_
timestamp 1644511149
transform 1 0 21988 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1024_
timestamp 1644511149
transform 1 0 22264 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1025_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1644511149
transform 1 0 22264 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1644511149
transform 1 0 24104 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1028_
timestamp 1644511149
transform 1 0 22724 0 1 40256
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1029_
timestamp 1644511149
transform 1 0 20700 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1644511149
transform 1 0 20424 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1644511149
transform 1 0 20056 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1032_
timestamp 1644511149
transform 1 0 17296 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1033_
timestamp 1644511149
transform 1 0 20424 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1644511149
transform 1 0 22264 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1035_
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1036_
timestamp 1644511149
transform 1 0 21896 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1037_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1038_
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1039_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1040_
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1041_
timestamp 1644511149
transform 1 0 21988 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1042_
timestamp 1644511149
transform 1 0 22816 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1644511149
transform 1 0 20792 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1044_
timestamp 1644511149
transform 1 0 22908 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1045_
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1046_
timestamp 1644511149
transform 1 0 23092 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1047_
timestamp 1644511149
transform 1 0 22172 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1048_
timestamp 1644511149
transform 1 0 20608 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1644511149
transform 1 0 25300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1050_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1051_
timestamp 1644511149
transform 1 0 22264 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1052_
timestamp 1644511149
transform 1 0 20792 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1644511149
transform 1 0 21804 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1054_
timestamp 1644511149
transform 1 0 20516 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1055_
timestamp 1644511149
transform 1 0 21804 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1056_
timestamp 1644511149
transform 1 0 22172 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1057_
timestamp 1644511149
transform 1 0 20792 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1058_
timestamp 1644511149
transform 1 0 20516 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1059_
timestamp 1644511149
transform 1 0 20608 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1060_
timestamp 1644511149
transform 1 0 20976 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1061_
timestamp 1644511149
transform 1 0 21160 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1644511149
transform 1 0 13340 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1063_
timestamp 1644511149
transform 1 0 12144 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1064_
timestamp 1644511149
transform 1 0 12788 0 -1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1644511149
transform 1 0 20608 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1644511149
transform 1 0 13616 0 -1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1644511149
transform 1 0 21804 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1644511149
transform 1 0 12788 0 1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1069_
timestamp 1644511149
transform 1 0 21804 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1070_
timestamp 1644511149
transform 1 0 12788 0 1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1071_
timestamp 1644511149
transform 1 0 21160 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1072_
timestamp 1644511149
transform 1 0 19964 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1073_
timestamp 1644511149
transform 1 0 12788 0 -1 71808
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1074_
timestamp 1644511149
transform 1 0 21804 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1075_
timestamp 1644511149
transform 1 0 20884 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1644511149
transform 1 0 13708 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 1644511149
transform 1 0 14444 0 -1 76160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1078_
timestamp 1644511149
transform 1 0 20608 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1644511149
transform 1 0 14352 0 1 75072
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1080_
timestamp 1644511149
transform 1 0 21804 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1644511149
transform 1 0 14444 0 -1 75072
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1644511149
transform 1 0 19688 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1644511149
transform 1 0 15272 0 -1 75072
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1644511149
transform 1 0 20608 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1085_
timestamp 1644511149
transform 1 0 16836 0 -1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1086_
timestamp 1644511149
transform 1 0 14536 0 1 73984
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1087_
timestamp 1644511149
transform 1 0 17940 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1088_
timestamp 1644511149
transform 1 0 16468 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1644511149
transform 1 0 13340 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1090_
timestamp 1644511149
transform 1 0 14628 0 -1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1091_
timestamp 1644511149
transform 1 0 17296 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1092_
timestamp 1644511149
transform 1 0 14628 0 1 71808
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1093_
timestamp 1644511149
transform 1 0 16836 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1094_
timestamp 1644511149
transform 1 0 14628 0 1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp 1644511149
transform 1 0 16652 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1644511149
transform 1 0 15456 0 1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1097_
timestamp 1644511149
transform 1 0 16744 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1098_
timestamp 1644511149
transform 1 0 16560 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1644511149
transform 1 0 14628 0 1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 1644511149
transform 1 0 17112 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1101_
timestamp 1644511149
transform 1 0 15180 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1644511149
transform 1 0 12696 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1103_
timestamp 1644511149
transform 1 0 12788 0 -1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1104_
timestamp 1644511149
transform 1 0 14628 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1644511149
transform 1 0 12696 0 1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1106_
timestamp 1644511149
transform 1 0 14812 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1644511149
transform 1 0 12604 0 1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1108_
timestamp 1644511149
transform 1 0 13800 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1644511149
transform 1 0 12604 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1110_
timestamp 1644511149
transform 1 0 14076 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1111_
timestamp 1644511149
transform 1 0 15824 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1644511149
transform 1 0 12604 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1113_
timestamp 1644511149
transform 1 0 13524 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1114_
timestamp 1644511149
transform 1 0 16652 0 -1 62016
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1115_
timestamp 1644511149
transform 1 0 12696 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1644511149
transform 1 0 12788 0 -1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1644511149
transform 1 0 13340 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1644511149
transform 1 0 12788 0 1 63104
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1119_
timestamp 1644511149
transform 1 0 14904 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1120_
timestamp 1644511149
transform 1 0 12696 0 1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1121_
timestamp 1644511149
transform 1 0 15824 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1644511149
transform 1 0 11960 0 -1 64192
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1644511149
transform 1 0 17296 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1124_
timestamp 1644511149
transform 1 0 17848 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1644511149
transform 1 0 12604 0 -1 63104
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1126_
timestamp 1644511149
transform 1 0 17204 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1644511149
transform 1 0 19596 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1128_
timestamp 1644511149
transform 1 0 12696 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1129_
timestamp 1644511149
transform 1 0 12512 0 -1 62016
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1130_
timestamp 1644511149
transform 1 0 18860 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1131_
timestamp 1644511149
transform 1 0 12512 0 -1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1132_
timestamp 1644511149
transform 1 0 19228 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1133_
timestamp 1644511149
transform 1 0 14076 0 1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1134_
timestamp 1644511149
transform 1 0 20332 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1644511149
transform 1 0 12512 0 1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1644511149
transform 1 0 19228 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1644511149
transform 1 0 12512 0 -1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1138_
timestamp 1644511149
transform 1 0 19504 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1139_
timestamp 1644511149
transform 1 0 13156 0 1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1140_
timestamp 1644511149
transform 1 0 21068 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1644511149
transform 1 0 13156 0 -1 58752
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1644511149
transform 1 0 22172 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1143_
timestamp 1644511149
transform 1 0 25576 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _1144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1145_
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1147_
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1148_
timestamp 1644511149
transform 1 0 27968 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1644511149
transform 1 0 27508 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1151_
timestamp 1644511149
transform 1 0 26956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26404 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1154_
timestamp 1644511149
transform 1 0 23460 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1155_
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _1156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1157_
timestamp 1644511149
transform 1 0 23552 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1158_
timestamp 1644511149
transform 1 0 23460 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1159_
timestamp 1644511149
transform 1 0 22356 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1162_
timestamp 1644511149
transform 1 0 25760 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1163_
timestamp 1644511149
transform 1 0 26772 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1164_
timestamp 1644511149
transform 1 0 27324 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1165_
timestamp 1644511149
transform 1 0 18216 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1166_
timestamp 1644511149
transform 1 0 25944 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1167_
timestamp 1644511149
transform 1 0 25852 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1168_
timestamp 1644511149
transform 1 0 20332 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1169_
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1172_
timestamp 1644511149
transform 1 0 16468 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1174_
timestamp 1644511149
transform 1 0 20792 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1175_
timestamp 1644511149
transform 1 0 19964 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1176_
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1177_
timestamp 1644511149
transform 1 0 23184 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1178_
timestamp 1644511149
transform 1 0 20976 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1179_
timestamp 1644511149
transform 1 0 23092 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1180_
timestamp 1644511149
transform 1 0 24288 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1181_
timestamp 1644511149
transform 1 0 22264 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1182_
timestamp 1644511149
transform 1 0 21988 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1183_
timestamp 1644511149
transform 1 0 27140 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1184_
timestamp 1644511149
transform 1 0 28060 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1185_
timestamp 1644511149
transform 1 0 29532 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27508 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1187_
timestamp 1644511149
transform 1 0 27140 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1188_
timestamp 1644511149
transform 1 0 26864 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1189__1
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190__5
timestamp 1644511149
transform 1 0 19964 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190__6
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190__7
timestamp 1644511149
transform 1 0 19228 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190__8
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190__9
timestamp 1644511149
transform 1 0 22908 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21712 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193__10
timestamp 1644511149
transform 1 0 22540 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193__11
timestamp 1644511149
transform 1 0 22356 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1194_
timestamp 1644511149
transform 1 0 21804 0 -1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1195_
timestamp 1644511149
transform 1 0 1656 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1196_
timestamp 1644511149
transform 1 0 20240 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1197_
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198__12
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198__13
timestamp 1644511149
transform 1 0 17848 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1199_
timestamp 1644511149
transform 1 0 29348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1200_
timestamp 1644511149
transform 1 0 28428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1201_
timestamp 1644511149
transform 1 0 29348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1202_
timestamp 1644511149
transform 1 0 29808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1203_
timestamp 1644511149
transform 1 0 28244 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1204_
timestamp 1644511149
transform 1 0 29808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1206_
timestamp 1644511149
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1207_
timestamp 1644511149
transform 1 0 29348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1208_
timestamp 1644511149
transform 1 0 28612 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1209_
timestamp 1644511149
transform 1 0 28152 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1210_
timestamp 1644511149
transform 1 0 27876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1211_
timestamp 1644511149
transform 1 0 28060 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1212_
timestamp 1644511149
transform 1 0 27324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1213_
timestamp 1644511149
transform 1 0 28244 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1214_
timestamp 1644511149
transform 1 0 28152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1215_
timestamp 1644511149
transform 1 0 27048 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1216_
timestamp 1644511149
transform 1 0 29808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1217_
timestamp 1644511149
transform 1 0 29808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1218_
timestamp 1644511149
transform 1 0 28244 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1219_
timestamp 1644511149
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1220_
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1221_
timestamp 1644511149
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1222_
timestamp 1644511149
transform 1 0 28244 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1224_
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1225_
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1226_
timestamp 1644511149
transform 1 0 27048 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1227_
timestamp 1644511149
transform 1 0 27784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1228_
timestamp 1644511149
transform 1 0 27968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1229_
timestamp 1644511149
transform 1 0 27048 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1230_
timestamp 1644511149
transform 1 0 26128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1231_
timestamp 1644511149
transform 1 0 27232 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1232_
timestamp 1644511149
transform 1 0 26496 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1233_
timestamp 1644511149
transform 1 0 26956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1234_
timestamp 1644511149
transform 1 0 27324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1235_
timestamp 1644511149
transform 1 0 27784 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1236_
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp 1644511149
transform 1 0 27048 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1238_
timestamp 1644511149
transform 1 0 27048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1239_
timestamp 1644511149
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1240_
timestamp 1644511149
transform 1 0 27968 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1241_
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1242_
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1243_
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1244_
timestamp 1644511149
transform 1 0 27048 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1245_
timestamp 1644511149
transform 1 0 2300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1246_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1247_
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1248_
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1250_
timestamp 1644511149
transform 1 0 26036 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1251_
timestamp 1644511149
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1252_
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1254_
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1256_
timestamp 1644511149
transform 1 0 29348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1257_
timestamp 1644511149
transform 1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1258_
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1260_
timestamp 1644511149
transform 1 0 29348 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1262_
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1263_
timestamp 1644511149
transform 1 0 26680 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1264_
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1265_
timestamp 1644511149
transform 1 0 28060 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1644511149
transform 1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1267_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1268_
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1269_
timestamp 1644511149
transform 1 0 26312 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1270_
timestamp 1644511149
transform 1 0 2116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1271_
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1272_
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1273_
timestamp 1644511149
transform 1 0 27232 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1274_
timestamp 1644511149
transform 1 0 29348 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1644511149
transform 1 0 2116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1276_
timestamp 1644511149
transform 1 0 29348 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1278_
timestamp 1644511149
transform 1 0 29348 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1280_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1282_
timestamp 1644511149
transform 1 0 25668 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1644511149
transform 1 0 2116 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1284_
timestamp 1644511149
transform 1 0 28152 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1285_
timestamp 1644511149
transform 1 0 26772 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1286_
timestamp 1644511149
transform 1 0 1656 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1287_
timestamp 1644511149
transform 1 0 27048 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1288_
timestamp 1644511149
transform 1 0 2116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1289_
timestamp 1644511149
transform 1 0 29072 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1290_
timestamp 1644511149
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1291_
timestamp 1644511149
transform 1 0 28980 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1293_
timestamp 1644511149
transform 1 0 27968 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1295_
timestamp 1644511149
transform 1 0 28152 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _1296_
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1297_
timestamp 1644511149
transform 1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_8  _1298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1644511149
transform 1 0 1656 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_8  _1300_
timestamp 1644511149
transform 1 0 27968 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1301_
timestamp 1644511149
transform 1 0 2116 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_8  _1302_
timestamp 1644511149
transform 1 0 28244 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1303_
timestamp 1644511149
transform 1 0 2116 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_8  _1304_
timestamp 1644511149
transform 1 0 28244 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1644511149
transform 1 0 2116 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1306_
timestamp 1644511149
transform 1 0 23000 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1307_
timestamp 1644511149
transform 1 0 28704 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1308_
timestamp 1644511149
transform 1 0 29348 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1309_
timestamp 1644511149
transform 1 0 1656 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1310_
timestamp 1644511149
transform 1 0 29348 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1311_
timestamp 1644511149
transform 1 0 2116 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1312_
timestamp 1644511149
transform 1 0 29348 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1313_
timestamp 1644511149
transform 1 0 2116 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1314_
timestamp 1644511149
transform 1 0 28152 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1315_
timestamp 1644511149
transform 1 0 2116 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1316_
timestamp 1644511149
transform 1 0 26128 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1317_
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1318_
timestamp 1644511149
transform 1 0 26772 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1319_
timestamp 1644511149
transform 1 0 22632 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1320_
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1322_
timestamp 1644511149
transform 1 0 27232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1323_
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1324_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1325_
timestamp 1644511149
transform 1 0 25576 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1326_
timestamp 1644511149
transform 1 0 25576 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1327_
timestamp 1644511149
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1328_
timestamp 1644511149
transform 1 0 26496 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1329_
timestamp 1644511149
transform 1 0 24656 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1330_
timestamp 1644511149
transform 1 0 23368 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1331_
timestamp 1644511149
transform 1 0 23276 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1332_
timestamp 1644511149
transform 1 0 25852 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1333_
timestamp 1644511149
transform 1 0 25760 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1334_
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1335_
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_1  _1336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25576 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1339_
timestamp 1644511149
transform 1 0 25668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1340_
timestamp 1644511149
transform 1 0 25668 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1341_
timestamp 1644511149
transform 1 0 25576 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1342_
timestamp 1644511149
transform 1 0 26036 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1343_
timestamp 1644511149
transform 1 0 24656 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1344_
timestamp 1644511149
transform 1 0 19596 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1345_
timestamp 1644511149
transform 1 0 23000 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1346_
timestamp 1644511149
transform 1 0 25668 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1347_
timestamp 1644511149
transform 1 0 24288 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_1  _1348_
timestamp 1644511149
transform 1 0 24932 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1349_
timestamp 1644511149
transform 1 0 24564 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1350_
timestamp 1644511149
transform 1 0 25208 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1351_
timestamp 1644511149
transform 1 0 24656 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1352_
timestamp 1644511149
transform 1 0 24840 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1353_
timestamp 1644511149
transform 1 0 24472 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1354_
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1355_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1644511149
transform 1 0 23736 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1358_
timestamp 1644511149
transform 1 0 28060 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1359_
timestamp 1644511149
transform 1 0 27324 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1360_
timestamp 1644511149
transform 1 0 27140 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1361_
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _1363_
timestamp 1644511149
transform 1 0 23092 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1364_
timestamp 1644511149
transform 1 0 27692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1365_
timestamp 1644511149
transform 1 0 28244 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1366_
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1367_
timestamp 1644511149
transform 1 0 28244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1368_
timestamp 1644511149
transform 1 0 23828 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1369_
timestamp 1644511149
transform 1 0 22816 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1644511149
transform 1 0 28244 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1371_
timestamp 1644511149
transform 1 0 27416 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1372_
timestamp 1644511149
transform 1 0 28336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1373_
timestamp 1644511149
transform 1 0 23736 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1375_
timestamp 1644511149
transform 1 0 27600 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1376_
timestamp 1644511149
transform 1 0 29348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1377_
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1378_
timestamp 1644511149
transform 1 0 23736 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1379_
timestamp 1644511149
transform 1 0 24380 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__a41o_1  _1380_
timestamp 1644511149
transform 1 0 25392 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1381_
timestamp 1644511149
transform 1 0 25208 0 -1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1382_
timestamp 1644511149
transform 1 0 25024 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1383_
timestamp 1644511149
transform 1 0 25760 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1384_
timestamp 1644511149
transform 1 0 25300 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1385_
timestamp 1644511149
transform 1 0 24380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1386_
timestamp 1644511149
transform 1 0 24748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1387_
timestamp 1644511149
transform 1 0 23828 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1389_
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1390_
timestamp 1644511149
transform 1 0 23368 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1391_
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1392_
timestamp 1644511149
transform 1 0 23276 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1393_
timestamp 1644511149
transform 1 0 24472 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1394_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1395_
timestamp 1644511149
transform 1 0 25116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1396_
timestamp 1644511149
transform 1 0 24840 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1397_
timestamp 1644511149
transform 1 0 24380 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1398_
timestamp 1644511149
transform 1 0 24564 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1399_
timestamp 1644511149
transform 1 0 22816 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1400_
timestamp 1644511149
transform 1 0 28060 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1401_
timestamp 1644511149
transform 1 0 29440 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1402_
timestamp 1644511149
transform 1 0 27784 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1403_
timestamp 1644511149
transform 1 0 29072 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1404_
timestamp 1644511149
transform 1 0 22908 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1644511149
transform 1 0 29624 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1406_
timestamp 1644511149
transform 1 0 28244 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1407_
timestamp 1644511149
transform 1 0 28060 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1408_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1409_
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1410_
timestamp 1644511149
transform 1 0 28796 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _1411_
timestamp 1644511149
transform 1 0 22908 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp 1644511149
transform 1 0 29716 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1413_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1414_
timestamp 1644511149
transform 1 0 29440 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1415_
timestamp 1644511149
transform 1 0 23276 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1416_
timestamp 1644511149
transform 1 0 23276 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1417_
timestamp 1644511149
transform 1 0 29716 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1418_
timestamp 1644511149
transform 1 0 27416 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1419_
timestamp 1644511149
transform 1 0 29440 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1420_
timestamp 1644511149
transform 1 0 24288 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1421_
timestamp 1644511149
transform 1 0 24104 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1422_
timestamp 1644511149
transform 1 0 24932 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1423_
timestamp 1644511149
transform 1 0 24104 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1424_
timestamp 1644511149
transform 1 0 24380 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1425_
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1426_
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1427_
timestamp 1644511149
transform 1 0 24472 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1428_
timestamp 1644511149
transform 1 0 24748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1429_
timestamp 1644511149
transform 1 0 23736 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1430_
timestamp 1644511149
transform 1 0 23276 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1431_
timestamp 1644511149
transform 1 0 25300 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1432_
timestamp 1644511149
transform 1 0 25576 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1433_
timestamp 1644511149
transform 1 0 25576 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1434_
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1435_
timestamp 1644511149
transform 1 0 24748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1436_
timestamp 1644511149
transform 1 0 23184 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1437_
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1438_
timestamp 1644511149
transform 1 0 24656 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1439_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1440_
timestamp 1644511149
transform 1 0 24472 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1441_
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1442_
timestamp 1644511149
transform 1 0 25208 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1443_
timestamp 1644511149
transform 1 0 25668 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1444_
timestamp 1644511149
transform 1 0 23276 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1445_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1446_
timestamp 1644511149
transform 1 0 27416 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1447_
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1448_
timestamp 1644511149
transform 1 0 23276 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1644511149
transform 1 0 28060 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1450_
timestamp 1644511149
transform 1 0 29716 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1451_
timestamp 1644511149
transform 1 0 29532 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1452_
timestamp 1644511149
transform 1 0 28336 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1453_
timestamp 1644511149
transform 1 0 22356 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1454_
timestamp 1644511149
transform 1 0 29716 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1455_
timestamp 1644511149
transform 1 0 28152 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1456_
timestamp 1644511149
transform 1 0 27968 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1457_
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1458_
timestamp 1644511149
transform 1 0 28336 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1459_
timestamp 1644511149
transform 1 0 28152 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__and2_2  _1460_
timestamp 1644511149
transform 1 0 24380 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1461_
timestamp 1644511149
transform 1 0 28336 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1462_
timestamp 1644511149
transform 1 0 27416 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1463_
timestamp 1644511149
transform 1 0 29440 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1464_
timestamp 1644511149
transform 1 0 24932 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1465_
timestamp 1644511149
transform 1 0 24196 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1466_
timestamp 1644511149
transform 1 0 23184 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1467_
timestamp 1644511149
transform 1 0 24564 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1468_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1469_
timestamp 1644511149
transform 1 0 24380 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1470_
timestamp 1644511149
transform 1 0 24104 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1471_
timestamp 1644511149
transform 1 0 25116 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1472_
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1473_
timestamp 1644511149
transform 1 0 25300 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1474_
timestamp 1644511149
transform 1 0 24380 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1475_
timestamp 1644511149
transform 1 0 25760 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1476_
timestamp 1644511149
transform 1 0 26036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1477_
timestamp 1644511149
transform 1 0 25208 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1478_
timestamp 1644511149
transform 1 0 25484 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1479_
timestamp 1644511149
transform 1 0 25852 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1644511149
transform 1 0 23092 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1481_
timestamp 1644511149
transform 1 0 23368 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1644511149
transform 1 0 29716 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1483_
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1484_
timestamp 1644511149
transform 1 0 29440 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1485_
timestamp 1644511149
transform 1 0 23368 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1486_
timestamp 1644511149
transform 1 0 29716 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1487_
timestamp 1644511149
transform 1 0 28520 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1488_
timestamp 1644511149
transform 1 0 28336 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1489_
timestamp 1644511149
transform 1 0 23276 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1490_
timestamp 1644511149
transform 1 0 27968 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1491_
timestamp 1644511149
transform 1 0 27324 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1492_
timestamp 1644511149
transform 1 0 28244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1493_
timestamp 1644511149
transform 1 0 23276 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1494_
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1495_
timestamp 1644511149
transform 1 0 27232 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1496_
timestamp 1644511149
transform 1 0 26864 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1497_
timestamp 1644511149
transform 1 0 27784 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1498_
timestamp 1644511149
transform 1 0 28152 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1499_
timestamp 1644511149
transform 1 0 28060 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1500_
timestamp 1644511149
transform 1 0 28520 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1501_
timestamp 1644511149
transform 1 0 27968 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1502_
timestamp 1644511149
transform 1 0 27416 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1503_
timestamp 1644511149
transform 1 0 27416 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1504_
timestamp 1644511149
transform 1 0 27140 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1505_
timestamp 1644511149
transform 1 0 25944 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1506_
timestamp 1644511149
transform 1 0 26220 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1507_
timestamp 1644511149
transform 1 0 27140 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1508_
timestamp 1644511149
transform 1 0 27048 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1509_
timestamp 1644511149
transform 1 0 26496 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1510_
timestamp 1644511149
transform 1 0 27416 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1511_
timestamp 1644511149
transform 1 0 26956 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1512_
timestamp 1644511149
transform 1 0 26496 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1513_
timestamp 1644511149
transform 1 0 25944 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1514_
timestamp 1644511149
transform 1 0 27048 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1515_
timestamp 1644511149
transform 1 0 25944 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1516_
timestamp 1644511149
transform 1 0 24380 0 1 60928
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1517_
timestamp 1644511149
transform 1 0 25392 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1518_
timestamp 1644511149
transform 1 0 27416 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1519_
timestamp 1644511149
transform 1 0 29808 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1520_
timestamp 1644511149
transform 1 0 26220 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1521_
timestamp 1644511149
transform 1 0 28152 0 1 55488
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1522_
timestamp 1644511149
transform 1 0 27232 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1523_
timestamp 1644511149
transform 1 0 28152 0 -1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1524_
timestamp 1644511149
transform 1 0 26496 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1525_
timestamp 1644511149
transform 1 0 28244 0 1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1526_
timestamp 1644511149
transform 1 0 27968 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1527_
timestamp 1644511149
transform 1 0 27600 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1528_
timestamp 1644511149
transform 1 0 28520 0 -1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1529_
timestamp 1644511149
transform 1 0 26864 0 1 55488
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1530_
timestamp 1644511149
transform 1 0 28336 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1531_
timestamp 1644511149
transform 1 0 28244 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1532_
timestamp 1644511149
transform 1 0 29348 0 -1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1533_
timestamp 1644511149
transform 1 0 26680 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1534_
timestamp 1644511149
transform 1 0 24564 0 1 63104
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1535_
timestamp 1644511149
transform 1 0 24656 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1536_
timestamp 1644511149
transform 1 0 27416 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1537_
timestamp 1644511149
transform 1 0 27784 0 1 64192
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1538_
timestamp 1644511149
transform 1 0 26864 0 1 58752
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1539_
timestamp 1644511149
transform 1 0 25944 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1540_
timestamp 1644511149
transform 1 0 24656 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1541_
timestamp 1644511149
transform 1 0 26864 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1542_
timestamp 1644511149
transform 1 0 26956 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1543_
timestamp 1644511149
transform 1 0 24472 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1544_
timestamp 1644511149
transform 1 0 26956 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1545_
timestamp 1644511149
transform 1 0 26956 0 -1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1546_
timestamp 1644511149
transform 1 0 25852 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1547_
timestamp 1644511149
transform 1 0 23736 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1548_
timestamp 1644511149
transform 1 0 27232 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1549_
timestamp 1644511149
transform 1 0 29256 0 -1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1550_
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1551_
timestamp 1644511149
transform 1 0 29348 0 -1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1552_
timestamp 1644511149
transform 1 0 28888 0 -1 62016
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1553_
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1554_
timestamp 1644511149
transform 1 0 28152 0 -1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1555_
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1556_
timestamp 1644511149
transform 1 0 29348 0 -1 54400
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1557_
timestamp 1644511149
transform 1 0 28336 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1558_
timestamp 1644511149
transform 1 0 28336 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1559_
timestamp 1644511149
transform 1 0 26956 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1560_
timestamp 1644511149
transform 1 0 25668 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1561_
timestamp 1644511149
transform 1 0 24932 0 -1 64192
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1562_
timestamp 1644511149
transform 1 0 24656 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1563_
timestamp 1644511149
transform 1 0 26956 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1564_
timestamp 1644511149
transform 1 0 25944 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1565_
timestamp 1644511149
transform 1 0 26864 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1566_
timestamp 1644511149
transform 1 0 27416 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1567_
timestamp 1644511149
transform 1 0 27508 0 1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1568_
timestamp 1644511149
transform 1 0 25576 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1569_
timestamp 1644511149
transform 1 0 24932 0 1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1570_
timestamp 1644511149
transform 1 0 24840 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1571_
timestamp 1644511149
transform 1 0 26220 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1572_
timestamp 1644511149
transform 1 0 26496 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1573_
timestamp 1644511149
transform 1 0 25760 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1574_
timestamp 1644511149
transform 1 0 25760 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1575_
timestamp 1644511149
transform 1 0 27324 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1576_
timestamp 1644511149
transform 1 0 28152 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1577_
timestamp 1644511149
transform 1 0 29532 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1578_
timestamp 1644511149
transform 1 0 29348 0 -1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1644511149
transform 1 0 29256 0 -1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1580_
timestamp 1644511149
transform 1 0 29532 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1581_
timestamp 1644511149
transform 1 0 29348 0 -1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1582_
timestamp 1644511149
transform 1 0 27968 0 -1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1583_
timestamp 1644511149
transform 1 0 29532 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1584_
timestamp 1644511149
transform 1 0 29348 0 -1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1585_
timestamp 1644511149
transform 1 0 28520 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1586_
timestamp 1644511149
transform 1 0 29348 0 -1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1587_
timestamp 1644511149
transform 1 0 25668 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1588_
timestamp 1644511149
transform 1 0 24840 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1589_
timestamp 1644511149
transform 1 0 26956 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1590_
timestamp 1644511149
transform 1 0 25852 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1591_
timestamp 1644511149
transform 1 0 25300 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1592_
timestamp 1644511149
transform 1 0 26956 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1593_
timestamp 1644511149
transform 1 0 25944 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1594_
timestamp 1644511149
transform 1 0 25024 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1595_
timestamp 1644511149
transform 1 0 26404 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1596_
timestamp 1644511149
transform 1 0 26956 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1597_
timestamp 1644511149
transform 1 0 25668 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1598_
timestamp 1644511149
transform 1 0 27692 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1599_
timestamp 1644511149
transform 1 0 28520 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1600_
timestamp 1644511149
transform 1 0 28152 0 -1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1601_
timestamp 1644511149
transform 1 0 28520 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1602_
timestamp 1644511149
transform 1 0 28244 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1603_
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1604_
timestamp 1644511149
transform 1 0 26588 0 1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1605_
timestamp 1644511149
transform 1 0 27600 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1606_
timestamp 1644511149
transform 1 0 27784 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1607_
timestamp 1644511149
transform 1 0 17296 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1608_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1609_
timestamp 1644511149
transform 1 0 23276 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1610_
timestamp 1644511149
transform 1 0 22724 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1644511149
transform 1 0 21804 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1612_
timestamp 1644511149
transform 1 0 19412 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1613_
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1614_
timestamp 1644511149
transform 1 0 17664 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1615_
timestamp 1644511149
transform 1 0 17756 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1616_
timestamp 1644511149
transform 1 0 19872 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1617_
timestamp 1644511149
transform 1 0 19228 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1618_
timestamp 1644511149
transform 1 0 18400 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1619_
timestamp 1644511149
transform 1 0 19228 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1620_
timestamp 1644511149
transform 1 0 18492 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1621_
timestamp 1644511149
transform 1 0 17664 0 -1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1622_
timestamp 1644511149
transform 1 0 19688 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1623_
timestamp 1644511149
transform 1 0 20424 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1624_
timestamp 1644511149
transform 1 0 19504 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1625_
timestamp 1644511149
transform 1 0 19228 0 1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1626_
timestamp 1644511149
transform 1 0 18308 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1627_
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1628_
timestamp 1644511149
transform 1 0 17020 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1629_
timestamp 1644511149
transform 1 0 17572 0 1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1630_
timestamp 1644511149
transform 1 0 17848 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1631_
timestamp 1644511149
transform 1 0 17848 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1632_
timestamp 1644511149
transform 1 0 17112 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1633_
timestamp 1644511149
transform 1 0 17112 0 1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1634_
timestamp 1644511149
transform 1 0 18492 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1635_
timestamp 1644511149
transform 1 0 16652 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1636_
timestamp 1644511149
transform 1 0 17664 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1637_
timestamp 1644511149
transform 1 0 15732 0 1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1638_
timestamp 1644511149
transform 1 0 16284 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1639_
timestamp 1644511149
transform 1 0 16652 0 -1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1640_
timestamp 1644511149
transform 1 0 16652 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1641_
timestamp 1644511149
transform 1 0 15640 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1642_
timestamp 1644511149
transform 1 0 15916 0 1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1643_
timestamp 1644511149
transform 1 0 15180 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1644_
timestamp 1644511149
transform 1 0 16008 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1645_
timestamp 1644511149
transform 1 0 17020 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1646_
timestamp 1644511149
transform 1 0 14076 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1647_
timestamp 1644511149
transform 1 0 14076 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1648_
timestamp 1644511149
transform 1 0 13892 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1649_
timestamp 1644511149
transform 1 0 13340 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1650_
timestamp 1644511149
transform 1 0 13892 0 -1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1651_
timestamp 1644511149
transform 1 0 13708 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1652_
timestamp 1644511149
transform 1 0 14076 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1653_
timestamp 1644511149
transform 1 0 13156 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1654_
timestamp 1644511149
transform 1 0 22448 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1655_
timestamp 1644511149
transform 1 0 17940 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1656_
timestamp 1644511149
transform 1 0 15364 0 -1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1657_
timestamp 1644511149
transform 1 0 15272 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1658_
timestamp 1644511149
transform 1 0 18400 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1659_
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1660_
timestamp 1644511149
transform 1 0 18216 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1661_
timestamp 1644511149
transform 1 0 17204 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1662_
timestamp 1644511149
transform 1 0 15732 0 1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1663_
timestamp 1644511149
transform 1 0 15548 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1664_
timestamp 1644511149
transform 1 0 16744 0 1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1665_
timestamp 1644511149
transform 1 0 15916 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1666_
timestamp 1644511149
transform 1 0 16652 0 -1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1667_
timestamp 1644511149
transform 1 0 16836 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1668_
timestamp 1644511149
transform 1 0 15916 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1669_
timestamp 1644511149
transform 1 0 15824 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1670_
timestamp 1644511149
transform 1 0 19228 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1671_
timestamp 1644511149
transform 1 0 16928 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1672_
timestamp 1644511149
transform 1 0 14904 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1673_
timestamp 1644511149
transform 1 0 19228 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1674_
timestamp 1644511149
transform 1 0 19872 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1675_
timestamp 1644511149
transform 1 0 18584 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1676_
timestamp 1644511149
transform 1 0 18308 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1677_
timestamp 1644511149
transform 1 0 19228 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1678_
timestamp 1644511149
transform 1 0 17296 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1679_
timestamp 1644511149
transform 1 0 19136 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1680_
timestamp 1644511149
transform 1 0 20424 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1681_
timestamp 1644511149
transform 1 0 17940 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1682_
timestamp 1644511149
transform 1 0 19044 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1683_
timestamp 1644511149
transform 1 0 19228 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1684_
timestamp 1644511149
transform 1 0 19228 0 1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1685_
timestamp 1644511149
transform 1 0 20884 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1686_
timestamp 1644511149
transform 1 0 18492 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1687_
timestamp 1644511149
transform 1 0 20424 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1688_
timestamp 1644511149
transform 1 0 19872 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1689_
timestamp 1644511149
transform 1 0 20516 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1690_
timestamp 1644511149
transform 1 0 19964 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1691_
timestamp 1644511149
transform 1 0 21804 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1692_
timestamp 1644511149
transform 1 0 19872 0 1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1693_
timestamp 1644511149
transform 1 0 20516 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1694_
timestamp 1644511149
transform 1 0 19872 0 -1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1695_
timestamp 1644511149
transform 1 0 21068 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1696_
timestamp 1644511149
transform 1 0 19320 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1697_
timestamp 1644511149
transform 1 0 19780 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1698_
timestamp 1644511149
transform 1 0 20332 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1699_
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1700_
timestamp 1644511149
transform 1 0 20608 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1701_
timestamp 1644511149
transform 1 0 19504 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1702_
timestamp 1644511149
transform 1 0 19688 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1703_
timestamp 1644511149
transform 1 0 19412 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1704_
timestamp 1644511149
transform 1 0 19780 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1705_
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1706_
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1707_
timestamp 1644511149
transform 1 0 20424 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1708_
timestamp 1644511149
transform 1 0 19320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1709_
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1710_
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1711_
timestamp 1644511149
transform 1 0 19320 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1712_
timestamp 1644511149
transform 1 0 19872 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1713_
timestamp 1644511149
transform 1 0 21068 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1714_
timestamp 1644511149
transform 1 0 19412 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1715_
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1716_
timestamp 1644511149
transform 1 0 22540 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1717_
timestamp 1644511149
transform 1 0 22264 0 1 51136
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1718_
timestamp 1644511149
transform 1 0 25944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1719_
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1720_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1721_
timestamp 1644511149
transform 1 0 25116 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1722_
timestamp 1644511149
transform 1 0 24104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1724_
timestamp 1644511149
transform 1 0 22632 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1725_
timestamp 1644511149
transform 1 0 25852 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1726_
timestamp 1644511149
transform 1 0 25024 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1727_
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1728_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1729_
timestamp 1644511149
transform 1 0 22724 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1730_
timestamp 1644511149
transform 1 0 23828 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1731_
timestamp 1644511149
transform 1 0 22632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1732_
timestamp 1644511149
transform 1 0 23736 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1733_
timestamp 1644511149
transform 1 0 22724 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1734_
timestamp 1644511149
transform 1 0 25300 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1735_
timestamp 1644511149
transform 1 0 23368 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1736_
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1737_
timestamp 1644511149
transform 1 0 22448 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1738_
timestamp 1644511149
transform 1 0 24748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1739_
timestamp 1644511149
transform 1 0 24564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1740_
timestamp 1644511149
transform 1 0 23828 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1741_
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1742_
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _1743_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1744_
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1745_
timestamp 1644511149
transform 1 0 25392 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1746_
timestamp 1644511149
transform 1 0 24104 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1747_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1748_
timestamp 1644511149
transform 1 0 23644 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1749_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1750_
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1751_
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1752_
timestamp 1644511149
transform 1 0 23184 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1753_
timestamp 1644511149
transform 1 0 25300 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1754_
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1755_
timestamp 1644511149
transform 1 0 25208 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1756_
timestamp 1644511149
transform 1 0 25208 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1757_
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1758_
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _1759_
timestamp 1644511149
transform 1 0 19872 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1760_
timestamp 1644511149
transform 1 0 20240 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1761_
timestamp 1644511149
transform 1 0 20424 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1762_
timestamp 1644511149
transform 1 0 22448 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1763_
timestamp 1644511149
transform 1 0 19780 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1764_
timestamp 1644511149
transform 1 0 20608 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1765_
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1766_
timestamp 1644511149
transform 1 0 18124 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1767_
timestamp 1644511149
transform 1 0 19320 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1768_
timestamp 1644511149
transform 1 0 20516 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1769_
timestamp 1644511149
transform 1 0 15732 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1770_
timestamp 1644511149
transform 1 0 15824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1771_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1772_
timestamp 1644511149
transform 1 0 20240 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1773_
timestamp 1644511149
transform 1 0 17940 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1774_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1775_
timestamp 1644511149
transform 1 0 18400 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1776_
timestamp 1644511149
transform 1 0 17848 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1777_
timestamp 1644511149
transform 1 0 17756 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1778_
timestamp 1644511149
transform 1 0 19964 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1779_
timestamp 1644511149
transform 1 0 20424 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1780_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1781_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1782_
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1783_
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1784_
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1785_
timestamp 1644511149
transform 1 0 15088 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1786_
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1787_
timestamp 1644511149
transform 1 0 15364 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1788_
timestamp 1644511149
transform 1 0 15364 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1789_
timestamp 1644511149
transform 1 0 14904 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1790_
timestamp 1644511149
transform 1 0 14996 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1791_
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1792_
timestamp 1644511149
transform 1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1793_
timestamp 1644511149
transform 1 0 14076 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1794_
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1795_
timestamp 1644511149
transform 1 0 14720 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1796_
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1797_
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1798_
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1799_
timestamp 1644511149
transform 1 0 13156 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1800_
timestamp 1644511149
transform 1 0 12696 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1801_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1802_
timestamp 1644511149
transform 1 0 12420 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1803_
timestamp 1644511149
transform 1 0 12328 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1804_
timestamp 1644511149
transform 1 0 12512 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1805_
timestamp 1644511149
transform 1 0 13248 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1806_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1807_
timestamp 1644511149
transform 1 0 12144 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1808_
timestamp 1644511149
transform 1 0 11592 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1809_
timestamp 1644511149
transform 1 0 11592 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1810_
timestamp 1644511149
transform 1 0 12236 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1811_
timestamp 1644511149
transform 1 0 10580 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1812_
timestamp 1644511149
transform 1 0 11500 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1813_
timestamp 1644511149
transform 1 0 11500 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1814_
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1815_
timestamp 1644511149
transform 1 0 10304 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1816_
timestamp 1644511149
transform 1 0 11040 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1817_
timestamp 1644511149
transform 1 0 10212 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1818_
timestamp 1644511149
transform 1 0 10672 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1819_
timestamp 1644511149
transform 1 0 12144 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1820_
timestamp 1644511149
transform 1 0 10396 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1821_
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1822_
timestamp 1644511149
transform 1 0 11960 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1823_
timestamp 1644511149
transform 1 0 12972 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1824_
timestamp 1644511149
transform 1 0 10764 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1825_
timestamp 1644511149
transform 1 0 9476 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1826_
timestamp 1644511149
transform 1 0 11868 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1827_
timestamp 1644511149
transform 1 0 10212 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1828_
timestamp 1644511149
transform 1 0 11500 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1829_
timestamp 1644511149
transform 1 0 10304 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1830_
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1831_
timestamp 1644511149
transform 1 0 11500 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1832_
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1833_
timestamp 1644511149
transform 1 0 11776 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1834_
timestamp 1644511149
transform 1 0 11684 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1835_
timestamp 1644511149
transform 1 0 15180 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1836_
timestamp 1644511149
transform 1 0 15640 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1837_
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1838_
timestamp 1644511149
transform 1 0 12328 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1839_
timestamp 1644511149
transform 1 0 13340 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1840_
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1841_
timestamp 1644511149
transform 1 0 14536 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1842_
timestamp 1644511149
transform 1 0 12788 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1843_
timestamp 1644511149
transform 1 0 13984 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1844_
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1845_
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1846_
timestamp 1644511149
transform 1 0 14076 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1847_
timestamp 1644511149
transform 1 0 15180 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1848_
timestamp 1644511149
transform 1 0 15088 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1849_
timestamp 1644511149
transform 1 0 14628 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1850_
timestamp 1644511149
transform 1 0 15364 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1851_
timestamp 1644511149
transform 1 0 15456 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1852_
timestamp 1644511149
transform 1 0 15364 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1853_
timestamp 1644511149
transform 1 0 15548 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1854_
timestamp 1644511149
transform 1 0 15272 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1855_
timestamp 1644511149
transform 1 0 14444 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1856_
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1857_
timestamp 1644511149
transform 1 0 18308 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1858_
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1859_
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1860_
timestamp 1644511149
transform 1 0 18952 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1861_
timestamp 1644511149
transform 1 0 16376 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1862_
timestamp 1644511149
transform 1 0 17848 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _1863_
timestamp 1644511149
transform 1 0 16100 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1864_
timestamp 1644511149
transform 1 0 17020 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1865_
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1866_
timestamp 1644511149
transform 1 0 18584 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1867_
timestamp 1644511149
transform 1 0 16468 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1868_
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1869_
timestamp 1644511149
transform 1 0 16744 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1870_
timestamp 1644511149
transform 1 0 17296 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1871_
timestamp 1644511149
transform 1 0 17480 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1872_
timestamp 1644511149
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1873_
timestamp 1644511149
transform 1 0 16744 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1874_
timestamp 1644511149
transform 1 0 16652 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1875_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1876_
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1877_
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1878_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1644511149
transform 1 0 21804 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1644511149
transform 1 0 19688 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1882_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 -1 59840
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1644511149
transform 1 0 19228 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1644511149
transform 1 0 17020 0 -1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1644511149
transform 1 0 18492 0 -1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1644511149
transform 1 0 17296 0 1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1887_
timestamp 1644511149
transform 1 0 16652 0 -1 54400
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1888_
timestamp 1644511149
transform 1 0 16928 0 -1 60928
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1889_
timestamp 1644511149
transform 1 0 14628 0 -1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1890_
timestamp 1644511149
transform 1 0 14444 0 -1 60928
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1644511149
transform 1 0 14076 0 1 56576
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1644511149
transform 1 0 13708 0 -1 66368
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1644511149
transform 1 0 13892 0 -1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1644511149
transform 1 0 15272 0 1 66368
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1895_
timestamp 1644511149
transform 1 0 14720 0 1 69632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1896_
timestamp 1644511149
transform 1 0 17020 0 -1 66368
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1897_
timestamp 1644511149
transform 1 0 17112 0 1 75072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1898_
timestamp 1644511149
transform 1 0 15180 0 1 75072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1644511149
transform 1 0 16836 0 -1 70720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1644511149
transform 1 0 18124 0 -1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1644511149
transform 1 0 18216 0 -1 75072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1644511149
transform 1 0 21804 0 -1 75072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1903_
timestamp 1644511149
transform 1 0 19780 0 1 75072
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1644511149
transform 1 0 20424 0 1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1905_
timestamp 1644511149
transform 1 0 21160 0 1 73984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1644511149
transform 1 0 22264 0 1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1644511149
transform 1 0 21344 0 1 65280
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1644511149
transform 1 0 21804 0 -1 65280
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1644511149
transform 1 0 21068 0 1 62016
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1644511149
transform 1 0 20976 0 1 59840
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1644511149
transform 1 0 20332 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1644511149
transform 1 0 19780 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1644511149
transform 1 0 19504 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1644511149
transform 1 0 19596 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1644511149
transform 1 0 21896 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1644511149
transform 1 0 22356 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1644511149
transform 1 0 21528 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1644511149
transform 1 0 21528 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1644511149
transform 1 0 21804 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1923_
timestamp 1644511149
transform 1 0 21988 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1644511149
transform 1 0 21896 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1927_
timestamp 1644511149
transform 1 0 23276 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1928_
timestamp 1644511149
transform 1 0 22448 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1929_
timestamp 1644511149
transform 1 0 22448 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1930_
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1931_
timestamp 1644511149
transform 1 0 23920 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1932_
timestamp 1644511149
transform 1 0 25024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1933_
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1934_
timestamp 1644511149
transform 1 0 20884 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1935_
timestamp 1644511149
transform 1 0 21896 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1936_
timestamp 1644511149
transform 1 0 20884 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1937_
timestamp 1644511149
transform 1 0 22080 0 -1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1938_
timestamp 1644511149
transform 1 0 19412 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1939_
timestamp 1644511149
transform 1 0 18400 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1940_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1941_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1942_
timestamp 1644511149
transform 1 0 17572 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1943_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1944_
timestamp 1644511149
transform 1 0 15640 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1945_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1946_
timestamp 1644511149
transform 1 0 15088 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1947_
timestamp 1644511149
transform 1 0 14996 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1948_
timestamp 1644511149
transform 1 0 14168 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1949_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1950_
timestamp 1644511149
transform 1 0 13892 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1951_
timestamp 1644511149
transform 1 0 12052 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1952_
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1953_
timestamp 1644511149
transform 1 0 14076 0 -1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1954_
timestamp 1644511149
transform 1 0 11592 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1955_
timestamp 1644511149
transform 1 0 11592 0 1 39168
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1956_
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1957_
timestamp 1644511149
transform 1 0 9660 0 1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1958_
timestamp 1644511149
transform 1 0 9660 0 1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1959_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 1 42432
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1960_
timestamp 1644511149
transform 1 0 9936 0 1 48960
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1961_
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1962_
timestamp 1644511149
transform 1 0 11776 0 1 52224
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1963_
timestamp 1644511149
transform 1 0 11776 0 1 50048
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1964_
timestamp 1644511149
transform 1 0 12788 0 -1 43520
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1965_
timestamp 1644511149
transform 1 0 12972 0 -1 50048
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1966_
timestamp 1644511149
transform 1 0 12604 0 -1 52224
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1967_
timestamp 1644511149
transform 1 0 14720 0 1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1968_
timestamp 1644511149
transform 1 0 13892 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1969_
timestamp 1644511149
transform 1 0 15548 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1970_
timestamp 1644511149
transform 1 0 14720 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1971_
timestamp 1644511149
transform 1 0 14628 0 1 46784
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1972_
timestamp 1644511149
transform 1 0 17112 0 1 47872
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1973_
timestamp 1644511149
transform 1 0 17296 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1974_
timestamp 1644511149
transform 1 0 17388 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1975_
timestamp 1644511149
transform 1 0 17296 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1976_
timestamp 1644511149
transform 1 0 16468 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1977_
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1978_
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1979_
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1980_
timestamp 1644511149
transform 1 0 16836 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1981_
timestamp 1644511149
transform 1 0 17940 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0047_
timestamp 1644511149
transform 1 0 19504 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0053_
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0426_
timestamp 1644511149
transform 1 0 16928 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0427_
timestamp 1644511149
transform 1 0 18860 0 -1 52224
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0428_
timestamp 1644511149
transform 1 0 16560 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0434_
timestamp 1644511149
transform 1 0 17020 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0435_
timestamp 1644511149
transform 1 0 16928 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0437_
timestamp 1644511149
transform 1 0 17020 0 -1 57664
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0443_
timestamp 1644511149
transform 1 0 15456 0 1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0445_
timestamp 1644511149
transform 1 0 15088 0 1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0451_
timestamp 1644511149
transform 1 0 19596 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0452_
timestamp 1644511149
transform 1 0 16652 0 1 69632
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0454_
timestamp 1644511149
transform 1 0 16928 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0455_
timestamp 1644511149
transform 1 0 18860 0 -1 56576
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0456_
timestamp 1644511149
transform 1 0 16928 0 1 70720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0462_
timestamp 1644511149
transform 1 0 18676 0 -1 70720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0464_
timestamp 1644511149
transform 1 0 19596 0 1 70720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0470_
timestamp 1644511149
transform 1 0 19964 0 1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0472_
timestamp 1644511149
transform 1 0 19504 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0478_
timestamp 1644511149
transform 1 0 19964 0 1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0480_
timestamp 1644511149
transform 1 0 19504 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0486_
timestamp 1644511149
transform 1 0 19504 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0488_
timestamp 1644511149
transform 1 0 20240 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0520_
timestamp 1644511149
transform 1 0 15272 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0521_
timestamp 1644511149
transform 1 0 18952 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0523_
timestamp 1644511149
transform 1 0 13984 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0524_
timestamp 1644511149
transform 1 0 18216 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0529_
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0531_
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0538_
timestamp 1644511149
transform 1 0 13892 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0540_
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0546_
timestamp 1644511149
transform 1 0 11776 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0548_
timestamp 1644511149
transform 1 0 11868 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0554_
timestamp 1644511149
transform 1 0 11684 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0556_
timestamp 1644511149
transform 1 0 11868 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0562_
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0564_
timestamp 1644511149
transform 1 0 14444 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0570_
timestamp 1644511149
transform 1 0 15732 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0572_
timestamp 1644511149
transform 1 0 17020 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0578_
timestamp 1644511149
transform 1 0 17020 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0580_
timestamp 1644511149
transform 1 0 16928 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_a_clk_i
timestamp 1644511149
transform 1 0 21988 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_b_clk_i
timestamp 1644511149
transform 1 0 20056 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0010_
timestamp 1644511149
transform 1 0 21804 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0047_
timestamp 1644511149
transform 1 0 22172 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0053_
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0426_
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0427_
timestamp 1644511149
transform 1 0 16836 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0428_
timestamp 1644511149
transform 1 0 13892 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0434_
timestamp 1644511149
transform 1 0 16744 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0435_
timestamp 1644511149
transform 1 0 17572 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0437_
timestamp 1644511149
transform 1 0 15824 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0443_
timestamp 1644511149
transform 1 0 15824 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0445_
timestamp 1644511149
transform 1 0 14536 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0451_
timestamp 1644511149
transform 1 0 19228 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0452_
timestamp 1644511149
transform 1 0 17296 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0454_
timestamp 1644511149
transform 1 0 15824 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0455_
timestamp 1644511149
transform 1 0 18952 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0456_
timestamp 1644511149
transform 1 0 17204 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0462_
timestamp 1644511149
transform 1 0 18308 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0464_
timestamp 1644511149
transform 1 0 19228 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0470_
timestamp 1644511149
transform 1 0 19136 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0472_
timestamp 1644511149
transform 1 0 19688 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0478_
timestamp 1644511149
transform 1 0 19964 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0480_
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0486_
timestamp 1644511149
transform 1 0 19044 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0488_
timestamp 1644511149
transform 1 0 20976 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0520_
timestamp 1644511149
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0521_
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0523_
timestamp 1644511149
transform 1 0 14444 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0524_
timestamp 1644511149
transform 1 0 19228 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0529_
timestamp 1644511149
transform 1 0 16008 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0531_
timestamp 1644511149
transform 1 0 16744 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0538_
timestamp 1644511149
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0540_
timestamp 1644511149
transform 1 0 13064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0546_
timestamp 1644511149
transform 1 0 9476 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0548_
timestamp 1644511149
transform 1 0 12236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0554_
timestamp 1644511149
transform 1 0 11868 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0556_
timestamp 1644511149
transform 1 0 12880 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0562_
timestamp 1644511149
transform 1 0 13248 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0564_
timestamp 1644511149
transform 1 0 13248 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0570_
timestamp 1644511149
transform 1 0 13248 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0572_
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0578_
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__0580_
timestamp 1644511149
transform 1 0 15824 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_a_clk_i
timestamp 1644511149
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_b_clk_i
timestamp 1644511149
transform 1 0 18400 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0010_
timestamp 1644511149
transform 1 0 23276 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0047_
timestamp 1644511149
transform 1 0 19780 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0053_
timestamp 1644511149
transform 1 0 19964 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0426_
timestamp 1644511149
transform 1 0 15824 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0427_
timestamp 1644511149
transform 1 0 21804 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0428_
timestamp 1644511149
transform 1 0 18216 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0434_
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0435_
timestamp 1644511149
transform 1 0 18308 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0437_
timestamp 1644511149
transform 1 0 17756 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0443_
timestamp 1644511149
transform 1 0 14720 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0445_
timestamp 1644511149
transform 1 0 15272 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0451_
timestamp 1644511149
transform 1 0 18768 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0452_
timestamp 1644511149
transform 1 0 17020 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0454_
timestamp 1644511149
transform 1 0 17940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0455_
timestamp 1644511149
transform 1 0 19596 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0456_
timestamp 1644511149
transform 1 0 15824 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0462_
timestamp 1644511149
transform 1 0 19596 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0464_
timestamp 1644511149
transform 1 0 18400 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0470_
timestamp 1644511149
transform 1 0 20056 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0472_
timestamp 1644511149
transform 1 0 21068 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0478_
timestamp 1644511149
transform 1 0 20608 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0480_
timestamp 1644511149
transform 1 0 20700 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0486_
timestamp 1644511149
transform 1 0 20516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0488_
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0520_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0521_
timestamp 1644511149
transform 1 0 19228 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0523_
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0524_
timestamp 1644511149
transform 1 0 19136 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0529_
timestamp 1644511149
transform 1 0 17388 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0531_
timestamp 1644511149
transform 1 0 16008 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0538_
timestamp 1644511149
transform 1 0 13064 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0540_
timestamp 1644511149
transform 1 0 13156 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0546_
timestamp 1644511149
transform 1 0 15180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0548_
timestamp 1644511149
transform 1 0 10304 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0554_
timestamp 1644511149
transform 1 0 10672 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0556_
timestamp 1644511149
transform 1 0 13064 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0562_
timestamp 1644511149
transform 1 0 13248 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0564_
timestamp 1644511149
transform 1 0 14444 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0570_
timestamp 1644511149
transform 1 0 17848 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0572_
timestamp 1644511149
transform 1 0 16008 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0578_
timestamp 1644511149
transform 1 0 17480 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__0580_
timestamp 1644511149
transform 1 0 15824 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_a_clk_i
timestamp 1644511149
transform 1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_b_clk_i
timestamp 1644511149
transform 1 0 22356 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold5
timestamp 1644511149
transform 1 0 17848 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold6
timestamp 1644511149
transform 1 0 21252 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold8
timestamp 1644511149
transform 1 0 20240 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold9
timestamp 1644511149
transform 1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1644511149
transform 1 0 22356 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1644511149
transform 1 0 22080 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 2024 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 2392 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 2024 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 3220 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 2392 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 1380 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 2024 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 1380 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 1380 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 1380 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 1380 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 1380 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 1380 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 1380 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 1380 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 1380 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1644511149
transform 1 0 1380 0 1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 1380 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 1380 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 1380 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 1380 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 1380 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 1380 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 1380 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 1380 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 2668 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1644511149
transform 1 0 1380 0 -1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 1380 0 1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1644511149
transform 1 0 1380 0 1 76160
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 1380 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1644511149
transform 1 0 2668 0 -1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform 1 0 3772 0 1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 1380 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1644511149
transform 1 0 1380 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 1380 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 1380 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform 1 0 1380 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 1380 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1644511149
transform 1 0 1380 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input65
timestamp 1644511149
transform 1 0 29624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 29808 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input67
timestamp 1644511149
transform 1 0 29624 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1644511149
transform 1 0 29900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1644511149
transform 1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 26772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1644511149
transform 1 0 29808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1644511149
transform 1 0 29808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1644511149
transform 1 0 29808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1644511149
transform 1 0 28704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1644511149
transform 1 0 28704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1644511149
transform 1 0 29808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1644511149
transform 1 0 29808 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1644511149
transform 1 0 29808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1644511149
transform 1 0 29900 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1644511149
transform 1 0 29808 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input85
timestamp 1644511149
transform 1 0 29808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1644511149
transform 1 0 29808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1644511149
transform 1 0 28704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1644511149
transform 1 0 29256 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1644511149
transform 1 0 29072 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1644511149
transform 1 0 28704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1644511149
transform 1 0 28060 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1644511149
transform 1 0 27416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1644511149
transform 1 0 29808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input94
timestamp 1644511149
transform 1 0 28704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1644511149
transform 1 0 29808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1644511149
transform 1 0 29072 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1644511149
transform 1 0 28428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1644511149
transform 1 0 29256 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input102
timestamp 1644511149
transform 1 0 28152 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input103
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1644511149
transform 1 0 28612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1644511149
transform 1 0 29256 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1644511149
transform 1 0 29808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1644511149
transform 1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1644511149
transform 1 0 27968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1644511149
transform 1 0 27968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input113
timestamp 1644511149
transform 1 0 28888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input114
timestamp 1644511149
transform 1 0 29624 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input115
timestamp 1644511149
transform 1 0 29624 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input116
timestamp 1644511149
transform 1 0 29624 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input117
timestamp 1644511149
transform 1 0 29624 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input118
timestamp 1644511149
transform 1 0 28520 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input119
timestamp 1644511149
transform 1 0 28704 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input120
timestamp 1644511149
transform 1 0 28888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input121
timestamp 1644511149
transform 1 0 28888 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input122
timestamp 1644511149
transform 1 0 27968 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1644511149
transform 1 0 28428 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input124
timestamp 1644511149
transform 1 0 29624 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input125
timestamp 1644511149
transform 1 0 29624 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input126
timestamp 1644511149
transform 1 0 29624 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input127
timestamp 1644511149
transform 1 0 29808 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input128
timestamp 1644511149
transform 1 0 28612 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input129
timestamp 1644511149
transform 1 0 29808 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input130
timestamp 1644511149
transform 1 0 28888 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input131
timestamp 1644511149
transform 1 0 29624 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input132
timestamp 1644511149
transform 1 0 29624 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input133
timestamp 1644511149
transform 1 0 29624 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input134
timestamp 1644511149
transform 1 0 28520 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input135
timestamp 1644511149
transform 1 0 29624 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input136
timestamp 1644511149
transform 1 0 28888 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input137
timestamp 1644511149
transform 1 0 26864 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input138
timestamp 1644511149
transform 1 0 28152 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input139
timestamp 1644511149
transform 1 0 29808 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input140
timestamp 1644511149
transform 1 0 29624 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input141
timestamp 1644511149
transform 1 0 28520 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input142
timestamp 1644511149
transform 1 0 26956 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input143
timestamp 1644511149
transform 1 0 27324 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input144
timestamp 1644511149
transform 1 0 26772 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input145
timestamp 1644511149
transform 1 0 29808 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input146
timestamp 1644511149
transform 1 0 29624 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input147
timestamp 1644511149
transform 1 0 29808 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input148
timestamp 1644511149
transform 1 0 28612 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input149
timestamp 1644511149
transform 1 0 29624 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input150
timestamp 1644511149
transform 1 0 28704 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input151
timestamp 1644511149
transform 1 0 28704 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input152
timestamp 1644511149
transform 1 0 27968 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1644511149
transform 1 0 25760 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input154
timestamp 1644511149
transform 1 0 29624 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input155
timestamp 1644511149
transform 1 0 28520 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1644511149
transform 1 0 29808 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input157
timestamp 1644511149
transform 1 0 29808 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input158
timestamp 1644511149
transform 1 0 28704 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input159
timestamp 1644511149
transform 1 0 29072 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1644511149
transform 1 0 27784 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1644511149
transform 1 0 29808 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input162
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net199_2
timestamp 1644511149
transform 1 0 17940 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net199_3
timestamp 1644511149
transform 1 0 20976 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net199_4
timestamp 1644511149
transform 1 0 23552 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 1380 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 1380 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 1380 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output179
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output180
timestamp 1644511149
transform 1 0 2024 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1644511149
transform 1 0 28704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1644511149
transform 1 0 29808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1644511149
transform 1 0 29808 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1644511149
transform 1 0 29808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1644511149
transform 1 0 29808 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1644511149
transform 1 0 29808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1644511149
transform 1 0 28704 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1644511149
transform 1 0 29808 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1644511149
transform 1 0 29072 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1644511149
transform 1 0 28704 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1644511149
transform 1 0 29808 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1644511149
transform 1 0 28704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1644511149
transform 1 0 28704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1644511149
transform 1 0 27968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1644511149
transform 1 0 29808 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1644511149
transform 1 0 29808 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1644511149
transform 1 0 29808 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1644511149
transform 1 0 29072 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1644511149
transform 1 0 29808 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1644511149
transform 1 0 28336 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1644511149
transform 1 0 28704 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1644511149
transform 1 0 27968 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1644511149
transform 1 0 28704 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1644511149
transform 1 0 26128 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1644511149
transform 1 0 25116 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1644511149
transform 1 0 29808 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1644511149
transform 1 0 28428 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1644511149
transform 1 0 27508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1644511149
transform 1 0 28704 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1644511149
transform 1 0 26864 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1644511149
transform 1 0 27508 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1644511149
transform 1 0 29072 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1644511149
transform 1 0 29808 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1644511149
transform 1 0 29808 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1644511149
transform 1 0 29808 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1644511149
transform 1 0 29808 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1644511149
transform 1 0 29808 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1644511149
transform 1 0 29808 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1644511149
transform 1 0 29808 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1644511149
transform 1 0 29808 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1644511149
transform 1 0 29808 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1644511149
transform 1 0 29808 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1644511149
transform 1 0 29808 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1644511149
transform 1 0 27876 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1644511149
transform 1 0 29808 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1644511149
transform 1 0 29808 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1644511149
transform 1 0 29808 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1644511149
transform 1 0 29072 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1644511149
transform 1 0 29808 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1644511149
transform 1 0 29808 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1644511149
transform 1 0 28704 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1644511149
transform 1 0 29072 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1644511149
transform 1 0 27968 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1644511149
transform 1 0 28336 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1644511149
transform 1 0 29808 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1644511149
transform 1 0 28704 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1644511149
transform 1 0 27232 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1644511149
transform 1 0 29072 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output280
timestamp 1644511149
transform 1 0 29808 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1644511149
transform 1 0 28704 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1644511149
transform 1 0 29808 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output283
timestamp 1644511149
transform 1 0 29808 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output284
timestamp 1644511149
transform 1 0 28704 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1644511149
transform 1 0 29072 0 -1 69632
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 4904 800 5024 6 ram_addr0[0]
port 0 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 ram_addr0[1]
port 1 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 ram_addr0[2]
port 2 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 ram_addr0[3]
port 3 nsew signal tristate
rlabel metal3 s 0 7488 800 7608 6 ram_addr0[4]
port 4 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 ram_addr0[5]
port 5 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 ram_addr0[6]
port 6 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 ram_addr0[7]
port 7 nsew signal tristate
rlabel metal3 s 0 53728 800 53848 6 ram_addr1[0]
port 8 nsew signal tristate
rlabel metal3 s 0 54408 800 54528 6 ram_addr1[1]
port 9 nsew signal tristate
rlabel metal3 s 0 55088 800 55208 6 ram_addr1[2]
port 10 nsew signal tristate
rlabel metal3 s 0 55768 800 55888 6 ram_addr1[3]
port 11 nsew signal tristate
rlabel metal3 s 0 56448 800 56568 6 ram_addr1[4]
port 12 nsew signal tristate
rlabel metal3 s 0 56992 800 57112 6 ram_addr1[5]
port 13 nsew signal tristate
rlabel metal3 s 0 57672 800 57792 6 ram_addr1[6]
port 14 nsew signal tristate
rlabel metal3 s 0 58352 800 58472 6 ram_addr1[7]
port 15 nsew signal tristate
rlabel metal3 s 0 280 800 400 6 ram_clk0
port 16 nsew signal tristate
rlabel metal3 s 0 52368 800 52488 6 ram_clk1
port 17 nsew signal tristate
rlabel metal3 s 0 824 800 944 6 ram_csb0
port 18 nsew signal tristate
rlabel metal3 s 0 53048 800 53168 6 ram_csb1
port 19 nsew signal tristate
rlabel metal3 s 0 10072 800 10192 6 ram_din0[0]
port 20 nsew signal tristate
rlabel metal3 s 0 16736 800 16856 6 ram_din0[10]
port 21 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 ram_din0[11]
port 22 nsew signal tristate
rlabel metal3 s 0 18096 800 18216 6 ram_din0[12]
port 23 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 ram_din0[13]
port 24 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 ram_din0[14]
port 25 nsew signal tristate
rlabel metal3 s 0 20000 800 20120 6 ram_din0[15]
port 26 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 ram_din0[16]
port 27 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 ram_din0[17]
port 28 nsew signal tristate
rlabel metal3 s 0 22040 800 22160 6 ram_din0[18]
port 29 nsew signal tristate
rlabel metal3 s 0 22720 800 22840 6 ram_din0[19]
port 30 nsew signal tristate
rlabel metal3 s 0 10752 800 10872 6 ram_din0[1]
port 31 nsew signal tristate
rlabel metal3 s 0 23400 800 23520 6 ram_din0[20]
port 32 nsew signal tristate
rlabel metal3 s 0 23944 800 24064 6 ram_din0[21]
port 33 nsew signal tristate
rlabel metal3 s 0 24624 800 24744 6 ram_din0[22]
port 34 nsew signal tristate
rlabel metal3 s 0 25304 800 25424 6 ram_din0[23]
port 35 nsew signal tristate
rlabel metal3 s 0 25984 800 26104 6 ram_din0[24]
port 36 nsew signal tristate
rlabel metal3 s 0 26664 800 26784 6 ram_din0[25]
port 37 nsew signal tristate
rlabel metal3 s 0 27344 800 27464 6 ram_din0[26]
port 38 nsew signal tristate
rlabel metal3 s 0 28024 800 28144 6 ram_din0[27]
port 39 nsew signal tristate
rlabel metal3 s 0 28568 800 28688 6 ram_din0[28]
port 40 nsew signal tristate
rlabel metal3 s 0 29248 800 29368 6 ram_din0[29]
port 41 nsew signal tristate
rlabel metal3 s 0 11432 800 11552 6 ram_din0[2]
port 42 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 ram_din0[30]
port 43 nsew signal tristate
rlabel metal3 s 0 30608 800 30728 6 ram_din0[31]
port 44 nsew signal tristate
rlabel metal3 s 0 12112 800 12232 6 ram_din0[3]
port 45 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 ram_din0[4]
port 46 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 ram_din0[5]
port 47 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 ram_din0[6]
port 48 nsew signal tristate
rlabel metal3 s 0 14696 800 14816 6 ram_din0[7]
port 49 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 ram_din0[8]
port 50 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 ram_din0[9]
port 51 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 ram_dout0[0]
port 52 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 ram_dout0[10]
port 53 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 ram_dout0[11]
port 54 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 ram_dout0[12]
port 55 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 ram_dout0[13]
port 56 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 ram_dout0[14]
port 57 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 ram_dout0[15]
port 58 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 ram_dout0[16]
port 59 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 ram_dout0[17]
port 60 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 ram_dout0[18]
port 61 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 ram_dout0[19]
port 62 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 ram_dout0[1]
port 63 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 ram_dout0[20]
port 64 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 ram_dout0[21]
port 65 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 ram_dout0[22]
port 66 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 ram_dout0[23]
port 67 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 ram_dout0[24]
port 68 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 ram_dout0[25]
port 69 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 ram_dout0[26]
port 70 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 ram_dout0[27]
port 71 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 ram_dout0[28]
port 72 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 ram_dout0[29]
port 73 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 ram_dout0[2]
port 74 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 ram_dout0[30]
port 75 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 ram_dout0[31]
port 76 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 ram_dout0[3]
port 77 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 ram_dout0[4]
port 78 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 ram_dout0[5]
port 79 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 ram_dout0[6]
port 80 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 ram_dout0[7]
port 81 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 ram_dout0[8]
port 82 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 ram_dout0[9]
port 83 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 ram_dout1[0]
port 84 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 ram_dout1[10]
port 85 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 ram_dout1[11]
port 86 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 ram_dout1[12]
port 87 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 ram_dout1[13]
port 88 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 ram_dout1[14]
port 89 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 ram_dout1[15]
port 90 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 ram_dout1[16]
port 91 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 ram_dout1[17]
port 92 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 ram_dout1[18]
port 93 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 ram_dout1[19]
port 94 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 ram_dout1[1]
port 95 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 ram_dout1[20]
port 96 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 ram_dout1[21]
port 97 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 ram_dout1[22]
port 98 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 ram_dout1[23]
port 99 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 ram_dout1[24]
port 100 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 ram_dout1[25]
port 101 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 ram_dout1[26]
port 102 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 ram_dout1[27]
port 103 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 ram_dout1[28]
port 104 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 ram_dout1[29]
port 105 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 ram_dout1[2]
port 106 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 ram_dout1[30]
port 107 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 ram_dout1[31]
port 108 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 ram_dout1[3]
port 109 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 ram_dout1[4]
port 110 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 ram_dout1[5]
port 111 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 ram_dout1[6]
port 112 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 ram_dout1[7]
port 113 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 ram_dout1[8]
port 114 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 ram_dout1[9]
port 115 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 ram_web0
port 116 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 ram_wmask0[0]
port 117 nsew signal tristate
rlabel metal3 s 0 2864 800 2984 6 ram_wmask0[1]
port 118 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 ram_wmask0[2]
port 119 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 ram_wmask0[3]
port 120 nsew signal tristate
rlabel metal4 s 5910 2128 6230 77840 6 vccd1
port 121 nsew power input
rlabel metal4 s 15840 2128 16160 77840 6 vccd1
port 121 nsew power input
rlabel metal4 s 25771 2128 26091 77840 6 vccd1
port 121 nsew power input
rlabel metal4 s 10874 2128 11194 77840 6 vssd1
port 122 nsew ground input
rlabel metal4 s 20805 2128 21125 77840 6 vssd1
port 122 nsew ground input
rlabel metal3 s 31200 552 32000 672 6 wb_a_clk_i
port 123 nsew signal input
rlabel metal3 s 31200 960 32000 1080 6 wb_a_rst_i
port 124 nsew signal input
rlabel metal3 s 31200 40536 32000 40656 6 wb_b_clk_i
port 125 nsew signal input
rlabel metal3 s 31200 40944 32000 41064 6 wb_b_rst_i
port 126 nsew signal input
rlabel metal3 s 31200 2864 32000 2984 6 wbs_a_ack_o
port 127 nsew signal tristate
rlabel metal3 s 31200 5312 32000 5432 6 wbs_a_adr_i[0]
port 128 nsew signal input
rlabel metal3 s 31200 9936 32000 10056 6 wbs_a_adr_i[10]
port 129 nsew signal input
rlabel metal3 s 31200 5720 32000 5840 6 wbs_a_adr_i[1]
port 130 nsew signal input
rlabel metal3 s 31200 6128 32000 6248 6 wbs_a_adr_i[2]
port 131 nsew signal input
rlabel metal3 s 31200 6672 32000 6792 6 wbs_a_adr_i[3]
port 132 nsew signal input
rlabel metal3 s 31200 7080 32000 7200 6 wbs_a_adr_i[4]
port 133 nsew signal input
rlabel metal3 s 31200 7624 32000 7744 6 wbs_a_adr_i[5]
port 134 nsew signal input
rlabel metal3 s 31200 8032 32000 8152 6 wbs_a_adr_i[6]
port 135 nsew signal input
rlabel metal3 s 31200 8576 32000 8696 6 wbs_a_adr_i[7]
port 136 nsew signal input
rlabel metal3 s 31200 8984 32000 9104 6 wbs_a_adr_i[8]
port 137 nsew signal input
rlabel metal3 s 31200 9528 32000 9648 6 wbs_a_adr_i[9]
port 138 nsew signal input
rlabel metal3 s 31200 1912 32000 2032 6 wbs_a_cyc_i
port 139 nsew signal input
rlabel metal3 s 31200 10480 32000 10600 6 wbs_a_dat_i[0]
port 140 nsew signal input
rlabel metal3 s 31200 15104 32000 15224 6 wbs_a_dat_i[10]
port 141 nsew signal input
rlabel metal3 s 31200 15648 32000 15768 6 wbs_a_dat_i[11]
port 142 nsew signal input
rlabel metal3 s 31200 16056 32000 16176 6 wbs_a_dat_i[12]
port 143 nsew signal input
rlabel metal3 s 31200 16600 32000 16720 6 wbs_a_dat_i[13]
port 144 nsew signal input
rlabel metal3 s 31200 17008 32000 17128 6 wbs_a_dat_i[14]
port 145 nsew signal input
rlabel metal3 s 31200 17416 32000 17536 6 wbs_a_dat_i[15]
port 146 nsew signal input
rlabel metal3 s 31200 17960 32000 18080 6 wbs_a_dat_i[16]
port 147 nsew signal input
rlabel metal3 s 31200 18368 32000 18488 6 wbs_a_dat_i[17]
port 148 nsew signal input
rlabel metal3 s 31200 18912 32000 19032 6 wbs_a_dat_i[18]
port 149 nsew signal input
rlabel metal3 s 31200 19320 32000 19440 6 wbs_a_dat_i[19]
port 150 nsew signal input
rlabel metal3 s 31200 10888 32000 11008 6 wbs_a_dat_i[1]
port 151 nsew signal input
rlabel metal3 s 31200 19864 32000 19984 6 wbs_a_dat_i[20]
port 152 nsew signal input
rlabel metal3 s 31200 20272 32000 20392 6 wbs_a_dat_i[21]
port 153 nsew signal input
rlabel metal3 s 31200 20816 32000 20936 6 wbs_a_dat_i[22]
port 154 nsew signal input
rlabel metal3 s 31200 21224 32000 21344 6 wbs_a_dat_i[23]
port 155 nsew signal input
rlabel metal3 s 31200 21768 32000 21888 6 wbs_a_dat_i[24]
port 156 nsew signal input
rlabel metal3 s 31200 22176 32000 22296 6 wbs_a_dat_i[25]
port 157 nsew signal input
rlabel metal3 s 31200 22720 32000 22840 6 wbs_a_dat_i[26]
port 158 nsew signal input
rlabel metal3 s 31200 23128 32000 23248 6 wbs_a_dat_i[27]
port 159 nsew signal input
rlabel metal3 s 31200 23536 32000 23656 6 wbs_a_dat_i[28]
port 160 nsew signal input
rlabel metal3 s 31200 24080 32000 24200 6 wbs_a_dat_i[29]
port 161 nsew signal input
rlabel metal3 s 31200 11432 32000 11552 6 wbs_a_dat_i[2]
port 162 nsew signal input
rlabel metal3 s 31200 24488 32000 24608 6 wbs_a_dat_i[30]
port 163 nsew signal input
rlabel metal3 s 31200 25032 32000 25152 6 wbs_a_dat_i[31]
port 164 nsew signal input
rlabel metal3 s 31200 11840 32000 11960 6 wbs_a_dat_i[3]
port 165 nsew signal input
rlabel metal3 s 31200 12248 32000 12368 6 wbs_a_dat_i[4]
port 166 nsew signal input
rlabel metal3 s 31200 12792 32000 12912 6 wbs_a_dat_i[5]
port 167 nsew signal input
rlabel metal3 s 31200 13200 32000 13320 6 wbs_a_dat_i[6]
port 168 nsew signal input
rlabel metal3 s 31200 13744 32000 13864 6 wbs_a_dat_i[7]
port 169 nsew signal input
rlabel metal3 s 31200 14152 32000 14272 6 wbs_a_dat_i[8]
port 170 nsew signal input
rlabel metal3 s 31200 14696 32000 14816 6 wbs_a_dat_i[9]
port 171 nsew signal input
rlabel metal3 s 31200 25440 32000 25560 6 wbs_a_dat_o[0]
port 172 nsew signal tristate
rlabel metal3 s 31200 30200 32000 30320 6 wbs_a_dat_o[10]
port 173 nsew signal tristate
rlabel metal3 s 31200 30608 32000 30728 6 wbs_a_dat_o[11]
port 174 nsew signal tristate
rlabel metal3 s 31200 31152 32000 31272 6 wbs_a_dat_o[12]
port 175 nsew signal tristate
rlabel metal3 s 31200 31560 32000 31680 6 wbs_a_dat_o[13]
port 176 nsew signal tristate
rlabel metal3 s 31200 32104 32000 32224 6 wbs_a_dat_o[14]
port 177 nsew signal tristate
rlabel metal3 s 31200 32512 32000 32632 6 wbs_a_dat_o[15]
port 178 nsew signal tristate
rlabel metal3 s 31200 33056 32000 33176 6 wbs_a_dat_o[16]
port 179 nsew signal tristate
rlabel metal3 s 31200 33464 32000 33584 6 wbs_a_dat_o[17]
port 180 nsew signal tristate
rlabel metal3 s 31200 34008 32000 34128 6 wbs_a_dat_o[18]
port 181 nsew signal tristate
rlabel metal3 s 31200 34416 32000 34536 6 wbs_a_dat_o[19]
port 182 nsew signal tristate
rlabel metal3 s 31200 25984 32000 26104 6 wbs_a_dat_o[1]
port 183 nsew signal tristate
rlabel metal3 s 31200 34824 32000 34944 6 wbs_a_dat_o[20]
port 184 nsew signal tristate
rlabel metal3 s 31200 35368 32000 35488 6 wbs_a_dat_o[21]
port 185 nsew signal tristate
rlabel metal3 s 31200 35776 32000 35896 6 wbs_a_dat_o[22]
port 186 nsew signal tristate
rlabel metal3 s 31200 36320 32000 36440 6 wbs_a_dat_o[23]
port 187 nsew signal tristate
rlabel metal3 s 31200 36728 32000 36848 6 wbs_a_dat_o[24]
port 188 nsew signal tristate
rlabel metal3 s 31200 37272 32000 37392 6 wbs_a_dat_o[25]
port 189 nsew signal tristate
rlabel metal3 s 31200 37680 32000 37800 6 wbs_a_dat_o[26]
port 190 nsew signal tristate
rlabel metal3 s 31200 38224 32000 38344 6 wbs_a_dat_o[27]
port 191 nsew signal tristate
rlabel metal3 s 31200 38632 32000 38752 6 wbs_a_dat_o[28]
port 192 nsew signal tristate
rlabel metal3 s 31200 39176 32000 39296 6 wbs_a_dat_o[29]
port 193 nsew signal tristate
rlabel metal3 s 31200 26392 32000 26512 6 wbs_a_dat_o[2]
port 194 nsew signal tristate
rlabel metal3 s 31200 39584 32000 39704 6 wbs_a_dat_o[30]
port 195 nsew signal tristate
rlabel metal3 s 31200 40128 32000 40248 6 wbs_a_dat_o[31]
port 196 nsew signal tristate
rlabel metal3 s 31200 26936 32000 27056 6 wbs_a_dat_o[3]
port 197 nsew signal tristate
rlabel metal3 s 31200 27344 32000 27464 6 wbs_a_dat_o[4]
port 198 nsew signal tristate
rlabel metal3 s 31200 27888 32000 28008 6 wbs_a_dat_o[5]
port 199 nsew signal tristate
rlabel metal3 s 31200 28296 32000 28416 6 wbs_a_dat_o[6]
port 200 nsew signal tristate
rlabel metal3 s 31200 28704 32000 28824 6 wbs_a_dat_o[7]
port 201 nsew signal tristate
rlabel metal3 s 31200 29248 32000 29368 6 wbs_a_dat_o[8]
port 202 nsew signal tristate
rlabel metal3 s 31200 29656 32000 29776 6 wbs_a_dat_o[9]
port 203 nsew signal tristate
rlabel metal3 s 31200 3408 32000 3528 6 wbs_a_sel_i[0]
port 204 nsew signal input
rlabel metal3 s 31200 3816 32000 3936 6 wbs_a_sel_i[1]
port 205 nsew signal input
rlabel metal3 s 31200 4360 32000 4480 6 wbs_a_sel_i[2]
port 206 nsew signal input
rlabel metal3 s 31200 4768 32000 4888 6 wbs_a_sel_i[3]
port 207 nsew signal input
rlabel metal3 s 31200 1504 32000 1624 6 wbs_a_stb_i
port 208 nsew signal input
rlabel metal3 s 31200 2456 32000 2576 6 wbs_a_we_i
port 209 nsew signal input
rlabel metal3 s 31200 42848 32000 42968 6 wbs_b_ack_o
port 210 nsew signal tristate
rlabel metal3 s 31200 45296 32000 45416 6 wbs_b_adr_i[0]
port 211 nsew signal input
rlabel metal3 s 31200 45704 32000 45824 6 wbs_b_adr_i[1]
port 212 nsew signal input
rlabel metal3 s 31200 46112 32000 46232 6 wbs_b_adr_i[2]
port 213 nsew signal input
rlabel metal3 s 31200 46656 32000 46776 6 wbs_b_adr_i[3]
port 214 nsew signal input
rlabel metal3 s 31200 47064 32000 47184 6 wbs_b_adr_i[4]
port 215 nsew signal input
rlabel metal3 s 31200 47608 32000 47728 6 wbs_b_adr_i[5]
port 216 nsew signal input
rlabel metal3 s 31200 48016 32000 48136 6 wbs_b_adr_i[6]
port 217 nsew signal input
rlabel metal3 s 31200 48560 32000 48680 6 wbs_b_adr_i[7]
port 218 nsew signal input
rlabel metal3 s 31200 48968 32000 49088 6 wbs_b_adr_i[8]
port 219 nsew signal input
rlabel metal3 s 31200 49512 32000 49632 6 wbs_b_adr_i[9]
port 220 nsew signal input
rlabel metal3 s 31200 41896 32000 42016 6 wbs_b_cyc_i
port 221 nsew signal input
rlabel metal3 s 31200 49920 32000 50040 6 wbs_b_dat_i[0]
port 222 nsew signal input
rlabel metal3 s 31200 54680 32000 54800 6 wbs_b_dat_i[10]
port 223 nsew signal input
rlabel metal3 s 31200 55088 32000 55208 6 wbs_b_dat_i[11]
port 224 nsew signal input
rlabel metal3 s 31200 55632 32000 55752 6 wbs_b_dat_i[12]
port 225 nsew signal input
rlabel metal3 s 31200 56040 32000 56160 6 wbs_b_dat_i[13]
port 226 nsew signal input
rlabel metal3 s 31200 56584 32000 56704 6 wbs_b_dat_i[14]
port 227 nsew signal input
rlabel metal3 s 31200 56992 32000 57112 6 wbs_b_dat_i[15]
port 228 nsew signal input
rlabel metal3 s 31200 57400 32000 57520 6 wbs_b_dat_i[16]
port 229 nsew signal input
rlabel metal3 s 31200 57944 32000 58064 6 wbs_b_dat_i[17]
port 230 nsew signal input
rlabel metal3 s 31200 58352 32000 58472 6 wbs_b_dat_i[18]
port 231 nsew signal input
rlabel metal3 s 31200 58896 32000 59016 6 wbs_b_dat_i[19]
port 232 nsew signal input
rlabel metal3 s 31200 50464 32000 50584 6 wbs_b_dat_i[1]
port 233 nsew signal input
rlabel metal3 s 31200 59304 32000 59424 6 wbs_b_dat_i[20]
port 234 nsew signal input
rlabel metal3 s 31200 59848 32000 59968 6 wbs_b_dat_i[21]
port 235 nsew signal input
rlabel metal3 s 31200 60256 32000 60376 6 wbs_b_dat_i[22]
port 236 nsew signal input
rlabel metal3 s 31200 60800 32000 60920 6 wbs_b_dat_i[23]
port 237 nsew signal input
rlabel metal3 s 31200 61208 32000 61328 6 wbs_b_dat_i[24]
port 238 nsew signal input
rlabel metal3 s 31200 61752 32000 61872 6 wbs_b_dat_i[25]
port 239 nsew signal input
rlabel metal3 s 31200 62160 32000 62280 6 wbs_b_dat_i[26]
port 240 nsew signal input
rlabel metal3 s 31200 62704 32000 62824 6 wbs_b_dat_i[27]
port 241 nsew signal input
rlabel metal3 s 31200 63112 32000 63232 6 wbs_b_dat_i[28]
port 242 nsew signal input
rlabel metal3 s 31200 63520 32000 63640 6 wbs_b_dat_i[29]
port 243 nsew signal input
rlabel metal3 s 31200 50872 32000 50992 6 wbs_b_dat_i[2]
port 244 nsew signal input
rlabel metal3 s 31200 64064 32000 64184 6 wbs_b_dat_i[30]
port 245 nsew signal input
rlabel metal3 s 31200 64472 32000 64592 6 wbs_b_dat_i[31]
port 246 nsew signal input
rlabel metal3 s 31200 51416 32000 51536 6 wbs_b_dat_i[3]
port 247 nsew signal input
rlabel metal3 s 31200 51824 32000 51944 6 wbs_b_dat_i[4]
port 248 nsew signal input
rlabel metal3 s 31200 52232 32000 52352 6 wbs_b_dat_i[5]
port 249 nsew signal input
rlabel metal3 s 31200 52776 32000 52896 6 wbs_b_dat_i[6]
port 250 nsew signal input
rlabel metal3 s 31200 53184 32000 53304 6 wbs_b_dat_i[7]
port 251 nsew signal input
rlabel metal3 s 31200 53728 32000 53848 6 wbs_b_dat_i[8]
port 252 nsew signal input
rlabel metal3 s 31200 54136 32000 54256 6 wbs_b_dat_i[9]
port 253 nsew signal input
rlabel metal3 s 31200 65016 32000 65136 6 wbs_b_dat_o[0]
port 254 nsew signal tristate
rlabel metal3 s 31200 69640 32000 69760 6 wbs_b_dat_o[10]
port 255 nsew signal tristate
rlabel metal3 s 31200 70184 32000 70304 6 wbs_b_dat_o[11]
port 256 nsew signal tristate
rlabel metal3 s 31200 70592 32000 70712 6 wbs_b_dat_o[12]
port 257 nsew signal tristate
rlabel metal3 s 31200 71136 32000 71256 6 wbs_b_dat_o[13]
port 258 nsew signal tristate
rlabel metal3 s 31200 71544 32000 71664 6 wbs_b_dat_o[14]
port 259 nsew signal tristate
rlabel metal3 s 31200 72088 32000 72208 6 wbs_b_dat_o[15]
port 260 nsew signal tristate
rlabel metal3 s 31200 72496 32000 72616 6 wbs_b_dat_o[16]
port 261 nsew signal tristate
rlabel metal3 s 31200 73040 32000 73160 6 wbs_b_dat_o[17]
port 262 nsew signal tristate
rlabel metal3 s 31200 73448 32000 73568 6 wbs_b_dat_o[18]
port 263 nsew signal tristate
rlabel metal3 s 31200 73992 32000 74112 6 wbs_b_dat_o[19]
port 264 nsew signal tristate
rlabel metal3 s 31200 65424 32000 65544 6 wbs_b_dat_o[1]
port 265 nsew signal tristate
rlabel metal3 s 31200 74400 32000 74520 6 wbs_b_dat_o[20]
port 266 nsew signal tristate
rlabel metal3 s 31200 74808 32000 74928 6 wbs_b_dat_o[21]
port 267 nsew signal tristate
rlabel metal3 s 31200 75352 32000 75472 6 wbs_b_dat_o[22]
port 268 nsew signal tristate
rlabel metal3 s 31200 75760 32000 75880 6 wbs_b_dat_o[23]
port 269 nsew signal tristate
rlabel metal3 s 31200 76304 32000 76424 6 wbs_b_dat_o[24]
port 270 nsew signal tristate
rlabel metal3 s 31200 76712 32000 76832 6 wbs_b_dat_o[25]
port 271 nsew signal tristate
rlabel metal3 s 31200 77256 32000 77376 6 wbs_b_dat_o[26]
port 272 nsew signal tristate
rlabel metal3 s 31200 77664 32000 77784 6 wbs_b_dat_o[27]
port 273 nsew signal tristate
rlabel metal3 s 31200 78208 32000 78328 6 wbs_b_dat_o[28]
port 274 nsew signal tristate
rlabel metal3 s 31200 78616 32000 78736 6 wbs_b_dat_o[29]
port 275 nsew signal tristate
rlabel metal3 s 31200 65968 32000 66088 6 wbs_b_dat_o[2]
port 276 nsew signal tristate
rlabel metal3 s 31200 79160 32000 79280 6 wbs_b_dat_o[30]
port 277 nsew signal tristate
rlabel metal3 s 31200 79568 32000 79688 6 wbs_b_dat_o[31]
port 278 nsew signal tristate
rlabel metal3 s 31200 66376 32000 66496 6 wbs_b_dat_o[3]
port 279 nsew signal tristate
rlabel metal3 s 31200 66920 32000 67040 6 wbs_b_dat_o[4]
port 280 nsew signal tristate
rlabel metal3 s 31200 67328 32000 67448 6 wbs_b_dat_o[5]
port 281 nsew signal tristate
rlabel metal3 s 31200 67872 32000 67992 6 wbs_b_dat_o[6]
port 282 nsew signal tristate
rlabel metal3 s 31200 68280 32000 68400 6 wbs_b_dat_o[7]
port 283 nsew signal tristate
rlabel metal3 s 31200 68688 32000 68808 6 wbs_b_dat_o[8]
port 284 nsew signal tristate
rlabel metal3 s 31200 69232 32000 69352 6 wbs_b_dat_o[9]
port 285 nsew signal tristate
rlabel metal3 s 31200 43392 32000 43512 6 wbs_b_sel_i[0]
port 286 nsew signal input
rlabel metal3 s 31200 43800 32000 43920 6 wbs_b_sel_i[1]
port 287 nsew signal input
rlabel metal3 s 31200 44344 32000 44464 6 wbs_b_sel_i[2]
port 288 nsew signal input
rlabel metal3 s 31200 44752 32000 44872 6 wbs_b_sel_i[3]
port 289 nsew signal input
rlabel metal3 s 31200 41488 32000 41608 6 wbs_b_stb_i
port 290 nsew signal input
rlabel metal3 s 31200 42440 32000 42560 6 wbs_b_we_i
port 291 nsew signal input
rlabel metal3 s 31200 144 32000 264 6 writable_port_req
port 292 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32000 80000
<< end >>
