VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_openram_wrapper
  CLASS BLOCK ;
  FOREIGN wb_openram_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 300.000 ;
  PIN ram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END ram_addr0[0]
  PIN ram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END ram_addr0[1]
  PIN ram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END ram_addr0[2]
  PIN ram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END ram_addr0[3]
  PIN ram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END ram_addr0[4]
  PIN ram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END ram_addr0[5]
  PIN ram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END ram_addr0[6]
  PIN ram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END ram_addr0[7]
  PIN ram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END ram_clk0
  PIN ram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END ram_csb0
  PIN ram_din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END ram_din0[0]
  PIN ram_din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END ram_din0[10]
  PIN ram_din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END ram_din0[11]
  PIN ram_din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END ram_din0[12]
  PIN ram_din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END ram_din0[13]
  PIN ram_din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END ram_din0[14]
  PIN ram_din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END ram_din0[15]
  PIN ram_din0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END ram_din0[16]
  PIN ram_din0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END ram_din0[17]
  PIN ram_din0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END ram_din0[18]
  PIN ram_din0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END ram_din0[19]
  PIN ram_din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END ram_din0[1]
  PIN ram_din0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END ram_din0[20]
  PIN ram_din0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END ram_din0[21]
  PIN ram_din0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END ram_din0[22]
  PIN ram_din0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END ram_din0[23]
  PIN ram_din0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END ram_din0[24]
  PIN ram_din0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END ram_din0[25]
  PIN ram_din0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END ram_din0[26]
  PIN ram_din0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END ram_din0[27]
  PIN ram_din0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END ram_din0[28]
  PIN ram_din0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END ram_din0[29]
  PIN ram_din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END ram_din0[2]
  PIN ram_din0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END ram_din0[30]
  PIN ram_din0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END ram_din0[31]
  PIN ram_din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END ram_din0[3]
  PIN ram_din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END ram_din0[4]
  PIN ram_din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END ram_din0[5]
  PIN ram_din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END ram_din0[6]
  PIN ram_din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END ram_din0[7]
  PIN ram_din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END ram_din0[8]
  PIN ram_din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END ram_din0[9]
  PIN ram_dout0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END ram_dout0[0]
  PIN ram_dout0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END ram_dout0[10]
  PIN ram_dout0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END ram_dout0[11]
  PIN ram_dout0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END ram_dout0[12]
  PIN ram_dout0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END ram_dout0[13]
  PIN ram_dout0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END ram_dout0[14]
  PIN ram_dout0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END ram_dout0[15]
  PIN ram_dout0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END ram_dout0[16]
  PIN ram_dout0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END ram_dout0[17]
  PIN ram_dout0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END ram_dout0[18]
  PIN ram_dout0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END ram_dout0[19]
  PIN ram_dout0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END ram_dout0[1]
  PIN ram_dout0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END ram_dout0[20]
  PIN ram_dout0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END ram_dout0[21]
  PIN ram_dout0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END ram_dout0[22]
  PIN ram_dout0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END ram_dout0[23]
  PIN ram_dout0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END ram_dout0[24]
  PIN ram_dout0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END ram_dout0[25]
  PIN ram_dout0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END ram_dout0[26]
  PIN ram_dout0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END ram_dout0[27]
  PIN ram_dout0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END ram_dout0[28]
  PIN ram_dout0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END ram_dout0[29]
  PIN ram_dout0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END ram_dout0[2]
  PIN ram_dout0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END ram_dout0[30]
  PIN ram_dout0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END ram_dout0[31]
  PIN ram_dout0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END ram_dout0[3]
  PIN ram_dout0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END ram_dout0[4]
  PIN ram_dout0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END ram_dout0[5]
  PIN ram_dout0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END ram_dout0[6]
  PIN ram_dout0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END ram_dout0[7]
  PIN ram_dout0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END ram_dout0[8]
  PIN ram_dout0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END ram_dout0[9]
  PIN ram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END ram_web0
  PIN ram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END ram_wmask0[0]
  PIN ram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END ram_wmask0[1]
  PIN ram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END ram_wmask0[2]
  PIN ram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END ram_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.545 10.640 11.145 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.195 10.640 20.795 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.850 10.640 30.450 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.370 10.640 15.970 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.025 10.640 25.625 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 1.400 40.000 2.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 4.120 40.000 4.720 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 15.000 40.000 15.600 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 29.280 40.000 29.880 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 57.840 40.000 58.440 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 60.560 40.000 61.160 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 63.280 40.000 63.880 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 66.000 40.000 66.600 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 68.720 40.000 69.320 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 72.120 40.000 72.720 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 74.840 40.000 75.440 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 77.560 40.000 78.160 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 80.280 40.000 80.880 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 83.000 40.000 83.600 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 32.000 40.000 32.600 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 85.720 40.000 86.320 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 88.440 40.000 89.040 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 91.840 40.000 92.440 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 94.560 40.000 95.160 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 97.280 40.000 97.880 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 100.000 40.000 100.600 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 102.720 40.000 103.320 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 105.440 40.000 106.040 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 108.840 40.000 109.440 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 111.560 40.000 112.160 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 34.720 40.000 35.320 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 114.280 40.000 114.880 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 117.000 40.000 117.600 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 38.120 40.000 38.720 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 40.840 40.000 41.440 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 43.560 40.000 44.160 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 46.280 40.000 46.880 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 49.000 40.000 49.600 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 51.720 40.000 52.320 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 55.120 40.000 55.720 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 9.560 40.000 10.160 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 119.720 40.000 120.320 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 148.280 40.000 148.880 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 151.000 40.000 151.600 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 153.720 40.000 154.320 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 156.440 40.000 157.040 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 159.160 40.000 159.760 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 162.560 40.000 163.160 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 165.280 40.000 165.880 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 168.000 40.000 168.600 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 170.720 40.000 171.320 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 173.440 40.000 174.040 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 122.440 40.000 123.040 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 176.160 40.000 176.760 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 179.560 40.000 180.160 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 182.280 40.000 182.880 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 185.000 40.000 185.600 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 187.720 40.000 188.320 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 190.440 40.000 191.040 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 193.160 40.000 193.760 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 196.560 40.000 197.160 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 199.280 40.000 199.880 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 202.000 40.000 202.600 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 125.840 40.000 126.440 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 204.720 40.000 205.320 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 207.440 40.000 208.040 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 128.560 40.000 129.160 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 131.280 40.000 131.880 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 134.000 40.000 134.600 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 136.720 40.000 137.320 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 139.440 40.000 140.040 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 142.840 40.000 143.440 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 145.560 40.000 146.160 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 210.160 40.000 210.760 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 238.720 40.000 239.320 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 241.440 40.000 242.040 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 244.160 40.000 244.760 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 246.880 40.000 247.480 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 250.280 40.000 250.880 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 253.000 40.000 253.600 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 255.720 40.000 256.320 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 258.440 40.000 259.040 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 261.160 40.000 261.760 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 263.880 40.000 264.480 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 213.560 40.000 214.160 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 267.280 40.000 267.880 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 270.000 40.000 270.600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 272.720 40.000 273.320 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 275.440 40.000 276.040 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 278.160 40.000 278.760 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 280.880 40.000 281.480 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 284.280 40.000 284.880 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 287.000 40.000 287.600 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 289.720 40.000 290.320 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 292.440 40.000 293.040 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 216.280 40.000 216.880 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 295.160 40.000 295.760 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 297.880 40.000 298.480 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 219.000 40.000 219.600 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 221.720 40.000 222.320 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 224.440 40.000 225.040 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 227.160 40.000 227.760 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 229.880 40.000 230.480 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 233.280 40.000 233.880 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 236.000 40.000 236.600 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 17.720 40.000 18.320 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 21.120 40.000 21.720 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 23.840 40.000 24.440 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 26.560 40.000 27.160 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 6.840 40.000 7.440 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 12.280 40.000 12.880 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 4.745 10.795 39.875 288.405 ;
      LAYER met1 ;
        RECT 4.685 10.640 39.935 288.560 ;
      LAYER met2 ;
        RECT 5.620 1.515 39.460 298.365 ;
      LAYER met3 ;
        RECT 4.000 298.200 35.600 298.345 ;
        RECT 4.400 297.480 35.600 298.200 ;
        RECT 4.400 296.800 36.000 297.480 ;
        RECT 4.000 296.160 36.000 296.800 ;
        RECT 4.000 294.760 35.600 296.160 ;
        RECT 4.000 294.120 36.000 294.760 ;
        RECT 4.400 293.440 36.000 294.120 ;
        RECT 4.400 292.720 35.600 293.440 ;
        RECT 4.000 292.040 35.600 292.720 ;
        RECT 4.000 290.720 36.000 292.040 ;
        RECT 4.400 289.320 35.600 290.720 ;
        RECT 4.000 288.000 36.000 289.320 ;
        RECT 4.000 286.640 35.600 288.000 ;
        RECT 4.400 286.600 35.600 286.640 ;
        RECT 4.400 285.280 36.000 286.600 ;
        RECT 4.400 285.240 35.600 285.280 ;
        RECT 4.000 283.880 35.600 285.240 ;
        RECT 4.000 283.240 36.000 283.880 ;
        RECT 4.400 281.880 36.000 283.240 ;
        RECT 4.400 281.840 35.600 281.880 ;
        RECT 4.000 280.480 35.600 281.840 ;
        RECT 4.000 279.160 36.000 280.480 ;
        RECT 4.400 277.760 35.600 279.160 ;
        RECT 4.000 276.440 36.000 277.760 ;
        RECT 4.000 275.080 35.600 276.440 ;
        RECT 4.400 275.040 35.600 275.080 ;
        RECT 4.400 273.720 36.000 275.040 ;
        RECT 4.400 273.680 35.600 273.720 ;
        RECT 4.000 272.320 35.600 273.680 ;
        RECT 4.000 271.680 36.000 272.320 ;
        RECT 4.400 271.000 36.000 271.680 ;
        RECT 4.400 270.280 35.600 271.000 ;
        RECT 4.000 269.600 35.600 270.280 ;
        RECT 4.000 268.280 36.000 269.600 ;
        RECT 4.000 267.600 35.600 268.280 ;
        RECT 4.400 266.880 35.600 267.600 ;
        RECT 4.400 266.200 36.000 266.880 ;
        RECT 4.000 264.880 36.000 266.200 ;
        RECT 4.000 264.200 35.600 264.880 ;
        RECT 4.400 263.480 35.600 264.200 ;
        RECT 4.400 262.800 36.000 263.480 ;
        RECT 4.000 262.160 36.000 262.800 ;
        RECT 4.000 260.760 35.600 262.160 ;
        RECT 4.000 260.120 36.000 260.760 ;
        RECT 4.400 259.440 36.000 260.120 ;
        RECT 4.400 258.720 35.600 259.440 ;
        RECT 4.000 258.040 35.600 258.720 ;
        RECT 4.000 256.720 36.000 258.040 ;
        RECT 4.400 255.320 35.600 256.720 ;
        RECT 4.000 254.000 36.000 255.320 ;
        RECT 4.000 252.640 35.600 254.000 ;
        RECT 4.400 252.600 35.600 252.640 ;
        RECT 4.400 251.280 36.000 252.600 ;
        RECT 4.400 251.240 35.600 251.280 ;
        RECT 4.000 249.880 35.600 251.240 ;
        RECT 4.000 248.560 36.000 249.880 ;
        RECT 4.400 247.880 36.000 248.560 ;
        RECT 4.400 247.160 35.600 247.880 ;
        RECT 4.000 246.480 35.600 247.160 ;
        RECT 4.000 245.160 36.000 246.480 ;
        RECT 4.400 243.760 35.600 245.160 ;
        RECT 4.000 242.440 36.000 243.760 ;
        RECT 4.000 241.080 35.600 242.440 ;
        RECT 4.400 241.040 35.600 241.080 ;
        RECT 4.400 239.720 36.000 241.040 ;
        RECT 4.400 239.680 35.600 239.720 ;
        RECT 4.000 238.320 35.600 239.680 ;
        RECT 4.000 237.680 36.000 238.320 ;
        RECT 4.400 237.000 36.000 237.680 ;
        RECT 4.400 236.280 35.600 237.000 ;
        RECT 4.000 235.600 35.600 236.280 ;
        RECT 4.000 234.280 36.000 235.600 ;
        RECT 4.000 233.600 35.600 234.280 ;
        RECT 4.400 232.880 35.600 233.600 ;
        RECT 4.400 232.200 36.000 232.880 ;
        RECT 4.000 230.880 36.000 232.200 ;
        RECT 4.000 229.520 35.600 230.880 ;
        RECT 4.400 229.480 35.600 229.520 ;
        RECT 4.400 228.160 36.000 229.480 ;
        RECT 4.400 228.120 35.600 228.160 ;
        RECT 4.000 226.760 35.600 228.120 ;
        RECT 4.000 226.120 36.000 226.760 ;
        RECT 4.400 225.440 36.000 226.120 ;
        RECT 4.400 224.720 35.600 225.440 ;
        RECT 4.000 224.040 35.600 224.720 ;
        RECT 4.000 222.720 36.000 224.040 ;
        RECT 4.000 222.040 35.600 222.720 ;
        RECT 4.400 221.320 35.600 222.040 ;
        RECT 4.400 220.640 36.000 221.320 ;
        RECT 4.000 220.000 36.000 220.640 ;
        RECT 4.000 218.640 35.600 220.000 ;
        RECT 4.400 218.600 35.600 218.640 ;
        RECT 4.400 217.280 36.000 218.600 ;
        RECT 4.400 217.240 35.600 217.280 ;
        RECT 4.000 215.880 35.600 217.240 ;
        RECT 4.000 214.560 36.000 215.880 ;
        RECT 4.400 213.160 35.600 214.560 ;
        RECT 4.000 211.160 36.000 213.160 ;
        RECT 4.400 209.760 35.600 211.160 ;
        RECT 4.000 208.440 36.000 209.760 ;
        RECT 4.000 207.080 35.600 208.440 ;
        RECT 4.400 207.040 35.600 207.080 ;
        RECT 4.400 205.720 36.000 207.040 ;
        RECT 4.400 205.680 35.600 205.720 ;
        RECT 4.000 204.320 35.600 205.680 ;
        RECT 4.000 203.000 36.000 204.320 ;
        RECT 4.400 201.600 35.600 203.000 ;
        RECT 4.000 200.280 36.000 201.600 ;
        RECT 4.000 199.600 35.600 200.280 ;
        RECT 4.400 198.880 35.600 199.600 ;
        RECT 4.400 198.200 36.000 198.880 ;
        RECT 4.000 197.560 36.000 198.200 ;
        RECT 4.000 196.160 35.600 197.560 ;
        RECT 4.000 195.520 36.000 196.160 ;
        RECT 4.400 194.160 36.000 195.520 ;
        RECT 4.400 194.120 35.600 194.160 ;
        RECT 4.000 192.760 35.600 194.120 ;
        RECT 4.000 192.120 36.000 192.760 ;
        RECT 4.400 191.440 36.000 192.120 ;
        RECT 4.400 190.720 35.600 191.440 ;
        RECT 4.000 190.040 35.600 190.720 ;
        RECT 4.000 188.720 36.000 190.040 ;
        RECT 4.000 188.040 35.600 188.720 ;
        RECT 4.400 187.320 35.600 188.040 ;
        RECT 4.400 186.640 36.000 187.320 ;
        RECT 4.000 186.000 36.000 186.640 ;
        RECT 4.000 184.600 35.600 186.000 ;
        RECT 4.000 183.960 36.000 184.600 ;
        RECT 4.400 183.280 36.000 183.960 ;
        RECT 4.400 182.560 35.600 183.280 ;
        RECT 4.000 181.880 35.600 182.560 ;
        RECT 4.000 180.560 36.000 181.880 ;
        RECT 4.400 179.160 35.600 180.560 ;
        RECT 4.000 177.160 36.000 179.160 ;
        RECT 4.000 176.480 35.600 177.160 ;
        RECT 4.400 175.760 35.600 176.480 ;
        RECT 4.400 175.080 36.000 175.760 ;
        RECT 4.000 174.440 36.000 175.080 ;
        RECT 4.000 173.080 35.600 174.440 ;
        RECT 4.400 173.040 35.600 173.080 ;
        RECT 4.400 171.720 36.000 173.040 ;
        RECT 4.400 171.680 35.600 171.720 ;
        RECT 4.000 170.320 35.600 171.680 ;
        RECT 4.000 169.000 36.000 170.320 ;
        RECT 4.400 167.600 35.600 169.000 ;
        RECT 4.000 166.280 36.000 167.600 ;
        RECT 4.000 165.600 35.600 166.280 ;
        RECT 4.400 164.880 35.600 165.600 ;
        RECT 4.400 164.200 36.000 164.880 ;
        RECT 4.000 163.560 36.000 164.200 ;
        RECT 4.000 162.160 35.600 163.560 ;
        RECT 4.000 161.520 36.000 162.160 ;
        RECT 4.400 160.160 36.000 161.520 ;
        RECT 4.400 160.120 35.600 160.160 ;
        RECT 4.000 158.760 35.600 160.120 ;
        RECT 4.000 157.440 36.000 158.760 ;
        RECT 4.400 156.040 35.600 157.440 ;
        RECT 4.000 154.720 36.000 156.040 ;
        RECT 4.000 154.040 35.600 154.720 ;
        RECT 4.400 153.320 35.600 154.040 ;
        RECT 4.400 152.640 36.000 153.320 ;
        RECT 4.000 152.000 36.000 152.640 ;
        RECT 4.000 150.600 35.600 152.000 ;
        RECT 4.000 149.960 36.000 150.600 ;
        RECT 4.400 149.280 36.000 149.960 ;
        RECT 4.400 148.560 35.600 149.280 ;
        RECT 4.000 147.880 35.600 148.560 ;
        RECT 4.000 146.560 36.000 147.880 ;
        RECT 4.400 145.160 35.600 146.560 ;
        RECT 4.000 143.840 36.000 145.160 ;
        RECT 4.000 142.480 35.600 143.840 ;
        RECT 4.400 142.440 35.600 142.480 ;
        RECT 4.400 141.080 36.000 142.440 ;
        RECT 4.000 140.440 36.000 141.080 ;
        RECT 4.000 139.040 35.600 140.440 ;
        RECT 4.000 138.400 36.000 139.040 ;
        RECT 4.400 137.720 36.000 138.400 ;
        RECT 4.400 137.000 35.600 137.720 ;
        RECT 4.000 136.320 35.600 137.000 ;
        RECT 4.000 135.000 36.000 136.320 ;
        RECT 4.400 133.600 35.600 135.000 ;
        RECT 4.000 132.280 36.000 133.600 ;
        RECT 4.000 130.920 35.600 132.280 ;
        RECT 4.400 130.880 35.600 130.920 ;
        RECT 4.400 129.560 36.000 130.880 ;
        RECT 4.400 129.520 35.600 129.560 ;
        RECT 4.000 128.160 35.600 129.520 ;
        RECT 4.000 127.520 36.000 128.160 ;
        RECT 4.400 126.840 36.000 127.520 ;
        RECT 4.400 126.120 35.600 126.840 ;
        RECT 4.000 125.440 35.600 126.120 ;
        RECT 4.000 123.440 36.000 125.440 ;
        RECT 4.400 122.040 35.600 123.440 ;
        RECT 4.000 120.720 36.000 122.040 ;
        RECT 4.000 120.040 35.600 120.720 ;
        RECT 4.400 119.320 35.600 120.040 ;
        RECT 4.400 118.640 36.000 119.320 ;
        RECT 4.000 118.000 36.000 118.640 ;
        RECT 4.000 116.600 35.600 118.000 ;
        RECT 4.000 115.960 36.000 116.600 ;
        RECT 4.400 115.280 36.000 115.960 ;
        RECT 4.400 114.560 35.600 115.280 ;
        RECT 4.000 113.880 35.600 114.560 ;
        RECT 4.000 112.560 36.000 113.880 ;
        RECT 4.000 111.880 35.600 112.560 ;
        RECT 4.400 111.160 35.600 111.880 ;
        RECT 4.400 110.480 36.000 111.160 ;
        RECT 4.000 109.840 36.000 110.480 ;
        RECT 4.000 108.480 35.600 109.840 ;
        RECT 4.400 108.440 35.600 108.480 ;
        RECT 4.400 107.080 36.000 108.440 ;
        RECT 4.000 106.440 36.000 107.080 ;
        RECT 4.000 105.040 35.600 106.440 ;
        RECT 4.000 104.400 36.000 105.040 ;
        RECT 4.400 103.720 36.000 104.400 ;
        RECT 4.400 103.000 35.600 103.720 ;
        RECT 4.000 102.320 35.600 103.000 ;
        RECT 4.000 101.000 36.000 102.320 ;
        RECT 4.400 99.600 35.600 101.000 ;
        RECT 4.000 98.280 36.000 99.600 ;
        RECT 4.000 96.920 35.600 98.280 ;
        RECT 4.400 96.880 35.600 96.920 ;
        RECT 4.400 95.560 36.000 96.880 ;
        RECT 4.400 95.520 35.600 95.560 ;
        RECT 4.000 94.160 35.600 95.520 ;
        RECT 4.000 92.840 36.000 94.160 ;
        RECT 4.400 91.440 35.600 92.840 ;
        RECT 4.000 89.440 36.000 91.440 ;
        RECT 4.400 88.040 35.600 89.440 ;
        RECT 4.000 86.720 36.000 88.040 ;
        RECT 4.000 85.360 35.600 86.720 ;
        RECT 4.400 85.320 35.600 85.360 ;
        RECT 4.400 84.000 36.000 85.320 ;
        RECT 4.400 83.960 35.600 84.000 ;
        RECT 4.000 82.600 35.600 83.960 ;
        RECT 4.000 81.960 36.000 82.600 ;
        RECT 4.400 81.280 36.000 81.960 ;
        RECT 4.400 80.560 35.600 81.280 ;
        RECT 4.000 79.880 35.600 80.560 ;
        RECT 4.000 78.560 36.000 79.880 ;
        RECT 4.000 77.880 35.600 78.560 ;
        RECT 4.400 77.160 35.600 77.880 ;
        RECT 4.400 76.480 36.000 77.160 ;
        RECT 4.000 75.840 36.000 76.480 ;
        RECT 4.000 74.480 35.600 75.840 ;
        RECT 4.400 74.440 35.600 74.480 ;
        RECT 4.400 73.120 36.000 74.440 ;
        RECT 4.400 73.080 35.600 73.120 ;
        RECT 4.000 71.720 35.600 73.080 ;
        RECT 4.000 70.400 36.000 71.720 ;
        RECT 4.400 69.720 36.000 70.400 ;
        RECT 4.400 69.000 35.600 69.720 ;
        RECT 4.000 68.320 35.600 69.000 ;
        RECT 4.000 67.000 36.000 68.320 ;
        RECT 4.000 66.320 35.600 67.000 ;
        RECT 4.400 65.600 35.600 66.320 ;
        RECT 4.400 64.920 36.000 65.600 ;
        RECT 4.000 64.280 36.000 64.920 ;
        RECT 4.000 62.920 35.600 64.280 ;
        RECT 4.400 62.880 35.600 62.920 ;
        RECT 4.400 61.560 36.000 62.880 ;
        RECT 4.400 61.520 35.600 61.560 ;
        RECT 4.000 60.160 35.600 61.520 ;
        RECT 4.000 58.840 36.000 60.160 ;
        RECT 4.400 57.440 35.600 58.840 ;
        RECT 4.000 56.120 36.000 57.440 ;
        RECT 4.000 55.440 35.600 56.120 ;
        RECT 4.400 54.720 35.600 55.440 ;
        RECT 4.400 54.040 36.000 54.720 ;
        RECT 4.000 52.720 36.000 54.040 ;
        RECT 4.000 51.360 35.600 52.720 ;
        RECT 4.400 51.320 35.600 51.360 ;
        RECT 4.400 50.000 36.000 51.320 ;
        RECT 4.400 49.960 35.600 50.000 ;
        RECT 4.000 48.600 35.600 49.960 ;
        RECT 4.000 47.280 36.000 48.600 ;
        RECT 4.400 45.880 35.600 47.280 ;
        RECT 4.000 44.560 36.000 45.880 ;
        RECT 4.000 43.880 35.600 44.560 ;
        RECT 4.400 43.160 35.600 43.880 ;
        RECT 4.400 42.480 36.000 43.160 ;
        RECT 4.000 41.840 36.000 42.480 ;
        RECT 4.000 40.440 35.600 41.840 ;
        RECT 4.000 39.800 36.000 40.440 ;
        RECT 4.400 39.120 36.000 39.800 ;
        RECT 4.400 38.400 35.600 39.120 ;
        RECT 4.000 37.720 35.600 38.400 ;
        RECT 4.000 36.400 36.000 37.720 ;
        RECT 4.400 35.720 36.000 36.400 ;
        RECT 4.400 35.000 35.600 35.720 ;
        RECT 4.000 34.320 35.600 35.000 ;
        RECT 4.000 33.000 36.000 34.320 ;
        RECT 4.000 32.320 35.600 33.000 ;
        RECT 4.400 31.600 35.600 32.320 ;
        RECT 4.400 30.920 36.000 31.600 ;
        RECT 4.000 30.280 36.000 30.920 ;
        RECT 4.000 28.920 35.600 30.280 ;
        RECT 4.400 28.880 35.600 28.920 ;
        RECT 4.400 27.560 36.000 28.880 ;
        RECT 4.400 27.520 35.600 27.560 ;
        RECT 4.000 26.160 35.600 27.520 ;
        RECT 4.000 24.840 36.000 26.160 ;
        RECT 4.400 23.440 35.600 24.840 ;
        RECT 4.000 22.120 36.000 23.440 ;
        RECT 4.000 20.760 35.600 22.120 ;
        RECT 4.400 20.720 35.600 20.760 ;
        RECT 4.400 19.360 36.000 20.720 ;
        RECT 4.000 18.720 36.000 19.360 ;
        RECT 4.000 17.360 35.600 18.720 ;
        RECT 4.400 17.320 35.600 17.360 ;
        RECT 4.400 16.000 36.000 17.320 ;
        RECT 4.400 15.960 35.600 16.000 ;
        RECT 4.000 14.600 35.600 15.960 ;
        RECT 4.000 13.280 36.000 14.600 ;
        RECT 4.400 11.880 35.600 13.280 ;
        RECT 4.000 10.560 36.000 11.880 ;
        RECT 4.000 9.880 35.600 10.560 ;
        RECT 4.400 9.160 35.600 9.880 ;
        RECT 4.400 8.480 36.000 9.160 ;
        RECT 4.000 7.840 36.000 8.480 ;
        RECT 4.000 6.440 35.600 7.840 ;
        RECT 4.000 5.800 36.000 6.440 ;
        RECT 4.400 5.120 36.000 5.800 ;
        RECT 4.400 4.400 35.600 5.120 ;
        RECT 4.000 3.720 35.600 4.400 ;
        RECT 4.000 2.400 36.000 3.720 ;
        RECT 4.400 1.535 35.600 2.400 ;
      LAYER met4 ;
        RECT 12.255 10.640 13.970 288.560 ;
        RECT 16.370 10.640 18.795 288.560 ;
        RECT 21.195 10.640 23.625 288.560 ;
        RECT 26.025 10.640 28.225 288.560 ;
  END
END wb_openram_wrapper
END LIBRARY

