magic
tech sky130A
magscale 1 2
timestamp 1647558826
<< obsli1 >>
rect 1104 2159 30820 77809
<< obsm1 >>
rect 1104 1300 31984 77840
<< obsm2 >>
rect 1306 167 31984 79665
<< metal3 >>
rect 0 79568 800 79688
rect 31200 79568 32000 79688
rect 31200 79160 32000 79280
rect 0 78888 800 79008
rect 31200 78616 32000 78736
rect 0 78208 800 78328
rect 31200 78208 32000 78328
rect 0 77528 800 77648
rect 31200 77664 32000 77784
rect 31200 77256 32000 77376
rect 0 76848 800 76968
rect 31200 76712 32000 76832
rect 0 76168 800 76288
rect 31200 76304 32000 76424
rect 31200 75760 32000 75880
rect 0 75488 800 75608
rect 31200 75352 32000 75472
rect 0 74944 800 75064
rect 31200 74808 32000 74928
rect 0 74264 800 74384
rect 31200 74400 32000 74520
rect 31200 73992 32000 74112
rect 0 73584 800 73704
rect 31200 73448 32000 73568
rect 0 72904 800 73024
rect 31200 73040 32000 73160
rect 31200 72496 32000 72616
rect 0 72224 800 72344
rect 31200 72088 32000 72208
rect 0 71544 800 71664
rect 31200 71544 32000 71664
rect 31200 71136 32000 71256
rect 0 70864 800 70984
rect 31200 70592 32000 70712
rect 0 70320 800 70440
rect 31200 70184 32000 70304
rect 0 69640 800 69760
rect 31200 69640 32000 69760
rect 31200 69232 32000 69352
rect 0 68960 800 69080
rect 31200 68688 32000 68808
rect 0 68280 800 68400
rect 31200 68280 32000 68400
rect 31200 67872 32000 67992
rect 0 67600 800 67720
rect 31200 67328 32000 67448
rect 0 66920 800 67040
rect 31200 66920 32000 67040
rect 0 66240 800 66360
rect 31200 66376 32000 66496
rect 31200 65968 32000 66088
rect 0 65696 800 65816
rect 31200 65424 32000 65544
rect 0 65016 800 65136
rect 31200 65016 32000 65136
rect 0 64336 800 64456
rect 31200 64472 32000 64592
rect 31200 64064 32000 64184
rect 0 63656 800 63776
rect 31200 63520 32000 63640
rect 0 62976 800 63096
rect 31200 63112 32000 63232
rect 31200 62704 32000 62824
rect 0 62296 800 62416
rect 31200 62160 32000 62280
rect 0 61616 800 61736
rect 31200 61752 32000 61872
rect 0 61072 800 61192
rect 31200 61208 32000 61328
rect 31200 60800 32000 60920
rect 0 60392 800 60512
rect 31200 60256 32000 60376
rect 0 59712 800 59832
rect 31200 59848 32000 59968
rect 31200 59304 32000 59424
rect 0 59032 800 59152
rect 31200 58896 32000 59016
rect 0 58352 800 58472
rect 31200 58352 32000 58472
rect 31200 57944 32000 58064
rect 0 57672 800 57792
rect 31200 57400 32000 57520
rect 0 56992 800 57112
rect 31200 56992 32000 57112
rect 0 56448 800 56568
rect 31200 56584 32000 56704
rect 31200 56040 32000 56160
rect 0 55768 800 55888
rect 31200 55632 32000 55752
rect 0 55088 800 55208
rect 31200 55088 32000 55208
rect 31200 54680 32000 54800
rect 0 54408 800 54528
rect 31200 54136 32000 54256
rect 0 53728 800 53848
rect 31200 53728 32000 53848
rect 0 53048 800 53168
rect 31200 53184 32000 53304
rect 31200 52776 32000 52896
rect 0 52368 800 52488
rect 31200 52232 32000 52352
rect 0 51824 800 51944
rect 31200 51824 32000 51944
rect 31200 51416 32000 51536
rect 0 51144 800 51264
rect 31200 50872 32000 50992
rect 0 50464 800 50584
rect 31200 50464 32000 50584
rect 0 49784 800 49904
rect 31200 49920 32000 50040
rect 31200 49512 32000 49632
rect 0 49104 800 49224
rect 31200 48968 32000 49088
rect 0 48424 800 48544
rect 31200 48560 32000 48680
rect 31200 48016 32000 48136
rect 0 47744 800 47864
rect 31200 47608 32000 47728
rect 0 47200 800 47320
rect 31200 47064 32000 47184
rect 0 46520 800 46640
rect 31200 46656 32000 46776
rect 31200 46112 32000 46232
rect 0 45840 800 45960
rect 31200 45704 32000 45824
rect 0 45160 800 45280
rect 31200 45296 32000 45416
rect 31200 44752 32000 44872
rect 0 44480 800 44600
rect 31200 44344 32000 44464
rect 0 43800 800 43920
rect 31200 43800 32000 43920
rect 31200 43392 32000 43512
rect 0 43120 800 43240
rect 31200 42848 32000 42968
rect 0 42576 800 42696
rect 31200 42440 32000 42560
rect 0 41896 800 42016
rect 31200 41896 32000 42016
rect 31200 41488 32000 41608
rect 0 41216 800 41336
rect 31200 40944 32000 41064
rect 0 40536 800 40656
rect 31200 40536 32000 40656
rect 31200 40128 32000 40248
rect 0 39856 800 39976
rect 31200 39584 32000 39704
rect 0 39176 800 39296
rect 31200 39176 32000 39296
rect 0 38496 800 38616
rect 31200 38632 32000 38752
rect 31200 38224 32000 38344
rect 0 37816 800 37936
rect 31200 37680 32000 37800
rect 0 37272 800 37392
rect 31200 37272 32000 37392
rect 0 36592 800 36712
rect 31200 36728 32000 36848
rect 31200 36320 32000 36440
rect 0 35912 800 36032
rect 31200 35776 32000 35896
rect 0 35232 800 35352
rect 31200 35368 32000 35488
rect 31200 34824 32000 34944
rect 0 34552 800 34672
rect 31200 34416 32000 34536
rect 0 33872 800 33992
rect 31200 34008 32000 34128
rect 31200 33464 32000 33584
rect 0 33192 800 33312
rect 31200 33056 32000 33176
rect 0 32648 800 32768
rect 31200 32512 32000 32632
rect 0 31968 800 32088
rect 31200 32104 32000 32224
rect 31200 31560 32000 31680
rect 0 31288 800 31408
rect 31200 31152 32000 31272
rect 0 30608 800 30728
rect 31200 30608 32000 30728
rect 31200 30200 32000 30320
rect 0 29928 800 30048
rect 31200 29656 32000 29776
rect 0 29248 800 29368
rect 31200 29248 32000 29368
rect 0 28568 800 28688
rect 31200 28704 32000 28824
rect 31200 28296 32000 28416
rect 0 28024 800 28144
rect 31200 27888 32000 28008
rect 0 27344 800 27464
rect 31200 27344 32000 27464
rect 31200 26936 32000 27056
rect 0 26664 800 26784
rect 31200 26392 32000 26512
rect 0 25984 800 26104
rect 31200 25984 32000 26104
rect 0 25304 800 25424
rect 31200 25440 32000 25560
rect 31200 25032 32000 25152
rect 0 24624 800 24744
rect 31200 24488 32000 24608
rect 0 23944 800 24064
rect 31200 24080 32000 24200
rect 0 23400 800 23520
rect 31200 23536 32000 23656
rect 31200 23128 32000 23248
rect 0 22720 800 22840
rect 31200 22720 32000 22840
rect 0 22040 800 22160
rect 31200 22176 32000 22296
rect 31200 21768 32000 21888
rect 0 21360 800 21480
rect 31200 21224 32000 21344
rect 0 20680 800 20800
rect 31200 20816 32000 20936
rect 31200 20272 32000 20392
rect 0 20000 800 20120
rect 31200 19864 32000 19984
rect 0 19320 800 19440
rect 31200 19320 32000 19440
rect 0 18776 800 18896
rect 31200 18912 32000 19032
rect 31200 18368 32000 18488
rect 0 18096 800 18216
rect 31200 17960 32000 18080
rect 0 17416 800 17536
rect 31200 17416 32000 17536
rect 31200 17008 32000 17128
rect 0 16736 800 16856
rect 31200 16600 32000 16720
rect 0 16056 800 16176
rect 31200 16056 32000 16176
rect 31200 15648 32000 15768
rect 0 15376 800 15496
rect 31200 15104 32000 15224
rect 0 14696 800 14816
rect 31200 14696 32000 14816
rect 0 14152 800 14272
rect 31200 14152 32000 14272
rect 31200 13744 32000 13864
rect 0 13472 800 13592
rect 31200 13200 32000 13320
rect 0 12792 800 12912
rect 31200 12792 32000 12912
rect 0 12112 800 12232
rect 31200 12248 32000 12368
rect 31200 11840 32000 11960
rect 0 11432 800 11552
rect 31200 11432 32000 11552
rect 0 10752 800 10872
rect 31200 10888 32000 11008
rect 31200 10480 32000 10600
rect 0 10072 800 10192
rect 31200 9936 32000 10056
rect 0 9528 800 9648
rect 31200 9528 32000 9648
rect 0 8848 800 8968
rect 31200 8984 32000 9104
rect 31200 8576 32000 8696
rect 0 8168 800 8288
rect 31200 8032 32000 8152
rect 0 7488 800 7608
rect 31200 7624 32000 7744
rect 31200 7080 32000 7200
rect 0 6808 800 6928
rect 31200 6672 32000 6792
rect 0 6128 800 6248
rect 31200 6128 32000 6248
rect 31200 5720 32000 5840
rect 0 5448 800 5568
rect 31200 5312 32000 5432
rect 0 4904 800 5024
rect 31200 4768 32000 4888
rect 0 4224 800 4344
rect 31200 4360 32000 4480
rect 31200 3816 32000 3936
rect 0 3544 800 3664
rect 31200 3408 32000 3528
rect 0 2864 800 2984
rect 31200 2864 32000 2984
rect 31200 2456 32000 2576
rect 0 2184 800 2304
rect 31200 1912 32000 2032
rect 0 1504 800 1624
rect 31200 1504 32000 1624
rect 0 824 800 944
rect 31200 960 32000 1080
rect 31200 552 32000 672
rect 0 280 800 400
rect 31200 144 32000 264
<< obsm3 >>
rect 880 79488 31120 79661
rect 800 79360 31962 79488
rect 800 79088 31120 79360
rect 880 79080 31120 79088
rect 880 78816 31962 79080
rect 880 78808 31120 78816
rect 800 78536 31120 78808
rect 800 78408 31962 78536
rect 880 78128 31120 78408
rect 800 77864 31962 78128
rect 800 77728 31120 77864
rect 880 77584 31120 77728
rect 880 77456 31962 77584
rect 880 77448 31120 77456
rect 800 77176 31120 77448
rect 800 77048 31962 77176
rect 880 76912 31962 77048
rect 880 76768 31120 76912
rect 800 76632 31120 76768
rect 800 76504 31962 76632
rect 800 76368 31120 76504
rect 880 76224 31120 76368
rect 880 76088 31962 76224
rect 800 75960 31962 76088
rect 800 75688 31120 75960
rect 880 75680 31120 75688
rect 880 75552 31962 75680
rect 880 75408 31120 75552
rect 800 75272 31120 75408
rect 800 75144 31962 75272
rect 880 75008 31962 75144
rect 880 74864 31120 75008
rect 800 74728 31120 74864
rect 800 74600 31962 74728
rect 800 74464 31120 74600
rect 880 74320 31120 74464
rect 880 74192 31962 74320
rect 880 74184 31120 74192
rect 800 73912 31120 74184
rect 800 73784 31962 73912
rect 880 73648 31962 73784
rect 880 73504 31120 73648
rect 800 73368 31120 73504
rect 800 73240 31962 73368
rect 800 73104 31120 73240
rect 880 72960 31120 73104
rect 880 72824 31962 72960
rect 800 72696 31962 72824
rect 800 72424 31120 72696
rect 880 72416 31120 72424
rect 880 72288 31962 72416
rect 880 72144 31120 72288
rect 800 72008 31120 72144
rect 800 71744 31962 72008
rect 880 71464 31120 71744
rect 800 71336 31962 71464
rect 800 71064 31120 71336
rect 880 71056 31120 71064
rect 880 70792 31962 71056
rect 880 70784 31120 70792
rect 800 70520 31120 70784
rect 880 70512 31120 70520
rect 880 70384 31962 70512
rect 880 70240 31120 70384
rect 800 70104 31120 70240
rect 800 69840 31962 70104
rect 880 69560 31120 69840
rect 800 69432 31962 69560
rect 800 69160 31120 69432
rect 880 69152 31120 69160
rect 880 68888 31962 69152
rect 880 68880 31120 68888
rect 800 68608 31120 68880
rect 800 68480 31962 68608
rect 880 68200 31120 68480
rect 800 68072 31962 68200
rect 800 67800 31120 68072
rect 880 67792 31120 67800
rect 880 67528 31962 67792
rect 880 67520 31120 67528
rect 800 67248 31120 67520
rect 800 67120 31962 67248
rect 880 66840 31120 67120
rect 800 66576 31962 66840
rect 800 66440 31120 66576
rect 880 66296 31120 66440
rect 880 66168 31962 66296
rect 880 66160 31120 66168
rect 800 65896 31120 66160
rect 880 65888 31120 65896
rect 880 65624 31962 65888
rect 880 65616 31120 65624
rect 800 65344 31120 65616
rect 800 65216 31962 65344
rect 880 64936 31120 65216
rect 800 64672 31962 64936
rect 800 64536 31120 64672
rect 880 64392 31120 64536
rect 880 64264 31962 64392
rect 880 64256 31120 64264
rect 800 63984 31120 64256
rect 800 63856 31962 63984
rect 880 63720 31962 63856
rect 880 63576 31120 63720
rect 800 63440 31120 63576
rect 800 63312 31962 63440
rect 800 63176 31120 63312
rect 880 63032 31120 63176
rect 880 62904 31962 63032
rect 880 62896 31120 62904
rect 800 62624 31120 62896
rect 800 62496 31962 62624
rect 880 62360 31962 62496
rect 880 62216 31120 62360
rect 800 62080 31120 62216
rect 800 61952 31962 62080
rect 800 61816 31120 61952
rect 880 61672 31120 61816
rect 880 61536 31962 61672
rect 800 61408 31962 61536
rect 800 61272 31120 61408
rect 880 61128 31120 61272
rect 880 61000 31962 61128
rect 880 60992 31120 61000
rect 800 60720 31120 60992
rect 800 60592 31962 60720
rect 880 60456 31962 60592
rect 880 60312 31120 60456
rect 800 60176 31120 60312
rect 800 60048 31962 60176
rect 800 59912 31120 60048
rect 880 59768 31120 59912
rect 880 59632 31962 59768
rect 800 59504 31962 59632
rect 800 59232 31120 59504
rect 880 59224 31120 59232
rect 880 59096 31962 59224
rect 880 58952 31120 59096
rect 800 58816 31120 58952
rect 800 58552 31962 58816
rect 880 58272 31120 58552
rect 800 58144 31962 58272
rect 800 57872 31120 58144
rect 880 57864 31120 57872
rect 880 57600 31962 57864
rect 880 57592 31120 57600
rect 800 57320 31120 57592
rect 800 57192 31962 57320
rect 880 56912 31120 57192
rect 800 56784 31962 56912
rect 800 56648 31120 56784
rect 880 56504 31120 56648
rect 880 56368 31962 56504
rect 800 56240 31962 56368
rect 800 55968 31120 56240
rect 880 55960 31120 55968
rect 880 55832 31962 55960
rect 880 55688 31120 55832
rect 800 55552 31120 55688
rect 800 55288 31962 55552
rect 880 55008 31120 55288
rect 800 54880 31962 55008
rect 800 54608 31120 54880
rect 880 54600 31120 54608
rect 880 54336 31962 54600
rect 880 54328 31120 54336
rect 800 54056 31120 54328
rect 800 53928 31962 54056
rect 880 53648 31120 53928
rect 800 53384 31962 53648
rect 800 53248 31120 53384
rect 880 53104 31120 53248
rect 880 52976 31962 53104
rect 880 52968 31120 52976
rect 800 52696 31120 52968
rect 800 52568 31962 52696
rect 880 52432 31962 52568
rect 880 52288 31120 52432
rect 800 52152 31120 52288
rect 800 52024 31962 52152
rect 880 51744 31120 52024
rect 800 51616 31962 51744
rect 800 51344 31120 51616
rect 880 51336 31120 51344
rect 880 51072 31962 51336
rect 880 51064 31120 51072
rect 800 50792 31120 51064
rect 800 50664 31962 50792
rect 880 50384 31120 50664
rect 800 50120 31962 50384
rect 800 49984 31120 50120
rect 880 49840 31120 49984
rect 880 49712 31962 49840
rect 880 49704 31120 49712
rect 800 49432 31120 49704
rect 800 49304 31962 49432
rect 880 49168 31962 49304
rect 880 49024 31120 49168
rect 800 48888 31120 49024
rect 800 48760 31962 48888
rect 800 48624 31120 48760
rect 880 48480 31120 48624
rect 880 48344 31962 48480
rect 800 48216 31962 48344
rect 800 47944 31120 48216
rect 880 47936 31120 47944
rect 880 47808 31962 47936
rect 880 47664 31120 47808
rect 800 47528 31120 47664
rect 800 47400 31962 47528
rect 880 47264 31962 47400
rect 880 47120 31120 47264
rect 800 46984 31120 47120
rect 800 46856 31962 46984
rect 800 46720 31120 46856
rect 880 46576 31120 46720
rect 880 46440 31962 46576
rect 800 46312 31962 46440
rect 800 46040 31120 46312
rect 880 46032 31120 46040
rect 880 45904 31962 46032
rect 880 45760 31120 45904
rect 800 45624 31120 45760
rect 800 45496 31962 45624
rect 800 45360 31120 45496
rect 880 45216 31120 45360
rect 880 45080 31962 45216
rect 800 44952 31962 45080
rect 800 44680 31120 44952
rect 880 44672 31120 44680
rect 880 44544 31962 44672
rect 880 44400 31120 44544
rect 800 44264 31120 44400
rect 800 44000 31962 44264
rect 880 43720 31120 44000
rect 800 43592 31962 43720
rect 800 43320 31120 43592
rect 880 43312 31120 43320
rect 880 43048 31962 43312
rect 880 43040 31120 43048
rect 800 42776 31120 43040
rect 880 42768 31120 42776
rect 880 42640 31962 42768
rect 880 42496 31120 42640
rect 800 42360 31120 42496
rect 800 42096 31962 42360
rect 880 41816 31120 42096
rect 800 41688 31962 41816
rect 800 41416 31120 41688
rect 880 41408 31120 41416
rect 880 41144 31962 41408
rect 880 41136 31120 41144
rect 800 40864 31120 41136
rect 800 40736 31962 40864
rect 880 40456 31120 40736
rect 800 40328 31962 40456
rect 800 40056 31120 40328
rect 880 40048 31120 40056
rect 880 39784 31962 40048
rect 880 39776 31120 39784
rect 800 39504 31120 39776
rect 800 39376 31962 39504
rect 880 39096 31120 39376
rect 800 38832 31962 39096
rect 800 38696 31120 38832
rect 880 38552 31120 38696
rect 880 38424 31962 38552
rect 880 38416 31120 38424
rect 800 38144 31120 38416
rect 800 38016 31962 38144
rect 880 37880 31962 38016
rect 880 37736 31120 37880
rect 800 37600 31120 37736
rect 800 37472 31962 37600
rect 880 37192 31120 37472
rect 800 36928 31962 37192
rect 800 36792 31120 36928
rect 880 36648 31120 36792
rect 880 36520 31962 36648
rect 880 36512 31120 36520
rect 800 36240 31120 36512
rect 800 36112 31962 36240
rect 880 35976 31962 36112
rect 880 35832 31120 35976
rect 800 35696 31120 35832
rect 800 35568 31962 35696
rect 800 35432 31120 35568
rect 880 35288 31120 35432
rect 880 35152 31962 35288
rect 800 35024 31962 35152
rect 800 34752 31120 35024
rect 880 34744 31120 34752
rect 880 34616 31962 34744
rect 880 34472 31120 34616
rect 800 34336 31120 34472
rect 800 34208 31962 34336
rect 800 34072 31120 34208
rect 880 33928 31120 34072
rect 880 33792 31962 33928
rect 800 33664 31962 33792
rect 800 33392 31120 33664
rect 880 33384 31120 33392
rect 880 33256 31962 33384
rect 880 33112 31120 33256
rect 800 32976 31120 33112
rect 800 32848 31962 32976
rect 880 32712 31962 32848
rect 880 32568 31120 32712
rect 800 32432 31120 32568
rect 800 32304 31962 32432
rect 800 32168 31120 32304
rect 880 32024 31120 32168
rect 880 31888 31962 32024
rect 800 31760 31962 31888
rect 800 31488 31120 31760
rect 880 31480 31120 31488
rect 880 31352 31962 31480
rect 880 31208 31120 31352
rect 800 31072 31120 31208
rect 800 30808 31962 31072
rect 880 30528 31120 30808
rect 800 30400 31962 30528
rect 800 30128 31120 30400
rect 880 30120 31120 30128
rect 880 29856 31962 30120
rect 880 29848 31120 29856
rect 800 29576 31120 29848
rect 800 29448 31962 29576
rect 880 29168 31120 29448
rect 800 28904 31962 29168
rect 800 28768 31120 28904
rect 880 28624 31120 28768
rect 880 28496 31962 28624
rect 880 28488 31120 28496
rect 800 28224 31120 28488
rect 880 28216 31120 28224
rect 880 28088 31962 28216
rect 880 27944 31120 28088
rect 800 27808 31120 27944
rect 800 27544 31962 27808
rect 880 27264 31120 27544
rect 800 27136 31962 27264
rect 800 26864 31120 27136
rect 880 26856 31120 26864
rect 880 26592 31962 26856
rect 880 26584 31120 26592
rect 800 26312 31120 26584
rect 800 26184 31962 26312
rect 880 25904 31120 26184
rect 800 25640 31962 25904
rect 800 25504 31120 25640
rect 880 25360 31120 25504
rect 880 25232 31962 25360
rect 880 25224 31120 25232
rect 800 24952 31120 25224
rect 800 24824 31962 24952
rect 880 24688 31962 24824
rect 880 24544 31120 24688
rect 800 24408 31120 24544
rect 800 24280 31962 24408
rect 800 24144 31120 24280
rect 880 24000 31120 24144
rect 880 23864 31962 24000
rect 800 23736 31962 23864
rect 800 23600 31120 23736
rect 880 23456 31120 23600
rect 880 23328 31962 23456
rect 880 23320 31120 23328
rect 800 23048 31120 23320
rect 800 22920 31962 23048
rect 880 22640 31120 22920
rect 800 22376 31962 22640
rect 800 22240 31120 22376
rect 880 22096 31120 22240
rect 880 21968 31962 22096
rect 880 21960 31120 21968
rect 800 21688 31120 21960
rect 800 21560 31962 21688
rect 880 21424 31962 21560
rect 880 21280 31120 21424
rect 800 21144 31120 21280
rect 800 21016 31962 21144
rect 800 20880 31120 21016
rect 880 20736 31120 20880
rect 880 20600 31962 20736
rect 800 20472 31962 20600
rect 800 20200 31120 20472
rect 880 20192 31120 20200
rect 880 20064 31962 20192
rect 880 19920 31120 20064
rect 800 19784 31120 19920
rect 800 19520 31962 19784
rect 880 19240 31120 19520
rect 800 19112 31962 19240
rect 800 18976 31120 19112
rect 880 18832 31120 18976
rect 880 18696 31962 18832
rect 800 18568 31962 18696
rect 800 18296 31120 18568
rect 880 18288 31120 18296
rect 880 18160 31962 18288
rect 880 18016 31120 18160
rect 800 17880 31120 18016
rect 800 17616 31962 17880
rect 880 17336 31120 17616
rect 800 17208 31962 17336
rect 800 16936 31120 17208
rect 880 16928 31120 16936
rect 880 16800 31962 16928
rect 880 16656 31120 16800
rect 800 16520 31120 16656
rect 800 16256 31962 16520
rect 880 15976 31120 16256
rect 800 15848 31962 15976
rect 800 15576 31120 15848
rect 880 15568 31120 15576
rect 880 15304 31962 15568
rect 880 15296 31120 15304
rect 800 15024 31120 15296
rect 800 14896 31962 15024
rect 880 14616 31120 14896
rect 800 14352 31962 14616
rect 880 14072 31120 14352
rect 800 13944 31962 14072
rect 800 13672 31120 13944
rect 880 13664 31120 13672
rect 880 13400 31962 13664
rect 880 13392 31120 13400
rect 800 13120 31120 13392
rect 800 12992 31962 13120
rect 880 12712 31120 12992
rect 800 12448 31962 12712
rect 800 12312 31120 12448
rect 880 12168 31120 12312
rect 880 12040 31962 12168
rect 880 12032 31120 12040
rect 800 11760 31120 12032
rect 800 11632 31962 11760
rect 880 11352 31120 11632
rect 800 11088 31962 11352
rect 800 10952 31120 11088
rect 880 10808 31120 10952
rect 880 10680 31962 10808
rect 880 10672 31120 10680
rect 800 10400 31120 10672
rect 800 10272 31962 10400
rect 880 10136 31962 10272
rect 880 9992 31120 10136
rect 800 9856 31120 9992
rect 800 9728 31962 9856
rect 880 9448 31120 9728
rect 800 9184 31962 9448
rect 800 9048 31120 9184
rect 880 8904 31120 9048
rect 880 8776 31962 8904
rect 880 8768 31120 8776
rect 800 8496 31120 8768
rect 800 8368 31962 8496
rect 880 8232 31962 8368
rect 880 8088 31120 8232
rect 800 7952 31120 8088
rect 800 7824 31962 7952
rect 800 7688 31120 7824
rect 880 7544 31120 7688
rect 880 7408 31962 7544
rect 800 7280 31962 7408
rect 800 7008 31120 7280
rect 880 7000 31120 7008
rect 880 6872 31962 7000
rect 880 6728 31120 6872
rect 800 6592 31120 6728
rect 800 6328 31962 6592
rect 880 6048 31120 6328
rect 800 5920 31962 6048
rect 800 5648 31120 5920
rect 880 5640 31120 5648
rect 880 5512 31962 5640
rect 880 5368 31120 5512
rect 800 5232 31120 5368
rect 800 5104 31962 5232
rect 880 4968 31962 5104
rect 880 4824 31120 4968
rect 800 4688 31120 4824
rect 800 4560 31962 4688
rect 800 4424 31120 4560
rect 880 4280 31120 4424
rect 880 4144 31962 4280
rect 800 4016 31962 4144
rect 800 3744 31120 4016
rect 880 3736 31120 3744
rect 880 3608 31962 3736
rect 880 3464 31120 3608
rect 800 3328 31120 3464
rect 800 3064 31962 3328
rect 880 2784 31120 3064
rect 800 2656 31962 2784
rect 800 2384 31120 2656
rect 880 2376 31120 2384
rect 880 2112 31962 2376
rect 880 2104 31120 2112
rect 800 1832 31120 2104
rect 800 1704 31962 1832
rect 880 1424 31120 1704
rect 800 1160 31962 1424
rect 800 1024 31120 1160
rect 880 880 31120 1024
rect 880 752 31962 880
rect 880 744 31120 752
rect 800 480 31120 744
rect 880 472 31120 480
rect 880 344 31962 472
rect 880 200 31120 344
rect 800 171 31120 200
<< metal4 >>
rect 5910 2128 6230 77840
rect 10874 2128 11194 77840
rect 15840 2128 16160 77840
rect 20805 2128 21125 77840
rect 25771 2128 26091 77840
<< obsm4 >>
rect 6310 2128 10794 77840
rect 11274 2128 15760 77840
rect 16240 2128 20725 77840
rect 21205 2128 25691 77840
rect 26171 2128 31957 77840
<< labels >>
rlabel metal3 s 0 4904 800 5024 6 ram_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 ram_addr0[1]
port 2 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 ram_addr0[2]
port 3 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 ram_addr0[3]
port 4 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 ram_addr0[4]
port 5 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 ram_addr0[5]
port 6 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 ram_addr0[6]
port 7 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 ram_addr0[7]
port 8 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 ram_addr1[0]
port 9 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 ram_addr1[1]
port 10 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 ram_addr1[2]
port 11 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 ram_addr1[3]
port 12 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 ram_addr1[4]
port 13 nsew signal output
rlabel metal3 s 0 56992 800 57112 6 ram_addr1[5]
port 14 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 ram_addr1[6]
port 15 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 ram_addr1[7]
port 16 nsew signal output
rlabel metal3 s 0 280 800 400 6 ram_clk0
port 17 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 ram_clk1
port 18 nsew signal output
rlabel metal3 s 0 824 800 944 6 ram_csb0
port 19 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 ram_csb1
port 20 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 ram_din0[0]
port 21 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 ram_din0[10]
port 22 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 ram_din0[11]
port 23 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 ram_din0[12]
port 24 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 ram_din0[13]
port 25 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 ram_din0[14]
port 26 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 ram_din0[15]
port 27 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 ram_din0[16]
port 28 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 ram_din0[17]
port 29 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 ram_din0[18]
port 30 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 ram_din0[19]
port 31 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 ram_din0[1]
port 32 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 ram_din0[20]
port 33 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 ram_din0[21]
port 34 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 ram_din0[22]
port 35 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 ram_din0[23]
port 36 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 ram_din0[24]
port 37 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 ram_din0[25]
port 38 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 ram_din0[26]
port 39 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 ram_din0[27]
port 40 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 ram_din0[28]
port 41 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 ram_din0[29]
port 42 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 ram_din0[2]
port 43 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 ram_din0[30]
port 44 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 ram_din0[31]
port 45 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 ram_din0[3]
port 46 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 ram_din0[4]
port 47 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 ram_din0[5]
port 48 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 ram_din0[6]
port 49 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 ram_din0[7]
port 50 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 ram_din0[8]
port 51 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 ram_din0[9]
port 52 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 ram_dout0[0]
port 53 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 ram_dout0[10]
port 54 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 ram_dout0[11]
port 55 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 ram_dout0[12]
port 56 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 ram_dout0[13]
port 57 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 ram_dout0[14]
port 58 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 ram_dout0[15]
port 59 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 ram_dout0[16]
port 60 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 ram_dout0[17]
port 61 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 ram_dout0[18]
port 62 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 ram_dout0[19]
port 63 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 ram_dout0[1]
port 64 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 ram_dout0[20]
port 65 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 ram_dout0[21]
port 66 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 ram_dout0[22]
port 67 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 ram_dout0[23]
port 68 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 ram_dout0[24]
port 69 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 ram_dout0[25]
port 70 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 ram_dout0[26]
port 71 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 ram_dout0[27]
port 72 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 ram_dout0[28]
port 73 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 ram_dout0[29]
port 74 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 ram_dout0[2]
port 75 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 ram_dout0[30]
port 76 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 ram_dout0[31]
port 77 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 ram_dout0[3]
port 78 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 ram_dout0[4]
port 79 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 ram_dout0[5]
port 80 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 ram_dout0[6]
port 81 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 ram_dout0[7]
port 82 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 ram_dout0[8]
port 83 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 ram_dout0[9]
port 84 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 ram_dout1[0]
port 85 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 ram_dout1[10]
port 86 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 ram_dout1[11]
port 87 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 ram_dout1[12]
port 88 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 ram_dout1[13]
port 89 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 ram_dout1[14]
port 90 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 ram_dout1[15]
port 91 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 ram_dout1[16]
port 92 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 ram_dout1[17]
port 93 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 ram_dout1[18]
port 94 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 ram_dout1[19]
port 95 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 ram_dout1[1]
port 96 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 ram_dout1[20]
port 97 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 ram_dout1[21]
port 98 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 ram_dout1[22]
port 99 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 ram_dout1[23]
port 100 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 ram_dout1[24]
port 101 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 ram_dout1[25]
port 102 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 ram_dout1[26]
port 103 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 ram_dout1[27]
port 104 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 ram_dout1[28]
port 105 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 ram_dout1[29]
port 106 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 ram_dout1[2]
port 107 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 ram_dout1[30]
port 108 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 ram_dout1[31]
port 109 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 ram_dout1[3]
port 110 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 ram_dout1[4]
port 111 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 ram_dout1[5]
port 112 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 ram_dout1[6]
port 113 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 ram_dout1[7]
port 114 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 ram_dout1[8]
port 115 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 ram_dout1[9]
port 116 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 ram_web0
port 117 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 ram_wmask0[0]
port 118 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 ram_wmask0[1]
port 119 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 ram_wmask0[2]
port 120 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 ram_wmask0[3]
port 121 nsew signal output
rlabel metal4 s 5910 2128 6230 77840 6 vccd1
port 122 nsew power input
rlabel metal4 s 15840 2128 16160 77840 6 vccd1
port 122 nsew power input
rlabel metal4 s 25771 2128 26091 77840 6 vccd1
port 122 nsew power input
rlabel metal4 s 10874 2128 11194 77840 6 vssd1
port 123 nsew ground input
rlabel metal4 s 20805 2128 21125 77840 6 vssd1
port 123 nsew ground input
rlabel metal3 s 31200 552 32000 672 6 wb_a_clk_i
port 124 nsew signal input
rlabel metal3 s 31200 960 32000 1080 6 wb_a_rst_i
port 125 nsew signal input
rlabel metal3 s 31200 40536 32000 40656 6 wb_b_clk_i
port 126 nsew signal input
rlabel metal3 s 31200 40944 32000 41064 6 wb_b_rst_i
port 127 nsew signal input
rlabel metal3 s 31200 2864 32000 2984 6 wbs_a_ack_o
port 128 nsew signal output
rlabel metal3 s 31200 5312 32000 5432 6 wbs_a_adr_i[0]
port 129 nsew signal input
rlabel metal3 s 31200 9936 32000 10056 6 wbs_a_adr_i[10]
port 130 nsew signal input
rlabel metal3 s 31200 5720 32000 5840 6 wbs_a_adr_i[1]
port 131 nsew signal input
rlabel metal3 s 31200 6128 32000 6248 6 wbs_a_adr_i[2]
port 132 nsew signal input
rlabel metal3 s 31200 6672 32000 6792 6 wbs_a_adr_i[3]
port 133 nsew signal input
rlabel metal3 s 31200 7080 32000 7200 6 wbs_a_adr_i[4]
port 134 nsew signal input
rlabel metal3 s 31200 7624 32000 7744 6 wbs_a_adr_i[5]
port 135 nsew signal input
rlabel metal3 s 31200 8032 32000 8152 6 wbs_a_adr_i[6]
port 136 nsew signal input
rlabel metal3 s 31200 8576 32000 8696 6 wbs_a_adr_i[7]
port 137 nsew signal input
rlabel metal3 s 31200 8984 32000 9104 6 wbs_a_adr_i[8]
port 138 nsew signal input
rlabel metal3 s 31200 9528 32000 9648 6 wbs_a_adr_i[9]
port 139 nsew signal input
rlabel metal3 s 31200 1912 32000 2032 6 wbs_a_cyc_i
port 140 nsew signal input
rlabel metal3 s 31200 10480 32000 10600 6 wbs_a_dat_i[0]
port 141 nsew signal input
rlabel metal3 s 31200 15104 32000 15224 6 wbs_a_dat_i[10]
port 142 nsew signal input
rlabel metal3 s 31200 15648 32000 15768 6 wbs_a_dat_i[11]
port 143 nsew signal input
rlabel metal3 s 31200 16056 32000 16176 6 wbs_a_dat_i[12]
port 144 nsew signal input
rlabel metal3 s 31200 16600 32000 16720 6 wbs_a_dat_i[13]
port 145 nsew signal input
rlabel metal3 s 31200 17008 32000 17128 6 wbs_a_dat_i[14]
port 146 nsew signal input
rlabel metal3 s 31200 17416 32000 17536 6 wbs_a_dat_i[15]
port 147 nsew signal input
rlabel metal3 s 31200 17960 32000 18080 6 wbs_a_dat_i[16]
port 148 nsew signal input
rlabel metal3 s 31200 18368 32000 18488 6 wbs_a_dat_i[17]
port 149 nsew signal input
rlabel metal3 s 31200 18912 32000 19032 6 wbs_a_dat_i[18]
port 150 nsew signal input
rlabel metal3 s 31200 19320 32000 19440 6 wbs_a_dat_i[19]
port 151 nsew signal input
rlabel metal3 s 31200 10888 32000 11008 6 wbs_a_dat_i[1]
port 152 nsew signal input
rlabel metal3 s 31200 19864 32000 19984 6 wbs_a_dat_i[20]
port 153 nsew signal input
rlabel metal3 s 31200 20272 32000 20392 6 wbs_a_dat_i[21]
port 154 nsew signal input
rlabel metal3 s 31200 20816 32000 20936 6 wbs_a_dat_i[22]
port 155 nsew signal input
rlabel metal3 s 31200 21224 32000 21344 6 wbs_a_dat_i[23]
port 156 nsew signal input
rlabel metal3 s 31200 21768 32000 21888 6 wbs_a_dat_i[24]
port 157 nsew signal input
rlabel metal3 s 31200 22176 32000 22296 6 wbs_a_dat_i[25]
port 158 nsew signal input
rlabel metal3 s 31200 22720 32000 22840 6 wbs_a_dat_i[26]
port 159 nsew signal input
rlabel metal3 s 31200 23128 32000 23248 6 wbs_a_dat_i[27]
port 160 nsew signal input
rlabel metal3 s 31200 23536 32000 23656 6 wbs_a_dat_i[28]
port 161 nsew signal input
rlabel metal3 s 31200 24080 32000 24200 6 wbs_a_dat_i[29]
port 162 nsew signal input
rlabel metal3 s 31200 11432 32000 11552 6 wbs_a_dat_i[2]
port 163 nsew signal input
rlabel metal3 s 31200 24488 32000 24608 6 wbs_a_dat_i[30]
port 164 nsew signal input
rlabel metal3 s 31200 25032 32000 25152 6 wbs_a_dat_i[31]
port 165 nsew signal input
rlabel metal3 s 31200 11840 32000 11960 6 wbs_a_dat_i[3]
port 166 nsew signal input
rlabel metal3 s 31200 12248 32000 12368 6 wbs_a_dat_i[4]
port 167 nsew signal input
rlabel metal3 s 31200 12792 32000 12912 6 wbs_a_dat_i[5]
port 168 nsew signal input
rlabel metal3 s 31200 13200 32000 13320 6 wbs_a_dat_i[6]
port 169 nsew signal input
rlabel metal3 s 31200 13744 32000 13864 6 wbs_a_dat_i[7]
port 170 nsew signal input
rlabel metal3 s 31200 14152 32000 14272 6 wbs_a_dat_i[8]
port 171 nsew signal input
rlabel metal3 s 31200 14696 32000 14816 6 wbs_a_dat_i[9]
port 172 nsew signal input
rlabel metal3 s 31200 25440 32000 25560 6 wbs_a_dat_o[0]
port 173 nsew signal output
rlabel metal3 s 31200 30200 32000 30320 6 wbs_a_dat_o[10]
port 174 nsew signal output
rlabel metal3 s 31200 30608 32000 30728 6 wbs_a_dat_o[11]
port 175 nsew signal output
rlabel metal3 s 31200 31152 32000 31272 6 wbs_a_dat_o[12]
port 176 nsew signal output
rlabel metal3 s 31200 31560 32000 31680 6 wbs_a_dat_o[13]
port 177 nsew signal output
rlabel metal3 s 31200 32104 32000 32224 6 wbs_a_dat_o[14]
port 178 nsew signal output
rlabel metal3 s 31200 32512 32000 32632 6 wbs_a_dat_o[15]
port 179 nsew signal output
rlabel metal3 s 31200 33056 32000 33176 6 wbs_a_dat_o[16]
port 180 nsew signal output
rlabel metal3 s 31200 33464 32000 33584 6 wbs_a_dat_o[17]
port 181 nsew signal output
rlabel metal3 s 31200 34008 32000 34128 6 wbs_a_dat_o[18]
port 182 nsew signal output
rlabel metal3 s 31200 34416 32000 34536 6 wbs_a_dat_o[19]
port 183 nsew signal output
rlabel metal3 s 31200 25984 32000 26104 6 wbs_a_dat_o[1]
port 184 nsew signal output
rlabel metal3 s 31200 34824 32000 34944 6 wbs_a_dat_o[20]
port 185 nsew signal output
rlabel metal3 s 31200 35368 32000 35488 6 wbs_a_dat_o[21]
port 186 nsew signal output
rlabel metal3 s 31200 35776 32000 35896 6 wbs_a_dat_o[22]
port 187 nsew signal output
rlabel metal3 s 31200 36320 32000 36440 6 wbs_a_dat_o[23]
port 188 nsew signal output
rlabel metal3 s 31200 36728 32000 36848 6 wbs_a_dat_o[24]
port 189 nsew signal output
rlabel metal3 s 31200 37272 32000 37392 6 wbs_a_dat_o[25]
port 190 nsew signal output
rlabel metal3 s 31200 37680 32000 37800 6 wbs_a_dat_o[26]
port 191 nsew signal output
rlabel metal3 s 31200 38224 32000 38344 6 wbs_a_dat_o[27]
port 192 nsew signal output
rlabel metal3 s 31200 38632 32000 38752 6 wbs_a_dat_o[28]
port 193 nsew signal output
rlabel metal3 s 31200 39176 32000 39296 6 wbs_a_dat_o[29]
port 194 nsew signal output
rlabel metal3 s 31200 26392 32000 26512 6 wbs_a_dat_o[2]
port 195 nsew signal output
rlabel metal3 s 31200 39584 32000 39704 6 wbs_a_dat_o[30]
port 196 nsew signal output
rlabel metal3 s 31200 40128 32000 40248 6 wbs_a_dat_o[31]
port 197 nsew signal output
rlabel metal3 s 31200 26936 32000 27056 6 wbs_a_dat_o[3]
port 198 nsew signal output
rlabel metal3 s 31200 27344 32000 27464 6 wbs_a_dat_o[4]
port 199 nsew signal output
rlabel metal3 s 31200 27888 32000 28008 6 wbs_a_dat_o[5]
port 200 nsew signal output
rlabel metal3 s 31200 28296 32000 28416 6 wbs_a_dat_o[6]
port 201 nsew signal output
rlabel metal3 s 31200 28704 32000 28824 6 wbs_a_dat_o[7]
port 202 nsew signal output
rlabel metal3 s 31200 29248 32000 29368 6 wbs_a_dat_o[8]
port 203 nsew signal output
rlabel metal3 s 31200 29656 32000 29776 6 wbs_a_dat_o[9]
port 204 nsew signal output
rlabel metal3 s 31200 3408 32000 3528 6 wbs_a_sel_i[0]
port 205 nsew signal input
rlabel metal3 s 31200 3816 32000 3936 6 wbs_a_sel_i[1]
port 206 nsew signal input
rlabel metal3 s 31200 4360 32000 4480 6 wbs_a_sel_i[2]
port 207 nsew signal input
rlabel metal3 s 31200 4768 32000 4888 6 wbs_a_sel_i[3]
port 208 nsew signal input
rlabel metal3 s 31200 1504 32000 1624 6 wbs_a_stb_i
port 209 nsew signal input
rlabel metal3 s 31200 2456 32000 2576 6 wbs_a_we_i
port 210 nsew signal input
rlabel metal3 s 31200 42848 32000 42968 6 wbs_b_ack_o
port 211 nsew signal output
rlabel metal3 s 31200 45296 32000 45416 6 wbs_b_adr_i[0]
port 212 nsew signal input
rlabel metal3 s 31200 45704 32000 45824 6 wbs_b_adr_i[1]
port 213 nsew signal input
rlabel metal3 s 31200 46112 32000 46232 6 wbs_b_adr_i[2]
port 214 nsew signal input
rlabel metal3 s 31200 46656 32000 46776 6 wbs_b_adr_i[3]
port 215 nsew signal input
rlabel metal3 s 31200 47064 32000 47184 6 wbs_b_adr_i[4]
port 216 nsew signal input
rlabel metal3 s 31200 47608 32000 47728 6 wbs_b_adr_i[5]
port 217 nsew signal input
rlabel metal3 s 31200 48016 32000 48136 6 wbs_b_adr_i[6]
port 218 nsew signal input
rlabel metal3 s 31200 48560 32000 48680 6 wbs_b_adr_i[7]
port 219 nsew signal input
rlabel metal3 s 31200 48968 32000 49088 6 wbs_b_adr_i[8]
port 220 nsew signal input
rlabel metal3 s 31200 49512 32000 49632 6 wbs_b_adr_i[9]
port 221 nsew signal input
rlabel metal3 s 31200 41896 32000 42016 6 wbs_b_cyc_i
port 222 nsew signal input
rlabel metal3 s 31200 49920 32000 50040 6 wbs_b_dat_i[0]
port 223 nsew signal input
rlabel metal3 s 31200 54680 32000 54800 6 wbs_b_dat_i[10]
port 224 nsew signal input
rlabel metal3 s 31200 55088 32000 55208 6 wbs_b_dat_i[11]
port 225 nsew signal input
rlabel metal3 s 31200 55632 32000 55752 6 wbs_b_dat_i[12]
port 226 nsew signal input
rlabel metal3 s 31200 56040 32000 56160 6 wbs_b_dat_i[13]
port 227 nsew signal input
rlabel metal3 s 31200 56584 32000 56704 6 wbs_b_dat_i[14]
port 228 nsew signal input
rlabel metal3 s 31200 56992 32000 57112 6 wbs_b_dat_i[15]
port 229 nsew signal input
rlabel metal3 s 31200 57400 32000 57520 6 wbs_b_dat_i[16]
port 230 nsew signal input
rlabel metal3 s 31200 57944 32000 58064 6 wbs_b_dat_i[17]
port 231 nsew signal input
rlabel metal3 s 31200 58352 32000 58472 6 wbs_b_dat_i[18]
port 232 nsew signal input
rlabel metal3 s 31200 58896 32000 59016 6 wbs_b_dat_i[19]
port 233 nsew signal input
rlabel metal3 s 31200 50464 32000 50584 6 wbs_b_dat_i[1]
port 234 nsew signal input
rlabel metal3 s 31200 59304 32000 59424 6 wbs_b_dat_i[20]
port 235 nsew signal input
rlabel metal3 s 31200 59848 32000 59968 6 wbs_b_dat_i[21]
port 236 nsew signal input
rlabel metal3 s 31200 60256 32000 60376 6 wbs_b_dat_i[22]
port 237 nsew signal input
rlabel metal3 s 31200 60800 32000 60920 6 wbs_b_dat_i[23]
port 238 nsew signal input
rlabel metal3 s 31200 61208 32000 61328 6 wbs_b_dat_i[24]
port 239 nsew signal input
rlabel metal3 s 31200 61752 32000 61872 6 wbs_b_dat_i[25]
port 240 nsew signal input
rlabel metal3 s 31200 62160 32000 62280 6 wbs_b_dat_i[26]
port 241 nsew signal input
rlabel metal3 s 31200 62704 32000 62824 6 wbs_b_dat_i[27]
port 242 nsew signal input
rlabel metal3 s 31200 63112 32000 63232 6 wbs_b_dat_i[28]
port 243 nsew signal input
rlabel metal3 s 31200 63520 32000 63640 6 wbs_b_dat_i[29]
port 244 nsew signal input
rlabel metal3 s 31200 50872 32000 50992 6 wbs_b_dat_i[2]
port 245 nsew signal input
rlabel metal3 s 31200 64064 32000 64184 6 wbs_b_dat_i[30]
port 246 nsew signal input
rlabel metal3 s 31200 64472 32000 64592 6 wbs_b_dat_i[31]
port 247 nsew signal input
rlabel metal3 s 31200 51416 32000 51536 6 wbs_b_dat_i[3]
port 248 nsew signal input
rlabel metal3 s 31200 51824 32000 51944 6 wbs_b_dat_i[4]
port 249 nsew signal input
rlabel metal3 s 31200 52232 32000 52352 6 wbs_b_dat_i[5]
port 250 nsew signal input
rlabel metal3 s 31200 52776 32000 52896 6 wbs_b_dat_i[6]
port 251 nsew signal input
rlabel metal3 s 31200 53184 32000 53304 6 wbs_b_dat_i[7]
port 252 nsew signal input
rlabel metal3 s 31200 53728 32000 53848 6 wbs_b_dat_i[8]
port 253 nsew signal input
rlabel metal3 s 31200 54136 32000 54256 6 wbs_b_dat_i[9]
port 254 nsew signal input
rlabel metal3 s 31200 65016 32000 65136 6 wbs_b_dat_o[0]
port 255 nsew signal output
rlabel metal3 s 31200 69640 32000 69760 6 wbs_b_dat_o[10]
port 256 nsew signal output
rlabel metal3 s 31200 70184 32000 70304 6 wbs_b_dat_o[11]
port 257 nsew signal output
rlabel metal3 s 31200 70592 32000 70712 6 wbs_b_dat_o[12]
port 258 nsew signal output
rlabel metal3 s 31200 71136 32000 71256 6 wbs_b_dat_o[13]
port 259 nsew signal output
rlabel metal3 s 31200 71544 32000 71664 6 wbs_b_dat_o[14]
port 260 nsew signal output
rlabel metal3 s 31200 72088 32000 72208 6 wbs_b_dat_o[15]
port 261 nsew signal output
rlabel metal3 s 31200 72496 32000 72616 6 wbs_b_dat_o[16]
port 262 nsew signal output
rlabel metal3 s 31200 73040 32000 73160 6 wbs_b_dat_o[17]
port 263 nsew signal output
rlabel metal3 s 31200 73448 32000 73568 6 wbs_b_dat_o[18]
port 264 nsew signal output
rlabel metal3 s 31200 73992 32000 74112 6 wbs_b_dat_o[19]
port 265 nsew signal output
rlabel metal3 s 31200 65424 32000 65544 6 wbs_b_dat_o[1]
port 266 nsew signal output
rlabel metal3 s 31200 74400 32000 74520 6 wbs_b_dat_o[20]
port 267 nsew signal output
rlabel metal3 s 31200 74808 32000 74928 6 wbs_b_dat_o[21]
port 268 nsew signal output
rlabel metal3 s 31200 75352 32000 75472 6 wbs_b_dat_o[22]
port 269 nsew signal output
rlabel metal3 s 31200 75760 32000 75880 6 wbs_b_dat_o[23]
port 270 nsew signal output
rlabel metal3 s 31200 76304 32000 76424 6 wbs_b_dat_o[24]
port 271 nsew signal output
rlabel metal3 s 31200 76712 32000 76832 6 wbs_b_dat_o[25]
port 272 nsew signal output
rlabel metal3 s 31200 77256 32000 77376 6 wbs_b_dat_o[26]
port 273 nsew signal output
rlabel metal3 s 31200 77664 32000 77784 6 wbs_b_dat_o[27]
port 274 nsew signal output
rlabel metal3 s 31200 78208 32000 78328 6 wbs_b_dat_o[28]
port 275 nsew signal output
rlabel metal3 s 31200 78616 32000 78736 6 wbs_b_dat_o[29]
port 276 nsew signal output
rlabel metal3 s 31200 65968 32000 66088 6 wbs_b_dat_o[2]
port 277 nsew signal output
rlabel metal3 s 31200 79160 32000 79280 6 wbs_b_dat_o[30]
port 278 nsew signal output
rlabel metal3 s 31200 79568 32000 79688 6 wbs_b_dat_o[31]
port 279 nsew signal output
rlabel metal3 s 31200 66376 32000 66496 6 wbs_b_dat_o[3]
port 280 nsew signal output
rlabel metal3 s 31200 66920 32000 67040 6 wbs_b_dat_o[4]
port 281 nsew signal output
rlabel metal3 s 31200 67328 32000 67448 6 wbs_b_dat_o[5]
port 282 nsew signal output
rlabel metal3 s 31200 67872 32000 67992 6 wbs_b_dat_o[6]
port 283 nsew signal output
rlabel metal3 s 31200 68280 32000 68400 6 wbs_b_dat_o[7]
port 284 nsew signal output
rlabel metal3 s 31200 68688 32000 68808 6 wbs_b_dat_o[8]
port 285 nsew signal output
rlabel metal3 s 31200 69232 32000 69352 6 wbs_b_dat_o[9]
port 286 nsew signal output
rlabel metal3 s 31200 43392 32000 43512 6 wbs_b_sel_i[0]
port 287 nsew signal input
rlabel metal3 s 31200 43800 32000 43920 6 wbs_b_sel_i[1]
port 288 nsew signal input
rlabel metal3 s 31200 44344 32000 44464 6 wbs_b_sel_i[2]
port 289 nsew signal input
rlabel metal3 s 31200 44752 32000 44872 6 wbs_b_sel_i[3]
port 290 nsew signal input
rlabel metal3 s 31200 41488 32000 41608 6 wbs_b_stb_i
port 291 nsew signal input
rlabel metal3 s 31200 42440 32000 42560 6 wbs_b_we_i
port 292 nsew signal input
rlabel metal3 s 31200 144 32000 264 6 writable_port_req
port 293 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4869946
string GDS_FILE /openlane/designs/wb_openram_wrapper/runs/RUN_2022.03.17_23.07.07/results/finishing/wb_openram_wrapper.magic.gds
string GDS_START 387950
<< end >>

