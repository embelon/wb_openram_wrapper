magic
tech sky130A
magscale 1 2
timestamp 1640039935
<< locali >>
rect 10885 74783 10919 74953
rect 10977 74919 11011 75701
rect 11069 74987 11103 76993
rect 11161 74919 11195 77469
rect 11069 74885 11195 74919
rect 10885 74749 11011 74783
rect 10977 73899 11011 74749
rect 10977 69207 11011 73729
rect 11069 72743 11103 74885
rect 11069 69547 11103 71553
rect 11161 71111 11195 74817
rect 9597 67167 9631 67337
rect 8493 64855 8527 64957
rect 10977 63835 11011 65705
rect 11069 63903 11103 69377
rect 11161 65127 11195 70941
rect 11253 70907 11287 76381
rect 11529 74239 11563 77537
rect 11253 67303 11287 69513
rect 10977 63801 11103 63835
rect 10977 56695 11011 63733
rect 11069 62407 11103 63801
rect 11161 62815 11195 64005
rect 11253 62815 11287 64957
rect 11069 60911 11103 62237
rect 11161 60979 11195 62781
rect 11253 60911 11287 62645
rect 11345 61047 11379 72029
rect 11437 70397 11471 71077
rect 11437 70363 11563 70397
rect 11437 60979 11471 67065
rect 11529 66011 11563 70363
rect 11621 68255 11655 72641
rect 11713 69479 11747 75293
rect 11253 60877 11379 60911
rect 10885 51323 10919 51561
rect 10977 51391 11011 52445
rect 11069 51391 11103 60605
rect 11161 60163 11195 60809
rect 11161 55199 11195 59993
rect 11161 51459 11195 55029
rect 11253 51527 11287 60741
rect 11345 59143 11379 60877
rect 11345 51391 11379 58973
rect 11437 53091 11471 60809
rect 11529 60299 11563 63189
rect 11621 60843 11655 68085
rect 11805 60843 11839 73185
rect 11897 62951 11931 68221
rect 11529 56083 11563 60129
rect 11621 55879 11655 60673
rect 11713 56967 11747 59109
rect 11805 55879 11839 60673
rect 11161 51357 11379 51391
rect 10885 51289 11011 51323
rect 10977 51077 11011 51289
rect 10885 51043 11011 51077
rect 10885 50711 10919 51043
rect 10977 49351 11011 50881
rect 10977 47243 11011 49113
rect 8953 43639 8987 43877
rect 10885 43639 10919 43945
rect 10977 41939 11011 47073
rect 10977 41259 11011 41565
rect 10919 41225 11011 41259
rect 9137 33303 9171 33473
rect 10977 32147 11011 41089
rect 11069 41055 11103 51017
rect 11161 50711 11195 51357
rect 11437 51051 11471 51425
rect 11529 51323 11563 55573
rect 11621 51323 11655 54553
rect 11161 47107 11195 49793
rect 11161 43843 11195 46937
rect 11069 40647 11103 40885
rect 11161 40715 11195 43673
rect 11253 42007 11287 50609
rect 11345 41531 11379 50949
rect 11529 50919 11563 51153
rect 11437 50885 11563 50919
rect 11437 47855 11471 50885
rect 11621 50779 11655 51153
rect 11713 50983 11747 55709
rect 11805 51391 11839 54009
rect 11897 53159 11931 61693
rect 11437 44455 11471 47685
rect 11253 41497 11379 41531
rect 11069 40613 11195 40647
rect 11069 32691 11103 40545
rect 11161 36839 11195 40613
rect 11161 35547 11195 36669
rect 10977 32113 11069 32147
rect 11161 32079 11195 33337
rect 10977 32045 11195 32079
rect 10977 32011 11011 32045
rect 10919 31977 11011 32011
rect 11069 31943 11103 31977
rect 10977 31909 11103 31943
rect 10977 26367 11011 31909
rect 11161 31807 11195 31909
rect 11069 31773 11195 31807
rect 10977 25279 11011 26197
rect 11069 22219 11103 31773
rect 11161 22627 11195 31569
rect 11253 24191 11287 41497
rect 11437 41259 11471 43741
rect 11529 41871 11563 50473
rect 11621 47991 11655 50609
rect 11345 33303 11379 41021
rect 11437 32895 11471 40069
rect 11345 30923 11379 32793
rect 11345 22219 11379 30753
rect 11437 22695 11471 32725
rect 11069 22185 11195 22219
rect 11345 22185 11471 22219
rect 11161 22097 11195 22185
rect 11069 22063 11195 22097
rect 9229 17187 9263 17289
rect 10977 8755 11011 21981
rect 11069 12437 11103 22063
rect 11345 21947 11379 22117
rect 11437 21947 11471 22185
rect 11529 22083 11563 41701
rect 11621 22287 11655 47821
rect 11713 41735 11747 50337
rect 11805 41939 11839 50677
rect 11897 41803 11931 52989
rect 11713 41701 11931 41735
rect 11713 31943 11747 41089
rect 11621 22015 11655 22117
rect 11529 21981 11655 22015
rect 11161 20995 11195 21913
rect 11529 21879 11563 21981
rect 11161 18819 11195 20825
rect 11161 18785 11287 18819
rect 11161 16303 11195 18717
rect 11253 17119 11287 18785
rect 11345 17391 11379 21777
rect 11161 13447 11195 16133
rect 11253 15487 11287 16541
rect 11069 12403 11195 12437
rect 10977 8721 11103 8755
rect 10977 6783 11011 8517
rect 11069 7531 11103 8721
rect 11161 5355 11195 12403
rect 11345 8075 11379 17221
rect 11437 8415 11471 21777
rect 11529 9027 11563 21709
rect 11621 18683 11655 21709
rect 11621 17187 11655 17357
rect 11713 17255 11747 31773
rect 11805 31671 11839 41633
rect 11897 40647 11931 41701
rect 11897 33371 11931 40477
rect 11897 31331 11931 32657
rect 11621 17153 11747 17187
rect 11621 10183 11655 17085
rect 11713 9163 11747 17153
rect 11805 8619 11839 31297
rect 11897 22763 11931 29665
rect 11897 13311 11931 21913
<< viali >>
rect 7573 77673 7607 77707
rect 8309 77673 8343 77707
rect 1409 77537 1443 77571
rect 1685 77537 1719 77571
rect 11529 77537 11563 77571
rect 2881 77469 2915 77503
rect 7389 77469 7423 77503
rect 8125 77469 8159 77503
rect 9137 77469 9171 77503
rect 9873 77469 9907 77503
rect 11161 77469 11195 77503
rect 2697 77333 2731 77367
rect 9321 77333 9355 77367
rect 10057 77333 10091 77367
rect 1409 77129 1443 77163
rect 8585 77129 8619 77163
rect 9321 77129 9355 77163
rect 1593 76993 1627 77027
rect 2237 76993 2271 77027
rect 2881 76993 2915 77027
rect 8401 76993 8435 77027
rect 9137 76993 9171 77027
rect 9873 76993 9907 77027
rect 11069 76993 11103 77027
rect 2053 76857 2087 76891
rect 2697 76789 2731 76823
rect 10057 76789 10091 76823
rect 9321 76585 9355 76619
rect 1593 76381 1627 76415
rect 9137 76381 9171 76415
rect 9873 76381 9907 76415
rect 1409 76245 1443 76279
rect 10057 76245 10091 76279
rect 9321 76041 9355 76075
rect 1685 75905 1719 75939
rect 9137 75905 9171 75939
rect 9873 75905 9907 75939
rect 1409 75837 1443 75871
rect 10057 75701 10091 75735
rect 10977 75701 11011 75735
rect 9873 75293 9907 75327
rect 1869 75225 1903 75259
rect 1961 75157 1995 75191
rect 10057 75157 10091 75191
rect 2697 74953 2731 74987
rect 3065 74953 3099 74987
rect 10885 74953 10919 74987
rect 1593 74817 1627 74851
rect 2237 74817 2271 74851
rect 9873 74817 9907 74851
rect 11069 74953 11103 74987
rect 10977 74885 11011 74919
rect 11253 76381 11287 76415
rect 3157 74749 3191 74783
rect 3249 74749 3283 74783
rect 1409 74681 1443 74715
rect 2053 74613 2087 74647
rect 10057 74613 10091 74647
rect 6101 74409 6135 74443
rect 9413 74409 9447 74443
rect 1961 74341 1995 74375
rect 2513 74273 2547 74307
rect 6745 74273 6779 74307
rect 10057 74273 10091 74307
rect 2421 74205 2455 74239
rect 9781 74205 9815 74239
rect 6469 74137 6503 74171
rect 2329 74069 2363 74103
rect 6561 74069 6595 74103
rect 9873 74069 9907 74103
rect 1593 73865 1627 73899
rect 3341 73865 3375 73899
rect 10977 73865 11011 73899
rect 1961 73729 1995 73763
rect 3709 73729 3743 73763
rect 3801 73729 3835 73763
rect 9137 73729 9171 73763
rect 9873 73729 9907 73763
rect 10977 73729 11011 73763
rect 2053 73661 2087 73695
rect 2237 73661 2271 73695
rect 3985 73661 4019 73695
rect 9321 73525 9355 73559
rect 10057 73525 10091 73559
rect 2145 73185 2179 73219
rect 7665 73185 7699 73219
rect 9965 73185 9999 73219
rect 1961 73117 1995 73151
rect 2881 73117 2915 73151
rect 10057 73117 10091 73151
rect 7573 73049 7607 73083
rect 9965 73049 9999 73083
rect 1501 72981 1535 73015
rect 1869 72981 1903 73015
rect 2697 72981 2731 73015
rect 7113 72981 7147 73015
rect 7481 72981 7515 73015
rect 9487 72981 9521 73015
rect 1777 72777 1811 72811
rect 2605 72777 2639 72811
rect 2973 72641 3007 72675
rect 9137 72641 9171 72675
rect 9873 72641 9907 72675
rect 1869 72573 1903 72607
rect 2053 72573 2087 72607
rect 3065 72573 3099 72607
rect 3157 72573 3191 72607
rect 1409 72505 1443 72539
rect 9321 72505 9355 72539
rect 10057 72437 10091 72471
rect 1409 72165 1443 72199
rect 6193 72165 6227 72199
rect 1593 72029 1627 72063
rect 2237 72029 2271 72063
rect 4077 72029 4111 72063
rect 4169 72029 4203 72063
rect 4353 72029 4387 72063
rect 6745 72029 6779 72063
rect 9137 72029 9171 72063
rect 9781 72029 9815 72063
rect 9873 72029 9907 72063
rect 4813 71961 4847 71995
rect 6469 71961 6503 71995
rect 6653 71961 6687 71995
rect 2053 71893 2087 71927
rect 9321 71893 9355 71927
rect 10057 71893 10091 71927
rect 1593 71553 1627 71587
rect 9873 71553 9907 71587
rect 1409 71349 1443 71383
rect 10057 71349 10091 71383
rect 1685 71009 1719 71043
rect 4445 71009 4479 71043
rect 1409 70941 1443 70975
rect 4169 70941 4203 70975
rect 9873 70941 9907 70975
rect 3801 70805 3835 70839
rect 4261 70805 4295 70839
rect 10057 70805 10091 70839
rect 2237 70465 2271 70499
rect 2329 70465 2363 70499
rect 2513 70465 2547 70499
rect 7481 70465 7515 70499
rect 7665 70465 7699 70499
rect 2973 70397 3007 70431
rect 7389 70397 7423 70431
rect 8125 70397 8159 70431
rect 9321 70397 9355 70431
rect 10241 70397 10275 70431
rect 9413 70057 9447 70091
rect 2881 69989 2915 70023
rect 10057 69921 10091 69955
rect 1685 69853 1719 69887
rect 1777 69853 1811 69887
rect 1961 69853 1995 69887
rect 3065 69853 3099 69887
rect 3985 69853 4019 69887
rect 2421 69785 2455 69819
rect 9781 69785 9815 69819
rect 3801 69717 3835 69751
rect 9229 69717 9263 69751
rect 9873 69717 9907 69751
rect 1501 69513 1535 69547
rect 1869 69513 1903 69547
rect 9229 69513 9263 69547
rect 10425 69513 10459 69547
rect 3065 69377 3099 69411
rect 3249 69377 3283 69411
rect 8401 69377 8435 69411
rect 9045 69377 9079 69411
rect 9781 69377 9815 69411
rect 10241 69377 10275 69411
rect 1961 69309 1995 69343
rect 2145 69309 2179 69343
rect 2973 69309 3007 69343
rect 3709 69309 3743 69343
rect 9873 69309 9907 69343
rect 10057 69309 10091 69343
rect 8585 69241 8619 69275
rect 11069 72709 11103 72743
rect 11161 74817 11195 74851
rect 11069 71553 11103 71587
rect 11161 71077 11195 71111
rect 11069 69513 11103 69547
rect 11161 70941 11195 70975
rect 9413 69173 9447 69207
rect 10977 69173 11011 69207
rect 11069 69377 11103 69411
rect 6837 68969 6871 69003
rect 2513 68833 2547 68867
rect 7481 68833 7515 68867
rect 1593 68765 1627 68799
rect 2605 68765 2639 68799
rect 2789 68765 2823 68799
rect 7205 68765 7239 68799
rect 8125 68765 8159 68799
rect 3249 68697 3283 68731
rect 7297 68697 7331 68731
rect 1409 68629 1443 68663
rect 8309 68629 8343 68663
rect 9229 68629 9263 68663
rect 10241 68629 10275 68663
rect 9965 68425 9999 68459
rect 9781 68357 9815 68391
rect 10057 68357 10091 68391
rect 1593 68289 1627 68323
rect 3525 68289 3559 68323
rect 3617 68289 3651 68323
rect 3801 68289 3835 68323
rect 8585 68289 8619 68323
rect 4261 68221 4295 68255
rect 1409 68085 1443 68119
rect 8769 68085 8803 68119
rect 9137 68085 9171 68119
rect 9505 68085 9539 68119
rect 9413 67813 9447 67847
rect 9965 67745 9999 67779
rect 1409 67677 1443 67711
rect 1685 67677 1719 67711
rect 8125 67677 8159 67711
rect 9689 67609 9723 67643
rect 9873 67609 9907 67643
rect 8309 67541 8343 67575
rect 1777 67337 1811 67371
rect 8677 67337 8711 67371
rect 9597 67337 9631 67371
rect 2789 67201 2823 67235
rect 8309 67201 8343 67235
rect 9045 67201 9079 67235
rect 9873 67201 9907 67235
rect 1869 67133 1903 67167
rect 2053 67133 2087 67167
rect 9137 67133 9171 67167
rect 9321 67133 9355 67167
rect 9597 67133 9631 67167
rect 1409 67065 1443 67099
rect 8493 67065 8527 67099
rect 9781 67065 9815 67099
rect 2605 66997 2639 67031
rect 10057 66997 10091 67031
rect 2053 66657 2087 66691
rect 2145 66589 2179 66623
rect 2329 66589 2363 66623
rect 7113 66589 7147 66623
rect 7205 66589 7239 66623
rect 7389 66589 7423 66623
rect 9413 66589 9447 66623
rect 9505 66589 9539 66623
rect 9689 66589 9723 66623
rect 2789 66521 2823 66555
rect 7849 66521 7883 66555
rect 10149 66521 10183 66555
rect 2421 66181 2455 66215
rect 3249 66181 3283 66215
rect 1777 66113 1811 66147
rect 1961 66113 1995 66147
rect 9137 66113 9171 66147
rect 9873 66113 9907 66147
rect 1685 66045 1719 66079
rect 3341 66045 3375 66079
rect 3525 66045 3559 66079
rect 2881 65909 2915 65943
rect 9321 65909 9355 65943
rect 10057 65909 10091 65943
rect 10977 65705 11011 65739
rect 1409 65637 1443 65671
rect 1593 65501 1627 65535
rect 2237 65501 2271 65535
rect 9413 65501 9447 65535
rect 9505 65501 9539 65535
rect 9689 65501 9723 65535
rect 10149 65433 10183 65467
rect 2053 65365 2087 65399
rect 7297 65161 7331 65195
rect 7665 65161 7699 65195
rect 8585 65161 8619 65195
rect 1869 65025 1903 65059
rect 7757 65025 7791 65059
rect 8769 65025 8803 65059
rect 9413 65025 9447 65059
rect 9873 65025 9907 65059
rect 7849 64957 7883 64991
rect 8493 64957 8527 64991
rect 10057 64889 10091 64923
rect 1961 64821 1995 64855
rect 8493 64821 8527 64855
rect 9229 64821 9263 64855
rect 1409 64413 1443 64447
rect 9413 64413 9447 64447
rect 9505 64413 9539 64447
rect 9689 64413 9723 64447
rect 10149 64345 10183 64379
rect 1593 64277 1627 64311
rect 9137 64073 9171 64107
rect 9229 64005 9263 64039
rect 1409 63937 1443 63971
rect 10149 63937 10183 63971
rect 9413 63869 9447 63903
rect 11529 74205 11563 74239
rect 11713 75293 11747 75327
rect 11621 72641 11655 72675
rect 11253 70873 11287 70907
rect 11345 72029 11379 72063
rect 11253 69513 11287 69547
rect 11253 67269 11287 67303
rect 11161 65093 11195 65127
rect 11253 64957 11287 64991
rect 11069 63869 11103 63903
rect 11161 64005 11195 64039
rect 8769 63801 8803 63835
rect 1593 63733 1627 63767
rect 9965 63733 9999 63767
rect 10977 63733 11011 63767
rect 2605 63461 2639 63495
rect 2973 63393 3007 63427
rect 3157 63393 3191 63427
rect 1409 63325 1443 63359
rect 9505 63325 9539 63359
rect 10149 63325 10183 63359
rect 1593 63189 1627 63223
rect 3065 63189 3099 63223
rect 9321 63189 9355 63223
rect 9965 63189 9999 63223
rect 2329 62985 2363 63019
rect 7849 62985 7883 63019
rect 9321 62985 9355 63019
rect 9413 62849 9447 62883
rect 10149 62849 10183 62883
rect 2421 62781 2455 62815
rect 2513 62781 2547 62815
rect 7849 62781 7883 62815
rect 7941 62781 7975 62815
rect 9321 62781 9355 62815
rect 1961 62713 1995 62747
rect 7389 62645 7423 62679
rect 8861 62645 8895 62679
rect 9965 62645 9999 62679
rect 7665 62441 7699 62475
rect 8309 62305 8343 62339
rect 8033 62237 8067 62271
rect 9321 62237 9355 62271
rect 9597 62237 9631 62271
rect 1869 62169 1903 62203
rect 2053 62169 2087 62203
rect 8125 62101 8159 62135
rect 1869 61761 1903 61795
rect 9321 61693 9355 61727
rect 9597 61693 9631 61727
rect 2053 61625 2087 61659
rect 2237 61217 2271 61251
rect 2329 61149 2363 61183
rect 2513 61149 2547 61183
rect 9413 61149 9447 61183
rect 9505 61149 9539 61183
rect 9689 61149 9723 61183
rect 2973 61081 3007 61115
rect 10149 61081 10183 61115
rect 2053 60809 2087 60843
rect 2145 60741 2179 60775
rect 8677 60741 8711 60775
rect 2789 60673 2823 60707
rect 9321 60673 9355 60707
rect 2053 60605 2087 60639
rect 9597 60605 9631 60639
rect 2973 60537 3007 60571
rect 1593 60469 1627 60503
rect 8769 60469 8803 60503
rect 7757 60197 7791 60231
rect 8217 60129 8251 60163
rect 8309 60129 8343 60163
rect 9965 60061 9999 60095
rect 1869 59993 1903 60027
rect 10149 59993 10183 60027
rect 1961 59925 1995 59959
rect 8217 59925 8251 59959
rect 9229 59653 9263 59687
rect 1869 59585 1903 59619
rect 9965 59585 9999 59619
rect 10149 59449 10183 59483
rect 1961 59381 1995 59415
rect 9321 59381 9355 59415
rect 10149 58973 10183 59007
rect 9965 58905 9999 58939
rect 1409 58497 1443 58531
rect 9965 58497 9999 58531
rect 1593 58361 1627 58395
rect 10149 58361 10183 58395
rect 1409 57885 1443 57919
rect 9965 57817 9999 57851
rect 1593 57749 1627 57783
rect 9781 57749 9815 57783
rect 10057 57749 10091 57783
rect 1409 57409 1443 57443
rect 9229 57409 9263 57443
rect 9873 57409 9907 57443
rect 1593 57205 1627 57239
rect 9321 57205 9355 57239
rect 10057 57205 10091 57239
rect 9505 56933 9539 56967
rect 9965 56865 9999 56899
rect 1409 56797 1443 56831
rect 10057 56729 10091 56763
rect 11069 62373 11103 62407
rect 11161 62781 11195 62815
rect 11253 62781 11287 62815
rect 11069 62237 11103 62271
rect 11161 60945 11195 60979
rect 11253 62645 11287 62679
rect 11069 60877 11103 60911
rect 11437 71077 11471 71111
rect 11345 61013 11379 61047
rect 11437 67065 11471 67099
rect 11713 69445 11747 69479
rect 11805 73185 11839 73219
rect 11621 68221 11655 68255
rect 11529 65977 11563 66011
rect 11621 68085 11655 68119
rect 11437 60945 11471 60979
rect 11529 63189 11563 63223
rect 11161 60809 11195 60843
rect 1593 56661 1627 56695
rect 9965 56661 9999 56695
rect 10977 56661 11011 56695
rect 11069 60605 11103 60639
rect 1409 56321 1443 56355
rect 9873 56321 9907 56355
rect 1593 56117 1627 56151
rect 10057 56117 10091 56151
rect 1409 55709 1443 55743
rect 9873 55709 9907 55743
rect 1593 55573 1627 55607
rect 9781 55573 9815 55607
rect 10057 55573 10091 55607
rect 1409 55233 1443 55267
rect 9873 55233 9907 55267
rect 1593 55029 1627 55063
rect 10057 55029 10091 55063
rect 1685 54825 1719 54859
rect 2145 54689 2179 54723
rect 2237 54553 2271 54587
rect 9965 54553 9999 54587
rect 10149 54553 10183 54587
rect 2145 54485 2179 54519
rect 2421 54281 2455 54315
rect 2237 54145 2271 54179
rect 9137 54145 9171 54179
rect 9873 54145 9907 54179
rect 2513 54077 2547 54111
rect 9781 54009 9815 54043
rect 10057 54009 10091 54043
rect 1961 53941 1995 53975
rect 9321 53941 9355 53975
rect 1593 53737 1627 53771
rect 1409 53533 1443 53567
rect 9137 53533 9171 53567
rect 9873 53533 9907 53567
rect 9321 53397 9355 53431
rect 9781 53397 9815 53431
rect 10057 53397 10091 53431
rect 1593 53193 1627 53227
rect 9965 53193 9999 53227
rect 1409 53057 1443 53091
rect 9781 53057 9815 53091
rect 10057 52989 10091 53023
rect 9505 52853 9539 52887
rect 1685 52649 1719 52683
rect 2789 52581 2823 52615
rect 9321 52581 9355 52615
rect 1961 52445 1995 52479
rect 2237 52445 2271 52479
rect 2973 52445 3007 52479
rect 9137 52445 9171 52479
rect 9873 52445 9907 52479
rect 10977 52445 11011 52479
rect 2145 52377 2179 52411
rect 9781 52309 9815 52343
rect 10057 52309 10091 52343
rect 1961 52105 1995 52139
rect 1869 51969 1903 52003
rect 9137 51969 9171 52003
rect 9873 51969 9907 52003
rect 9321 51765 9355 51799
rect 10057 51765 10091 51799
rect 1593 51561 1627 51595
rect 8953 51561 8987 51595
rect 10885 51561 10919 51595
rect 9505 51425 9539 51459
rect 1409 51357 1443 51391
rect 10977 51357 11011 51391
rect 11161 60129 11195 60163
rect 11253 60741 11287 60775
rect 11161 59993 11195 60027
rect 11161 55165 11195 55199
rect 11161 55029 11195 55063
rect 11345 59109 11379 59143
rect 11437 60809 11471 60843
rect 11253 51493 11287 51527
rect 11345 58973 11379 59007
rect 11161 51425 11195 51459
rect 11621 60809 11655 60843
rect 11897 68221 11931 68255
rect 11897 62917 11931 62951
rect 11805 60809 11839 60843
rect 11897 61693 11931 61727
rect 11529 60265 11563 60299
rect 11621 60673 11655 60707
rect 11529 60129 11563 60163
rect 11529 56049 11563 56083
rect 11805 60673 11839 60707
rect 11713 59109 11747 59143
rect 11713 56933 11747 56967
rect 11621 55845 11655 55879
rect 11805 55845 11839 55879
rect 11713 55709 11747 55743
rect 11437 53057 11471 53091
rect 11529 55573 11563 55607
rect 11069 51357 11103 51391
rect 11437 51425 11471 51459
rect 9321 51289 9355 51323
rect 9413 51221 9447 51255
rect 1961 51017 1995 51051
rect 2513 51017 2547 51051
rect 8769 51017 8803 51051
rect 1869 50881 1903 50915
rect 2697 50881 2731 50915
rect 9137 50881 9171 50915
rect 10149 50881 10183 50915
rect 9229 50813 9263 50847
rect 9413 50813 9447 50847
rect 11069 51017 11103 51051
rect 9965 50677 9999 50711
rect 10885 50677 10919 50711
rect 10977 50881 11011 50915
rect 1961 50473 1995 50507
rect 9137 50473 9171 50507
rect 9781 50337 9815 50371
rect 8125 50269 8159 50303
rect 1869 50201 1903 50235
rect 8309 50133 8343 50167
rect 9505 50133 9539 50167
rect 9597 50133 9631 50167
rect 8861 49929 8895 49963
rect 9965 49929 9999 49963
rect 8677 49793 8711 49827
rect 10057 49793 10091 49827
rect 9965 49725 9999 49759
rect 9505 49657 9539 49691
rect 8217 49385 8251 49419
rect 2053 49317 2087 49351
rect 10977 49317 11011 49351
rect 9229 49249 9263 49283
rect 1869 49181 1903 49215
rect 8401 49181 8435 49215
rect 9321 49181 9355 49215
rect 9505 49181 9539 49215
rect 9965 49113 9999 49147
rect 10977 49113 11011 49147
rect 8125 48841 8159 48875
rect 2053 48773 2087 48807
rect 1869 48705 1903 48739
rect 8309 48705 8343 48739
rect 9137 48705 9171 48739
rect 9321 48705 9355 48739
rect 9045 48637 9079 48671
rect 9781 48637 9815 48671
rect 2053 48229 2087 48263
rect 8401 48093 8435 48127
rect 9321 48093 9355 48127
rect 9413 48093 9447 48127
rect 9597 48093 9631 48127
rect 1869 48025 1903 48059
rect 10057 48025 10091 48059
rect 8217 47957 8251 47991
rect 1961 47753 1995 47787
rect 4721 47753 4755 47787
rect 5089 47753 5123 47787
rect 9045 47753 9079 47787
rect 9689 47685 9723 47719
rect 1869 47617 1903 47651
rect 8861 47617 8895 47651
rect 9229 47617 9263 47651
rect 9781 47617 9815 47651
rect 10333 47617 10367 47651
rect 5181 47549 5215 47583
rect 5365 47549 5399 47583
rect 9965 47549 9999 47583
rect 9321 47481 9355 47515
rect 8677 47413 8711 47447
rect 10149 47413 10183 47447
rect 1961 47209 1995 47243
rect 9413 47209 9447 47243
rect 10977 47209 11011 47243
rect 8217 47141 8251 47175
rect 9965 47073 9999 47107
rect 10977 47073 11011 47107
rect 8401 47005 8435 47039
rect 1869 46937 1903 46971
rect 9781 46937 9815 46971
rect 9873 46869 9907 46903
rect 9413 46665 9447 46699
rect 9781 46665 9815 46699
rect 8677 46597 8711 46631
rect 5089 46529 5123 46563
rect 5273 46529 5307 46563
rect 8493 46529 8527 46563
rect 4997 46461 5031 46495
rect 5733 46461 5767 46495
rect 8769 46461 8803 46495
rect 9873 46461 9907 46495
rect 9965 46461 9999 46495
rect 8217 46393 8251 46427
rect 1961 46121 1995 46155
rect 9505 46053 9539 46087
rect 1869 45917 1903 45951
rect 9781 45849 9815 45883
rect 10057 45849 10091 45883
rect 9965 45781 9999 45815
rect 10333 45577 10367 45611
rect 3341 45509 3375 45543
rect 1409 45441 1443 45475
rect 3433 45441 3467 45475
rect 8677 45441 8711 45475
rect 3617 45373 3651 45407
rect 2973 45305 3007 45339
rect 9229 45305 9263 45339
rect 1593 45237 1627 45271
rect 8861 45237 8895 45271
rect 2053 44965 2087 44999
rect 9413 44829 9447 44863
rect 9505 44829 9539 44863
rect 9689 44829 9723 44863
rect 1869 44761 1903 44795
rect 10149 44761 10183 44795
rect 2053 44421 2087 44455
rect 1869 44353 1903 44387
rect 8401 44353 8435 44387
rect 9505 44353 9539 44387
rect 9689 44353 9723 44387
rect 9414 44285 9448 44319
rect 10149 44285 10183 44319
rect 8585 44149 8619 44183
rect 10885 43945 10919 43979
rect 8953 43877 8987 43911
rect 8217 43809 8251 43843
rect 4077 43741 4111 43775
rect 4169 43741 4203 43775
rect 4353 43741 4387 43775
rect 8033 43741 8067 43775
rect 4813 43673 4847 43707
rect 9413 43741 9447 43775
rect 9505 43741 9539 43775
rect 9689 43741 9723 43775
rect 10149 43673 10183 43707
rect 7665 43605 7699 43639
rect 8125 43605 8159 43639
rect 8953 43605 8987 43639
rect 10885 43605 10919 43639
rect 1961 43401 1995 43435
rect 9321 43401 9355 43435
rect 1869 43265 1903 43299
rect 8401 43265 8435 43299
rect 9137 43265 9171 43299
rect 9873 43265 9907 43299
rect 8585 43061 8619 43095
rect 9781 43061 9815 43095
rect 10057 43061 10091 43095
rect 6561 42789 6595 42823
rect 7113 42721 7147 42755
rect 9965 42721 9999 42755
rect 1409 42653 1443 42687
rect 9487 42653 9521 42687
rect 10057 42653 10091 42687
rect 6837 42585 6871 42619
rect 9137 42585 9171 42619
rect 9321 42585 9355 42619
rect 9965 42585 9999 42619
rect 1593 42517 1627 42551
rect 7021 42517 7055 42551
rect 10333 42517 10367 42551
rect 1593 42313 1627 42347
rect 5273 42245 5307 42279
rect 1409 42177 1443 42211
rect 5365 42177 5399 42211
rect 9137 42177 9171 42211
rect 9965 42177 9999 42211
rect 5181 42109 5215 42143
rect 4813 42041 4847 42075
rect 10149 42041 10183 42075
rect 9321 41973 9355 42007
rect 10977 41905 11011 41939
rect 1593 41769 1627 41803
rect 1409 41565 1443 41599
rect 10977 41565 11011 41599
rect 9965 41497 9999 41531
rect 10057 41429 10091 41463
rect 10885 41225 10919 41259
rect 2053 41157 2087 41191
rect 1869 41089 1903 41123
rect 9965 41089 9999 41123
rect 10977 41089 11011 41123
rect 10149 40953 10183 40987
rect 2053 40613 2087 40647
rect 9137 40477 9171 40511
rect 9873 40477 9907 40511
rect 1869 40409 1903 40443
rect 9321 40341 9355 40375
rect 10057 40341 10091 40375
rect 9495 40137 9529 40171
rect 6837 40069 6871 40103
rect 9965 40069 9999 40103
rect 1685 40001 1719 40035
rect 8493 40001 8527 40035
rect 9137 40001 9171 40035
rect 9321 40001 9355 40035
rect 1409 39933 1443 39967
rect 6929 39933 6963 39967
rect 7021 39933 7055 39967
rect 9965 39933 9999 39967
rect 10057 39933 10091 39967
rect 6469 39865 6503 39899
rect 8677 39797 8711 39831
rect 10333 39797 10367 39831
rect 1869 39593 1903 39627
rect 9229 39593 9263 39627
rect 2329 39457 2363 39491
rect 5273 39457 5307 39491
rect 5181 39389 5215 39423
rect 2421 39321 2455 39355
rect 9505 39321 9539 39355
rect 9781 39321 9815 39355
rect 2329 39253 2363 39287
rect 4721 39253 4755 39287
rect 5089 39253 5123 39287
rect 9689 39253 9723 39287
rect 1593 39049 1627 39083
rect 9597 38981 9631 39015
rect 9689 38981 9723 39015
rect 1409 38913 1443 38947
rect 8309 38913 8343 38947
rect 9505 38845 9539 38879
rect 9137 38777 9171 38811
rect 8493 38709 8527 38743
rect 1593 38505 1627 38539
rect 9045 38505 9079 38539
rect 9413 38369 9447 38403
rect 9597 38369 9631 38403
rect 1409 38301 1443 38335
rect 8125 38301 8159 38335
rect 8309 38165 8343 38199
rect 9505 38165 9539 38199
rect 9045 37961 9079 37995
rect 9505 37961 9539 37995
rect 1409 37825 1443 37859
rect 8309 37825 8343 37859
rect 9413 37825 9447 37859
rect 9597 37757 9631 37791
rect 1593 37689 1627 37723
rect 8493 37621 8527 37655
rect 2421 37281 2455 37315
rect 9689 37281 9723 37315
rect 2145 37213 2179 37247
rect 8125 37213 8159 37247
rect 9597 37213 9631 37247
rect 9505 37145 9539 37179
rect 1777 37077 1811 37111
rect 2237 37077 2271 37111
rect 8309 37077 8343 37111
rect 9137 37077 9171 37111
rect 9965 36873 9999 36907
rect 10057 36805 10091 36839
rect 7941 36737 7975 36771
rect 8677 36737 8711 36771
rect 1409 36669 1443 36703
rect 1685 36669 1719 36703
rect 9321 36669 9355 36703
rect 9965 36669 9999 36703
rect 8125 36601 8159 36635
rect 8861 36533 8895 36567
rect 9505 36533 9539 36567
rect 10333 36533 10367 36567
rect 1409 36329 1443 36363
rect 8953 36261 8987 36295
rect 2329 36193 2363 36227
rect 3065 36193 3099 36227
rect 9413 36193 9447 36227
rect 9597 36193 9631 36227
rect 1593 36125 1627 36159
rect 2421 36125 2455 36159
rect 2605 36125 2639 36159
rect 9321 35989 9355 36023
rect 1409 35785 1443 35819
rect 1593 35649 1627 35683
rect 9137 35649 9171 35683
rect 9873 35649 9907 35683
rect 9321 35445 9355 35479
rect 10057 35445 10091 35479
rect 1409 35241 1443 35275
rect 9321 35241 9355 35275
rect 2513 35105 2547 35139
rect 2605 35105 2639 35139
rect 1593 35037 1627 35071
rect 2421 35037 2455 35071
rect 9137 35037 9171 35071
rect 9873 35037 9907 35071
rect 2053 34901 2087 34935
rect 10057 34901 10091 34935
rect 9413 34697 9447 34731
rect 3157 34629 3191 34663
rect 9873 34629 9907 34663
rect 2513 34561 2547 34595
rect 2697 34561 2731 34595
rect 9781 34561 9815 34595
rect 2421 34493 2455 34527
rect 9229 34493 9263 34527
rect 10057 34493 10091 34527
rect 1685 34017 1719 34051
rect 1409 33949 1443 33983
rect 9137 33949 9171 33983
rect 9873 33949 9907 33983
rect 9321 33813 9355 33847
rect 10057 33813 10091 33847
rect 9413 33609 9447 33643
rect 9873 33609 9907 33643
rect 1685 33473 1719 33507
rect 8677 33473 8711 33507
rect 9137 33473 9171 33507
rect 9781 33473 9815 33507
rect 1409 33405 1443 33439
rect 8861 33337 8895 33371
rect 10057 33405 10091 33439
rect 9137 33269 9171 33303
rect 9229 33269 9263 33303
rect 1409 33065 1443 33099
rect 10425 33065 10459 33099
rect 9413 32997 9447 33031
rect 2697 32929 2731 32963
rect 10057 32929 10091 32963
rect 1593 32861 1627 32895
rect 2605 32861 2639 32895
rect 9045 32861 9079 32895
rect 9873 32861 9907 32895
rect 10241 32861 10275 32895
rect 2145 32725 2179 32759
rect 2513 32725 2547 32759
rect 9229 32725 9263 32759
rect 9781 32725 9815 32759
rect 1409 32521 1443 32555
rect 1593 32385 1627 32419
rect 8677 32385 8711 32419
rect 9321 32317 9355 32351
rect 10241 32249 10275 32283
rect 8861 32181 8895 32215
rect 11529 51289 11563 51323
rect 11621 54553 11655 54587
rect 11621 51289 11655 51323
rect 11437 51017 11471 51051
rect 11529 51153 11563 51187
rect 11161 50677 11195 50711
rect 11345 50949 11379 50983
rect 11253 50609 11287 50643
rect 11161 49793 11195 49827
rect 11161 47073 11195 47107
rect 11161 46937 11195 46971
rect 11161 43809 11195 43843
rect 11069 41021 11103 41055
rect 11161 43673 11195 43707
rect 11069 40885 11103 40919
rect 11253 41973 11287 42007
rect 11621 51153 11655 51187
rect 11805 54009 11839 54043
rect 11897 53125 11931 53159
rect 11805 51357 11839 51391
rect 11897 52989 11931 53023
rect 11713 50949 11747 50983
rect 11621 50745 11655 50779
rect 11805 50677 11839 50711
rect 11621 50609 11655 50643
rect 11437 47821 11471 47855
rect 11529 50473 11563 50507
rect 11437 47685 11471 47719
rect 11437 44421 11471 44455
rect 11161 40681 11195 40715
rect 11437 43741 11471 43775
rect 11069 40545 11103 40579
rect 11161 36805 11195 36839
rect 11161 36669 11195 36703
rect 11161 35513 11195 35547
rect 11069 32657 11103 32691
rect 11161 33337 11195 33371
rect 11069 32113 11103 32147
rect 1409 31977 1443 32011
rect 10885 31977 10919 32011
rect 11069 31977 11103 32011
rect 11161 31909 11195 31943
rect 1593 31773 1627 31807
rect 9321 31773 9355 31807
rect 10241 31773 10275 31807
rect 9873 31433 9907 31467
rect 9781 31297 9815 31331
rect 10266 31297 10300 31331
rect 10057 31229 10091 31263
rect 9413 31093 9447 31127
rect 10425 31093 10459 31127
rect 1409 30685 1443 30719
rect 9873 30685 9907 30719
rect 1593 30549 1627 30583
rect 10057 30549 10091 30583
rect 1409 30209 1443 30243
rect 9873 30209 9907 30243
rect 1593 30005 1627 30039
rect 10057 30005 10091 30039
rect 1409 29597 1443 29631
rect 9137 29597 9171 29631
rect 9873 29597 9907 29631
rect 1593 29461 1627 29495
rect 9321 29461 9355 29495
rect 10057 29461 10091 29495
rect 9413 29257 9447 29291
rect 9873 29257 9907 29291
rect 1409 29121 1443 29155
rect 8677 29121 8711 29155
rect 9781 29121 9815 29155
rect 9229 29053 9263 29087
rect 9965 29053 9999 29087
rect 1593 28985 1627 29019
rect 8861 28985 8895 29019
rect 1409 28509 1443 28543
rect 9137 28509 9171 28543
rect 9873 28509 9907 28543
rect 1593 28373 1627 28407
rect 9321 28373 9355 28407
rect 10057 28373 10091 28407
rect 9781 28169 9815 28203
rect 9873 28033 9907 28067
rect 10057 27829 10091 27863
rect 1409 27421 1443 27455
rect 9873 27421 9907 27455
rect 1593 27285 1627 27319
rect 10057 27285 10091 27319
rect 1409 26945 1443 26979
rect 9873 26945 9907 26979
rect 1593 26741 1627 26775
rect 10057 26741 10091 26775
rect 1409 26333 1443 26367
rect 9873 26333 9907 26367
rect 10977 26333 11011 26367
rect 1593 26197 1627 26231
rect 10057 26197 10091 26231
rect 10977 26197 11011 26231
rect 10057 25993 10091 26027
rect 1409 25857 1443 25891
rect 9137 25857 9171 25891
rect 9873 25857 9907 25891
rect 1593 25653 1627 25687
rect 9321 25653 9355 25687
rect 9965 25313 9999 25347
rect 10977 25245 11011 25279
rect 9873 25177 9907 25211
rect 9413 25109 9447 25143
rect 9781 25109 9815 25143
rect 1409 24769 1443 24803
rect 9137 24769 9171 24803
rect 9965 24769 9999 24803
rect 10149 24769 10183 24803
rect 1593 24633 1627 24667
rect 9321 24633 9355 24667
rect 9321 24361 9355 24395
rect 10149 24293 10183 24327
rect 1409 24157 1443 24191
rect 9137 24157 9171 24191
rect 9965 24157 9999 24191
rect 1593 24021 1627 24055
rect 8861 23817 8895 23851
rect 9321 23817 9355 23851
rect 9873 23817 9907 23851
rect 1409 23681 1443 23715
rect 8769 23681 8803 23715
rect 9781 23681 9815 23715
rect 10057 23613 10091 23647
rect 9413 23545 9447 23579
rect 1593 23477 1627 23511
rect 9873 23137 9907 23171
rect 10057 23137 10091 23171
rect 1409 23069 1443 23103
rect 9781 23001 9815 23035
rect 1593 22933 1627 22967
rect 9413 22933 9447 22967
rect 8677 22729 8711 22763
rect 9873 22661 9907 22695
rect 1409 22593 1443 22627
rect 8585 22593 8619 22627
rect 9781 22593 9815 22627
rect 8861 22525 8895 22559
rect 10057 22525 10091 22559
rect 9413 22457 9447 22491
rect 1593 22389 1627 22423
rect 8217 22389 8251 22423
rect 11161 31569 11195 31603
rect 11621 47957 11655 47991
rect 11713 50337 11747 50371
rect 11529 41837 11563 41871
rect 11621 47821 11655 47855
rect 11437 41225 11471 41259
rect 11529 41701 11563 41735
rect 11345 41021 11379 41055
rect 11345 33269 11379 33303
rect 11437 40069 11471 40103
rect 11437 32861 11471 32895
rect 11345 32793 11379 32827
rect 11345 30889 11379 30923
rect 11437 32725 11471 32759
rect 11253 24157 11287 24191
rect 11345 30753 11379 30787
rect 11161 22593 11195 22627
rect 11437 22661 11471 22695
rect 8401 22049 8435 22083
rect 9597 22049 9631 22083
rect 11345 22117 11379 22151
rect 9321 21981 9355 22015
rect 10977 21981 11011 22015
rect 8217 21913 8251 21947
rect 8585 21641 8619 21675
rect 8493 21573 8527 21607
rect 1409 21505 1443 21539
rect 9597 21505 9631 21539
rect 8769 21437 8803 21471
rect 9321 21437 9355 21471
rect 1593 21369 1627 21403
rect 8125 21301 8159 21335
rect 9597 20961 9631 20995
rect 1409 20893 1443 20927
rect 9321 20893 9355 20927
rect 1593 20757 1627 20791
rect 8125 20553 8159 20587
rect 8769 20553 8803 20587
rect 9229 20485 9263 20519
rect 10241 20485 10275 20519
rect 1409 20417 1443 20451
rect 8309 20417 8343 20451
rect 8953 20417 8987 20451
rect 1593 20213 1627 20247
rect 8217 20009 8251 20043
rect 9873 19873 9907 19907
rect 9965 19873 9999 19907
rect 1409 19805 1443 19839
rect 8401 19805 8435 19839
rect 1593 19669 1627 19703
rect 9413 19669 9447 19703
rect 9781 19669 9815 19703
rect 8125 19465 8159 19499
rect 8769 19465 8803 19499
rect 9137 19465 9171 19499
rect 9965 19397 9999 19431
rect 10057 19397 10091 19431
rect 1409 19329 1443 19363
rect 8309 19329 8343 19363
rect 8953 19329 8987 19363
rect 9321 19329 9355 19363
rect 9781 19329 9815 19363
rect 9505 19193 9539 19227
rect 1593 19125 1627 19159
rect 7573 18921 7607 18955
rect 8217 18921 8251 18955
rect 10241 18921 10275 18955
rect 10057 18785 10091 18819
rect 7757 18717 7791 18751
rect 8401 18717 8435 18751
rect 9321 18717 9355 18751
rect 10425 18717 10459 18751
rect 9873 18649 9907 18683
rect 9413 18581 9447 18615
rect 9781 18581 9815 18615
rect 7113 18377 7147 18411
rect 9229 18377 9263 18411
rect 10241 18377 10275 18411
rect 1409 18241 1443 18275
rect 7297 18241 7331 18275
rect 8401 18241 8435 18275
rect 1593 18105 1627 18139
rect 8217 18037 8251 18071
rect 8401 17833 8435 17867
rect 9873 17697 9907 17731
rect 10057 17697 10091 17731
rect 1409 17629 1443 17663
rect 6561 17629 6595 17663
rect 7757 17629 7791 17663
rect 8242 17561 8276 17595
rect 1593 17493 1627 17527
rect 6653 17493 6687 17527
rect 8033 17493 8067 17527
rect 8125 17493 8159 17527
rect 9413 17493 9447 17527
rect 9781 17493 9815 17527
rect 9137 17289 9171 17323
rect 9229 17289 9263 17323
rect 9413 17289 9447 17323
rect 9873 17289 9907 17323
rect 10333 17221 10367 17255
rect 1409 17153 1443 17187
rect 6469 17153 6503 17187
rect 7113 17153 7147 17187
rect 8013 17153 8047 17187
rect 9229 17153 9263 17187
rect 9781 17153 9815 17187
rect 10241 17153 10275 17187
rect 7757 17085 7791 17119
rect 10057 17085 10091 17119
rect 6653 17017 6687 17051
rect 7297 17017 7331 17051
rect 1593 16949 1627 16983
rect 6469 16745 6503 16779
rect 7757 16609 7791 16643
rect 8125 16609 8159 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 1409 16541 1443 16575
rect 6469 16541 6503 16575
rect 6653 16541 6687 16575
rect 7113 16541 7147 16575
rect 9505 16541 9539 16575
rect 8242 16473 8276 16507
rect 1593 16405 1627 16439
rect 7205 16405 7239 16439
rect 8033 16405 8067 16439
rect 8401 16405 8435 16439
rect 9137 16405 9171 16439
rect 5641 16201 5675 16235
rect 8953 16201 8987 16235
rect 7840 16133 7874 16167
rect 9781 16133 9815 16167
rect 5825 16065 5859 16099
rect 7113 16065 7147 16099
rect 7573 16065 7607 16099
rect 9873 15997 9907 16031
rect 9965 15997 9999 16031
rect 6929 15861 6963 15895
rect 9413 15861 9447 15895
rect 8125 15657 8159 15691
rect 9321 15521 9355 15555
rect 10057 15521 10091 15555
rect 1409 15453 1443 15487
rect 6745 15453 6779 15487
rect 7389 15453 7423 15487
rect 8033 15453 8067 15487
rect 9873 15453 9907 15487
rect 7849 15385 7883 15419
rect 1593 15317 1627 15351
rect 6561 15317 6595 15351
rect 7205 15317 7239 15351
rect 9413 15317 9447 15351
rect 9781 15317 9815 15351
rect 6837 15113 6871 15147
rect 8677 15113 8711 15147
rect 9873 15113 9907 15147
rect 8585 15045 8619 15079
rect 1409 14977 1443 15011
rect 7021 14977 7055 15011
rect 7573 14977 7607 15011
rect 9321 14977 9355 15011
rect 9781 14977 9815 15011
rect 8769 14909 8803 14943
rect 9965 14909 9999 14943
rect 7757 14841 7791 14875
rect 1593 14773 1627 14807
rect 8217 14773 8251 14807
rect 9413 14773 9447 14807
rect 5273 14501 5307 14535
rect 7297 14433 7331 14467
rect 9873 14433 9907 14467
rect 9965 14433 9999 14467
rect 1409 14365 1443 14399
rect 5457 14365 5491 14399
rect 6101 14365 6135 14399
rect 6653 14365 6687 14399
rect 7665 14365 7699 14399
rect 7782 14365 7816 14399
rect 6837 14297 6871 14331
rect 9781 14297 9815 14331
rect 1593 14229 1627 14263
rect 5917 14229 5951 14263
rect 7573 14229 7607 14263
rect 7941 14229 7975 14263
rect 9413 14229 9447 14263
rect 5641 14025 5675 14059
rect 6377 14025 6411 14059
rect 7481 14025 7515 14059
rect 8217 14025 8251 14059
rect 8585 14025 8619 14059
rect 9873 14025 9907 14059
rect 1409 13889 1443 13923
rect 5825 13889 5859 13923
rect 6561 13889 6595 13923
rect 7389 13889 7423 13923
rect 8677 13889 8711 13923
rect 9781 13889 9815 13923
rect 7573 13821 7607 13855
rect 8861 13821 8895 13855
rect 9965 13821 9999 13855
rect 1593 13685 1627 13719
rect 7021 13685 7055 13719
rect 9413 13685 9447 13719
rect 6009 13481 6043 13515
rect 7665 13481 7699 13515
rect 5365 13345 5399 13379
rect 5641 13345 5675 13379
rect 7113 13345 7147 13379
rect 8217 13345 8251 13379
rect 9965 13345 9999 13379
rect 1409 13277 1443 13311
rect 5733 13277 5767 13311
rect 6837 13277 6871 13311
rect 9321 13277 9355 13311
rect 9873 13277 9907 13311
rect 5850 13209 5884 13243
rect 6929 13209 6963 13243
rect 1593 13141 1627 13175
rect 6469 13141 6503 13175
rect 8033 13141 8067 13175
rect 8125 13141 8159 13175
rect 9413 13141 9447 13175
rect 9781 13141 9815 13175
rect 7205 12937 7239 12971
rect 7573 12937 7607 12971
rect 7665 12937 7699 12971
rect 9689 12937 9723 12971
rect 8401 12869 8435 12903
rect 5641 12801 5675 12835
rect 6561 12801 6595 12835
rect 7849 12733 7883 12767
rect 5825 12665 5859 12699
rect 6653 12597 6687 12631
rect 8401 12393 8435 12427
rect 5733 12325 5767 12359
rect 7021 12257 7055 12291
rect 9873 12257 9907 12291
rect 9965 12257 9999 12291
rect 1409 12189 1443 12223
rect 5917 12189 5951 12223
rect 6377 12189 6411 12223
rect 6561 12189 6595 12223
rect 7266 12121 7300 12155
rect 1593 12053 1627 12087
rect 6469 12053 6503 12087
rect 9413 12053 9447 12087
rect 9781 12053 9815 12087
rect 9689 11849 9723 11883
rect 1409 11713 1443 11747
rect 6561 11713 6595 11747
rect 6828 11713 6862 11747
rect 8401 11713 8435 11747
rect 1593 11509 1627 11543
rect 7941 11509 7975 11543
rect 6469 11305 6503 11339
rect 8217 11305 8251 11339
rect 9229 11305 9263 11339
rect 10241 11305 10275 11339
rect 7113 11237 7147 11271
rect 1409 11101 1443 11135
rect 6653 11101 6687 11135
rect 7297 11101 7331 11135
rect 8125 11101 8159 11135
rect 1593 10965 1627 10999
rect 7113 10761 7147 10795
rect 7849 10761 7883 10795
rect 9781 10761 9815 10795
rect 9873 10761 9907 10795
rect 1409 10625 1443 10659
rect 6929 10625 6963 10659
rect 8033 10625 8067 10659
rect 8861 10625 8895 10659
rect 10425 10625 10459 10659
rect 8953 10557 8987 10591
rect 9137 10557 9171 10591
rect 9965 10557 9999 10591
rect 8493 10489 8527 10523
rect 9413 10489 9447 10523
rect 1593 10421 1627 10455
rect 10241 10421 10275 10455
rect 7205 10217 7239 10251
rect 9413 10217 9447 10251
rect 8217 10149 8251 10183
rect 9965 10081 9999 10115
rect 1409 10013 1443 10047
rect 7113 10013 7147 10047
rect 8401 10013 8435 10047
rect 9781 10013 9815 10047
rect 9873 9945 9907 9979
rect 1593 9877 1627 9911
rect 8677 9605 8711 9639
rect 8861 9605 8895 9639
rect 7849 9537 7883 9571
rect 9781 9537 9815 9571
rect 8033 9401 8067 9435
rect 9873 9333 9907 9367
rect 9321 9129 9355 9163
rect 10057 9129 10091 9163
rect 1409 8925 1443 8959
rect 9137 8925 9171 8959
rect 9873 8925 9907 8959
rect 1593 8789 1627 8823
rect 11161 21913 11195 21947
rect 11345 21913 11379 21947
rect 11805 41905 11839 41939
rect 11897 41769 11931 41803
rect 11805 41633 11839 41667
rect 11713 41089 11747 41123
rect 11713 31909 11747 31943
rect 11621 22253 11655 22287
rect 11713 31773 11747 31807
rect 11529 22049 11563 22083
rect 11621 22117 11655 22151
rect 11437 21913 11471 21947
rect 11529 21845 11563 21879
rect 11161 20961 11195 20995
rect 11345 21777 11379 21811
rect 11161 20825 11195 20859
rect 11161 18717 11195 18751
rect 11345 17357 11379 17391
rect 11437 21777 11471 21811
rect 11253 17085 11287 17119
rect 11345 17221 11379 17255
rect 11161 16269 11195 16303
rect 11253 16541 11287 16575
rect 11161 16133 11195 16167
rect 11253 15453 11287 15487
rect 11161 13413 11195 13447
rect 9229 8585 9263 8619
rect 10425 8585 10459 8619
rect 9137 8517 9171 8551
rect 9781 8517 9815 8551
rect 10977 8517 11011 8551
rect 1409 8449 1443 8483
rect 10241 8449 10275 8483
rect 10057 8381 10091 8415
rect 1593 8313 1627 8347
rect 10057 8041 10091 8075
rect 1409 7837 1443 7871
rect 9781 7769 9815 7803
rect 1593 7701 1627 7735
rect 9137 7497 9171 7531
rect 9873 7497 9907 7531
rect 1409 7361 1443 7395
rect 8953 7361 8987 7395
rect 9781 7361 9815 7395
rect 9965 7293 9999 7327
rect 9413 7225 9447 7259
rect 1593 7157 1627 7191
rect 9873 6817 9907 6851
rect 9965 6817 9999 6851
rect 11069 7497 11103 7531
rect 10977 6749 11011 6783
rect 9781 6681 9815 6715
rect 9413 6613 9447 6647
rect 9229 6409 9263 6443
rect 10241 6409 10275 6443
rect 1409 6273 1443 6307
rect 8769 6273 8803 6307
rect 1593 6137 1627 6171
rect 8861 6069 8895 6103
rect 9413 5729 9447 5763
rect 9597 5729 9631 5763
rect 1409 5661 1443 5695
rect 8125 5661 8159 5695
rect 8401 5593 8435 5627
rect 9321 5593 9355 5627
rect 1593 5525 1627 5559
rect 8953 5525 8987 5559
rect 11529 21709 11563 21743
rect 11621 21709 11655 21743
rect 11621 18649 11655 18683
rect 11621 17357 11655 17391
rect 11897 40613 11931 40647
rect 11897 40477 11931 40511
rect 11897 33337 11931 33371
rect 11805 31637 11839 31671
rect 11897 32657 11931 32691
rect 11713 17221 11747 17255
rect 11805 31297 11839 31331
rect 11897 31297 11931 31331
rect 11621 17085 11655 17119
rect 11621 10149 11655 10183
rect 11713 9129 11747 9163
rect 11529 8993 11563 9027
rect 11897 29665 11931 29699
rect 11897 22729 11931 22763
rect 11897 21913 11931 21947
rect 11897 13277 11931 13311
rect 11805 8585 11839 8619
rect 11437 8381 11471 8415
rect 11345 8041 11379 8075
rect 8125 5321 8159 5355
rect 9873 5321 9907 5355
rect 11161 5321 11195 5355
rect 9321 5253 9355 5287
rect 1409 5185 1443 5219
rect 8309 5185 8343 5219
rect 8953 5185 8987 5219
rect 9781 5185 9815 5219
rect 9965 5117 9999 5151
rect 9413 5049 9447 5083
rect 1593 4981 1627 5015
rect 8769 4981 8803 5015
rect 9321 4777 9355 4811
rect 9873 4641 9907 4675
rect 9965 4641 9999 4675
rect 1409 4573 1443 4607
rect 9781 4573 9815 4607
rect 1593 4437 1627 4471
rect 9413 4437 9447 4471
rect 1409 4097 1443 4131
rect 8861 4097 8895 4131
rect 9321 4097 9355 4131
rect 9597 4097 9631 4131
rect 8677 3961 8711 3995
rect 1593 3893 1627 3927
rect 8217 3689 8251 3723
rect 9597 3553 9631 3587
rect 1409 3485 1443 3519
rect 8401 3485 8435 3519
rect 9321 3485 9355 3519
rect 1593 3349 1627 3383
rect 9873 3145 9907 3179
rect 1409 3009 1443 3043
rect 7665 3009 7699 3043
rect 8401 3009 8435 3043
rect 7849 2873 7883 2907
rect 1593 2805 1627 2839
rect 7573 2465 7607 2499
rect 9597 2465 9631 2499
rect 1409 2397 1443 2431
rect 2145 2397 2179 2431
rect 3065 2397 3099 2431
rect 7849 2397 7883 2431
rect 9321 2397 9355 2431
rect 1593 2261 1627 2295
rect 2329 2261 2363 2295
rect 2881 2261 2915 2295
<< metal1 >>
rect 1104 77818 10856 77840
rect 1104 77766 2582 77818
rect 2634 77766 2646 77818
rect 2698 77766 2710 77818
rect 2762 77766 2774 77818
rect 2826 77766 2838 77818
rect 2890 77766 5845 77818
rect 5897 77766 5909 77818
rect 5961 77766 5973 77818
rect 6025 77766 6037 77818
rect 6089 77766 6101 77818
rect 6153 77766 9109 77818
rect 9161 77766 9173 77818
rect 9225 77766 9237 77818
rect 9289 77766 9301 77818
rect 9353 77766 9365 77818
rect 9417 77766 10856 77818
rect 1104 77744 10856 77766
rect 7558 77704 7564 77716
rect 7519 77676 7564 77704
rect 7558 77664 7564 77676
rect 7616 77664 7622 77716
rect 8202 77664 8208 77716
rect 8260 77704 8266 77716
rect 8297 77707 8355 77713
rect 8297 77704 8309 77707
rect 8260 77676 8309 77704
rect 8260 77664 8266 77676
rect 8297 77673 8309 77676
rect 8343 77673 8355 77707
rect 8297 77667 8355 77673
rect 1394 77568 1400 77580
rect 1355 77540 1400 77568
rect 1394 77528 1400 77540
rect 1452 77528 1458 77580
rect 1673 77571 1731 77577
rect 1673 77537 1685 77571
rect 1719 77568 1731 77571
rect 11517 77571 11575 77577
rect 11517 77568 11529 77571
rect 1719 77540 11529 77568
rect 1719 77537 1731 77540
rect 1673 77531 1731 77537
rect 11517 77537 11529 77540
rect 11563 77537 11575 77571
rect 11517 77531 11575 77537
rect 2866 77500 2872 77512
rect 2827 77472 2872 77500
rect 2866 77460 2872 77472
rect 2924 77460 2930 77512
rect 6178 77460 6184 77512
rect 6236 77500 6242 77512
rect 7377 77503 7435 77509
rect 7377 77500 7389 77503
rect 6236 77472 7389 77500
rect 6236 77460 6242 77472
rect 7377 77469 7389 77472
rect 7423 77469 7435 77503
rect 7377 77463 7435 77469
rect 8113 77503 8171 77509
rect 8113 77469 8125 77503
rect 8159 77469 8171 77503
rect 8113 77463 8171 77469
rect 3142 77392 3148 77444
rect 3200 77432 3206 77444
rect 8128 77432 8156 77463
rect 8938 77460 8944 77512
rect 8996 77500 9002 77512
rect 9125 77503 9183 77509
rect 9125 77500 9137 77503
rect 8996 77472 9137 77500
rect 8996 77460 9002 77472
rect 9125 77469 9137 77472
rect 9171 77469 9183 77503
rect 9125 77463 9183 77469
rect 9861 77503 9919 77509
rect 9861 77469 9873 77503
rect 9907 77500 9919 77503
rect 11149 77503 11207 77509
rect 11149 77500 11161 77503
rect 9907 77472 11161 77500
rect 9907 77469 9919 77472
rect 9861 77463 9919 77469
rect 11149 77469 11161 77472
rect 11195 77469 11207 77503
rect 11149 77463 11207 77469
rect 3200 77404 8156 77432
rect 3200 77392 3206 77404
rect 2685 77367 2743 77373
rect 2685 77333 2697 77367
rect 2731 77364 2743 77367
rect 3050 77364 3056 77376
rect 2731 77336 3056 77364
rect 2731 77333 2743 77336
rect 2685 77327 2743 77333
rect 3050 77324 3056 77336
rect 3108 77324 3114 77376
rect 9306 77364 9312 77376
rect 9267 77336 9312 77364
rect 9306 77324 9312 77336
rect 9364 77324 9370 77376
rect 10045 77367 10103 77373
rect 10045 77333 10057 77367
rect 10091 77364 10103 77367
rect 10134 77364 10140 77376
rect 10091 77336 10140 77364
rect 10091 77333 10103 77336
rect 10045 77327 10103 77333
rect 10134 77324 10140 77336
rect 10192 77324 10198 77376
rect 1104 77274 10856 77296
rect 1104 77222 4213 77274
rect 4265 77222 4277 77274
rect 4329 77222 4341 77274
rect 4393 77222 4405 77274
rect 4457 77222 4469 77274
rect 4521 77222 7477 77274
rect 7529 77222 7541 77274
rect 7593 77222 7605 77274
rect 7657 77222 7669 77274
rect 7721 77222 7733 77274
rect 7785 77222 10856 77274
rect 1104 77200 10856 77222
rect 1397 77163 1455 77169
rect 1397 77129 1409 77163
rect 1443 77160 1455 77163
rect 3694 77160 3700 77172
rect 1443 77132 3700 77160
rect 1443 77129 1455 77132
rect 1397 77123 1455 77129
rect 3694 77120 3700 77132
rect 3752 77120 3758 77172
rect 8570 77160 8576 77172
rect 8531 77132 8576 77160
rect 8570 77120 8576 77132
rect 8628 77120 8634 77172
rect 9309 77163 9367 77169
rect 9309 77129 9321 77163
rect 9355 77160 9367 77163
rect 9582 77160 9588 77172
rect 9355 77132 9588 77160
rect 9355 77129 9367 77132
rect 9309 77123 9367 77129
rect 9582 77120 9588 77132
rect 9640 77120 9646 77172
rect 2958 77092 2964 77104
rect 2792 77064 2964 77092
rect 1578 77024 1584 77036
rect 1539 76996 1584 77024
rect 1578 76984 1584 76996
rect 1636 76984 1642 77036
rect 2225 77027 2283 77033
rect 2225 76993 2237 77027
rect 2271 77024 2283 77027
rect 2792 77024 2820 77064
rect 2958 77052 2964 77064
rect 3016 77052 3022 77104
rect 2271 76996 2820 77024
rect 2869 77027 2927 77033
rect 2271 76993 2283 76996
rect 2225 76987 2283 76993
rect 2869 76993 2881 77027
rect 2915 77024 2927 77027
rect 3234 77024 3240 77036
rect 2915 76996 3240 77024
rect 2915 76993 2927 76996
rect 2869 76987 2927 76993
rect 3234 76984 3240 76996
rect 3292 76984 3298 77036
rect 8386 77024 8392 77036
rect 8347 76996 8392 77024
rect 8386 76984 8392 76996
rect 8444 76984 8450 77036
rect 9125 77027 9183 77033
rect 9125 76993 9137 77027
rect 9171 76993 9183 77027
rect 9125 76987 9183 76993
rect 9861 77027 9919 77033
rect 9861 76993 9873 77027
rect 9907 77024 9919 77027
rect 11057 77027 11115 77033
rect 11057 77024 11069 77027
rect 9907 76996 11069 77024
rect 9907 76993 9919 76996
rect 9861 76987 9919 76993
rect 11057 76993 11069 76996
rect 11103 76993 11115 77027
rect 11057 76987 11115 76993
rect 3326 76916 3332 76968
rect 3384 76956 3390 76968
rect 9140 76956 9168 76987
rect 3384 76928 9168 76956
rect 3384 76916 3390 76928
rect 2041 76891 2099 76897
rect 2041 76857 2053 76891
rect 2087 76888 2099 76891
rect 2958 76888 2964 76900
rect 2087 76860 2964 76888
rect 2087 76857 2099 76860
rect 2041 76851 2099 76857
rect 2958 76848 2964 76860
rect 3016 76848 3022 76900
rect 2685 76823 2743 76829
rect 2685 76789 2697 76823
rect 2731 76820 2743 76823
rect 6454 76820 6460 76832
rect 2731 76792 6460 76820
rect 2731 76789 2743 76792
rect 2685 76783 2743 76789
rect 6454 76780 6460 76792
rect 6512 76780 6518 76832
rect 10042 76820 10048 76832
rect 10003 76792 10048 76820
rect 10042 76780 10048 76792
rect 10100 76780 10106 76832
rect 1104 76730 10856 76752
rect 1104 76678 2582 76730
rect 2634 76678 2646 76730
rect 2698 76678 2710 76730
rect 2762 76678 2774 76730
rect 2826 76678 2838 76730
rect 2890 76678 5845 76730
rect 5897 76678 5909 76730
rect 5961 76678 5973 76730
rect 6025 76678 6037 76730
rect 6089 76678 6101 76730
rect 6153 76678 9109 76730
rect 9161 76678 9173 76730
rect 9225 76678 9237 76730
rect 9289 76678 9301 76730
rect 9353 76678 9365 76730
rect 9417 76678 10856 76730
rect 1104 76656 10856 76678
rect 9309 76619 9367 76625
rect 9309 76585 9321 76619
rect 9355 76616 9367 76619
rect 9490 76616 9496 76628
rect 9355 76588 9496 76616
rect 9355 76585 9367 76588
rect 9309 76579 9367 76585
rect 9490 76576 9496 76588
rect 9548 76576 9554 76628
rect 1578 76412 1584 76424
rect 1539 76384 1584 76412
rect 1578 76372 1584 76384
rect 1636 76372 1642 76424
rect 8294 76372 8300 76424
rect 8352 76412 8358 76424
rect 9125 76415 9183 76421
rect 9125 76412 9137 76415
rect 8352 76384 9137 76412
rect 8352 76372 8358 76384
rect 9125 76381 9137 76384
rect 9171 76381 9183 76415
rect 9125 76375 9183 76381
rect 9861 76415 9919 76421
rect 9861 76381 9873 76415
rect 9907 76412 9919 76415
rect 11241 76415 11299 76421
rect 11241 76412 11253 76415
rect 9907 76384 11253 76412
rect 9907 76381 9919 76384
rect 9861 76375 9919 76381
rect 11241 76381 11253 76384
rect 11287 76381 11299 76415
rect 11241 76375 11299 76381
rect 1397 76279 1455 76285
rect 1397 76245 1409 76279
rect 1443 76276 1455 76279
rect 2130 76276 2136 76288
rect 1443 76248 2136 76276
rect 1443 76245 1455 76248
rect 1397 76239 1455 76245
rect 2130 76236 2136 76248
rect 2188 76236 2194 76288
rect 10042 76276 10048 76288
rect 10003 76248 10048 76276
rect 10042 76236 10048 76248
rect 10100 76236 10106 76288
rect 1104 76186 10856 76208
rect 1104 76134 4213 76186
rect 4265 76134 4277 76186
rect 4329 76134 4341 76186
rect 4393 76134 4405 76186
rect 4457 76134 4469 76186
rect 4521 76134 7477 76186
rect 7529 76134 7541 76186
rect 7593 76134 7605 76186
rect 7657 76134 7669 76186
rect 7721 76134 7733 76186
rect 7785 76134 10856 76186
rect 1104 76112 10856 76134
rect 9306 76072 9312 76084
rect 9267 76044 9312 76072
rect 9306 76032 9312 76044
rect 9364 76032 9370 76084
rect 1673 75939 1731 75945
rect 1673 75905 1685 75939
rect 1719 75936 1731 75939
rect 1762 75936 1768 75948
rect 1719 75908 1768 75936
rect 1719 75905 1731 75908
rect 1673 75899 1731 75905
rect 1762 75896 1768 75908
rect 1820 75896 1826 75948
rect 8478 75896 8484 75948
rect 8536 75936 8542 75948
rect 9125 75939 9183 75945
rect 9125 75936 9137 75939
rect 8536 75908 9137 75936
rect 8536 75896 8542 75908
rect 9125 75905 9137 75908
rect 9171 75905 9183 75939
rect 9858 75936 9864 75948
rect 9819 75908 9864 75936
rect 9125 75899 9183 75905
rect 9858 75896 9864 75908
rect 9916 75896 9922 75948
rect 1394 75868 1400 75880
rect 1355 75840 1400 75868
rect 1394 75828 1400 75840
rect 1452 75828 1458 75880
rect 10045 75735 10103 75741
rect 10045 75701 10057 75735
rect 10091 75732 10103 75735
rect 10965 75735 11023 75741
rect 10965 75732 10977 75735
rect 10091 75704 10977 75732
rect 10091 75701 10103 75704
rect 10045 75695 10103 75701
rect 10965 75701 10977 75704
rect 11011 75701 11023 75735
rect 10965 75695 11023 75701
rect 1104 75642 10856 75664
rect 1104 75590 2582 75642
rect 2634 75590 2646 75642
rect 2698 75590 2710 75642
rect 2762 75590 2774 75642
rect 2826 75590 2838 75642
rect 2890 75590 5845 75642
rect 5897 75590 5909 75642
rect 5961 75590 5973 75642
rect 6025 75590 6037 75642
rect 6089 75590 6101 75642
rect 6153 75590 9109 75642
rect 9161 75590 9173 75642
rect 9225 75590 9237 75642
rect 9289 75590 9301 75642
rect 9353 75590 9365 75642
rect 9417 75590 10856 75642
rect 1104 75568 10856 75590
rect 9861 75327 9919 75333
rect 9861 75293 9873 75327
rect 9907 75324 9919 75327
rect 11701 75327 11759 75333
rect 11701 75324 11713 75327
rect 9907 75296 11713 75324
rect 9907 75293 9919 75296
rect 9861 75287 9919 75293
rect 11701 75293 11713 75296
rect 11747 75293 11759 75327
rect 11701 75287 11759 75293
rect 1854 75256 1860 75268
rect 1815 75228 1860 75256
rect 1854 75216 1860 75228
rect 1912 75216 1918 75268
rect 1946 75188 1952 75200
rect 1907 75160 1952 75188
rect 1946 75148 1952 75160
rect 2004 75148 2010 75200
rect 10045 75191 10103 75197
rect 10045 75157 10057 75191
rect 10091 75188 10103 75191
rect 10134 75188 10140 75200
rect 10091 75160 10140 75188
rect 10091 75157 10103 75160
rect 10045 75151 10103 75157
rect 10134 75148 10140 75160
rect 10192 75148 10198 75200
rect 1104 75098 10856 75120
rect 1104 75046 4213 75098
rect 4265 75046 4277 75098
rect 4329 75046 4341 75098
rect 4393 75046 4405 75098
rect 4457 75046 4469 75098
rect 4521 75046 7477 75098
rect 7529 75046 7541 75098
rect 7593 75046 7605 75098
rect 7657 75046 7669 75098
rect 7721 75046 7733 75098
rect 7785 75046 10856 75098
rect 1104 75024 10856 75046
rect 2685 74987 2743 74993
rect 2685 74953 2697 74987
rect 2731 74953 2743 74987
rect 3050 74984 3056 74996
rect 3011 74956 3056 74984
rect 2685 74947 2743 74953
rect 2700 74916 2728 74947
rect 3050 74944 3056 74956
rect 3108 74944 3114 74996
rect 10873 74987 10931 74993
rect 10873 74953 10885 74987
rect 10919 74984 10931 74987
rect 11057 74987 11115 74993
rect 11057 74984 11069 74987
rect 10919 74956 11069 74984
rect 10919 74953 10931 74956
rect 10873 74947 10931 74953
rect 11057 74953 11069 74956
rect 11103 74953 11115 74987
rect 11057 74947 11115 74953
rect 3142 74916 3148 74928
rect 2700 74888 3148 74916
rect 3142 74876 3148 74888
rect 3200 74876 3206 74928
rect 10962 74916 10968 74928
rect 10923 74888 10968 74916
rect 10962 74876 10968 74888
rect 11020 74876 11026 74928
rect 1578 74848 1584 74860
rect 1539 74820 1584 74848
rect 1578 74808 1584 74820
rect 1636 74808 1642 74860
rect 2222 74848 2228 74860
rect 2183 74820 2228 74848
rect 2222 74808 2228 74820
rect 2280 74808 2286 74860
rect 9861 74851 9919 74857
rect 9861 74817 9873 74851
rect 9907 74848 9919 74851
rect 11149 74851 11207 74857
rect 11149 74848 11161 74851
rect 9907 74820 11161 74848
rect 9907 74817 9919 74820
rect 9861 74811 9919 74817
rect 11149 74817 11161 74820
rect 11195 74817 11207 74851
rect 11149 74811 11207 74817
rect 2498 74740 2504 74792
rect 2556 74780 2562 74792
rect 3142 74780 3148 74792
rect 2556 74752 2774 74780
rect 3103 74752 3148 74780
rect 2556 74740 2562 74752
rect 1397 74715 1455 74721
rect 1397 74681 1409 74715
rect 1443 74712 1455 74715
rect 2746 74712 2774 74752
rect 3142 74740 3148 74752
rect 3200 74740 3206 74792
rect 3237 74783 3295 74789
rect 3237 74749 3249 74783
rect 3283 74749 3295 74783
rect 3237 74743 3295 74749
rect 3252 74712 3280 74743
rect 1443 74684 2636 74712
rect 2746 74684 3280 74712
rect 1443 74681 1455 74684
rect 1397 74675 1455 74681
rect 2038 74644 2044 74656
rect 1999 74616 2044 74644
rect 2038 74604 2044 74616
rect 2096 74604 2102 74656
rect 2608 74644 2636 74684
rect 4614 74644 4620 74656
rect 2608 74616 4620 74644
rect 4614 74604 4620 74616
rect 4672 74604 4678 74656
rect 10042 74644 10048 74656
rect 10003 74616 10048 74644
rect 10042 74604 10048 74616
rect 10100 74604 10106 74656
rect 1104 74554 10856 74576
rect 1104 74502 2582 74554
rect 2634 74502 2646 74554
rect 2698 74502 2710 74554
rect 2762 74502 2774 74554
rect 2826 74502 2838 74554
rect 2890 74502 5845 74554
rect 5897 74502 5909 74554
rect 5961 74502 5973 74554
rect 6025 74502 6037 74554
rect 6089 74502 6101 74554
rect 6153 74502 9109 74554
rect 9161 74502 9173 74554
rect 9225 74502 9237 74554
rect 9289 74502 9301 74554
rect 9353 74502 9365 74554
rect 9417 74502 10856 74554
rect 1104 74480 10856 74502
rect 6089 74443 6147 74449
rect 6089 74409 6101 74443
rect 6135 74440 6147 74443
rect 6178 74440 6184 74452
rect 6135 74412 6184 74440
rect 6135 74409 6147 74412
rect 6089 74403 6147 74409
rect 6178 74400 6184 74412
rect 6236 74400 6242 74452
rect 8386 74400 8392 74452
rect 8444 74440 8450 74452
rect 9401 74443 9459 74449
rect 9401 74440 9413 74443
rect 8444 74412 9413 74440
rect 8444 74400 8450 74412
rect 9401 74409 9413 74412
rect 9447 74409 9459 74443
rect 9401 74403 9459 74409
rect 1949 74375 2007 74381
rect 1949 74341 1961 74375
rect 1995 74372 2007 74375
rect 8938 74372 8944 74384
rect 1995 74344 8944 74372
rect 1995 74341 2007 74344
rect 1949 74335 2007 74341
rect 8938 74332 8944 74344
rect 8996 74332 9002 74384
rect 2498 74304 2504 74316
rect 2459 74276 2504 74304
rect 2498 74264 2504 74276
rect 2556 74264 2562 74316
rect 6733 74307 6791 74313
rect 6733 74273 6745 74307
rect 6779 74304 6791 74307
rect 6822 74304 6828 74316
rect 6779 74276 6828 74304
rect 6779 74273 6791 74276
rect 6733 74267 6791 74273
rect 6822 74264 6828 74276
rect 6880 74264 6886 74316
rect 10045 74307 10103 74313
rect 10045 74273 10057 74307
rect 10091 74304 10103 74307
rect 10226 74304 10232 74316
rect 10091 74276 10232 74304
rect 10091 74273 10103 74276
rect 10045 74267 10103 74273
rect 10226 74264 10232 74276
rect 10284 74264 10290 74316
rect 2314 74196 2320 74248
rect 2372 74236 2378 74248
rect 2409 74239 2467 74245
rect 2409 74236 2421 74239
rect 2372 74208 2421 74236
rect 2372 74196 2378 74208
rect 2409 74205 2421 74208
rect 2455 74205 2467 74239
rect 2409 74199 2467 74205
rect 9769 74239 9827 74245
rect 9769 74205 9781 74239
rect 9815 74236 9827 74239
rect 11517 74239 11575 74245
rect 11517 74236 11529 74239
rect 9815 74208 11529 74236
rect 9815 74205 9827 74208
rect 9769 74199 9827 74205
rect 9968 74180 9996 74208
rect 11517 74205 11529 74208
rect 11563 74205 11575 74239
rect 11517 74199 11575 74205
rect 6454 74168 6460 74180
rect 6367 74140 6460 74168
rect 6454 74128 6460 74140
rect 6512 74168 6518 74180
rect 6638 74168 6644 74180
rect 6512 74140 6644 74168
rect 6512 74128 6518 74140
rect 6638 74128 6644 74140
rect 6696 74128 6702 74180
rect 9950 74128 9956 74180
rect 10008 74128 10014 74180
rect 2130 74060 2136 74112
rect 2188 74100 2194 74112
rect 2317 74103 2375 74109
rect 2317 74100 2329 74103
rect 2188 74072 2329 74100
rect 2188 74060 2194 74072
rect 2317 74069 2329 74072
rect 2363 74069 2375 74103
rect 2317 74063 2375 74069
rect 6362 74060 6368 74112
rect 6420 74100 6426 74112
rect 6549 74103 6607 74109
rect 6549 74100 6561 74103
rect 6420 74072 6561 74100
rect 6420 74060 6426 74072
rect 6549 74069 6561 74072
rect 6595 74069 6607 74103
rect 6549 74063 6607 74069
rect 9861 74103 9919 74109
rect 9861 74069 9873 74103
rect 9907 74100 9919 74103
rect 10134 74100 10140 74112
rect 9907 74072 10140 74100
rect 9907 74069 9919 74072
rect 9861 74063 9919 74069
rect 10134 74060 10140 74072
rect 10192 74060 10198 74112
rect 1104 74010 10856 74032
rect 1104 73958 4213 74010
rect 4265 73958 4277 74010
rect 4329 73958 4341 74010
rect 4393 73958 4405 74010
rect 4457 73958 4469 74010
rect 4521 73958 7477 74010
rect 7529 73958 7541 74010
rect 7593 73958 7605 74010
rect 7657 73958 7669 74010
rect 7721 73958 7733 74010
rect 7785 73958 10856 74010
rect 1104 73936 10856 73958
rect 1581 73899 1639 73905
rect 1581 73865 1593 73899
rect 1627 73896 1639 73899
rect 3326 73896 3332 73908
rect 1627 73868 2774 73896
rect 3287 73868 3332 73896
rect 1627 73865 1639 73868
rect 1581 73859 1639 73865
rect 2746 73828 2774 73868
rect 3326 73856 3332 73868
rect 3384 73856 3390 73908
rect 10965 73899 11023 73905
rect 10965 73896 10977 73899
rect 6886 73868 10977 73896
rect 6886 73828 6914 73868
rect 10965 73865 10977 73868
rect 11011 73865 11023 73899
rect 10965 73859 11023 73865
rect 2746 73800 6914 73828
rect 1946 73760 1952 73772
rect 1859 73732 1952 73760
rect 1946 73720 1952 73732
rect 2004 73760 2010 73772
rect 2406 73760 2412 73772
rect 2004 73732 2412 73760
rect 2004 73720 2010 73732
rect 2406 73720 2412 73732
rect 2464 73720 2470 73772
rect 3694 73760 3700 73772
rect 3655 73732 3700 73760
rect 3694 73720 3700 73732
rect 3752 73720 3758 73772
rect 3789 73763 3847 73769
rect 3789 73729 3801 73763
rect 3835 73760 3847 73763
rect 4062 73760 4068 73772
rect 3835 73732 4068 73760
rect 3835 73729 3847 73732
rect 3789 73723 3847 73729
rect 4062 73720 4068 73732
rect 4120 73720 4126 73772
rect 8662 73720 8668 73772
rect 8720 73760 8726 73772
rect 9125 73763 9183 73769
rect 9125 73760 9137 73763
rect 8720 73732 9137 73760
rect 8720 73720 8726 73732
rect 9125 73729 9137 73732
rect 9171 73729 9183 73763
rect 9125 73723 9183 73729
rect 9861 73763 9919 73769
rect 9861 73729 9873 73763
rect 9907 73760 9919 73763
rect 10965 73763 11023 73769
rect 10965 73760 10977 73763
rect 9907 73732 10977 73760
rect 9907 73729 9919 73732
rect 9861 73723 9919 73729
rect 10965 73729 10977 73732
rect 11011 73729 11023 73763
rect 10965 73723 11023 73729
rect 2041 73695 2099 73701
rect 2041 73692 2053 73695
rect 1964 73664 2053 73692
rect 1964 73636 1992 73664
rect 2041 73661 2053 73664
rect 2087 73661 2099 73695
rect 2041 73655 2099 73661
rect 2225 73695 2283 73701
rect 2225 73661 2237 73695
rect 2271 73692 2283 73695
rect 2498 73692 2504 73704
rect 2271 73664 2504 73692
rect 2271 73661 2283 73664
rect 2225 73655 2283 73661
rect 2498 73652 2504 73664
rect 2556 73692 2562 73704
rect 3973 73695 4031 73701
rect 3973 73692 3985 73695
rect 2556 73664 3985 73692
rect 2556 73652 2562 73664
rect 3973 73661 3985 73664
rect 4019 73692 4031 73695
rect 6822 73692 6828 73704
rect 4019 73664 6828 73692
rect 4019 73661 4031 73664
rect 3973 73655 4031 73661
rect 6822 73652 6828 73664
rect 6880 73652 6886 73704
rect 1946 73584 1952 73636
rect 2004 73584 2010 73636
rect 9309 73559 9367 73565
rect 9309 73525 9321 73559
rect 9355 73556 9367 73559
rect 9490 73556 9496 73568
rect 9355 73528 9496 73556
rect 9355 73525 9367 73528
rect 9309 73519 9367 73525
rect 9490 73516 9496 73528
rect 9548 73516 9554 73568
rect 10042 73556 10048 73568
rect 10003 73528 10048 73556
rect 10042 73516 10048 73528
rect 10100 73516 10106 73568
rect 1104 73466 10856 73488
rect 1104 73414 2582 73466
rect 2634 73414 2646 73466
rect 2698 73414 2710 73466
rect 2762 73414 2774 73466
rect 2826 73414 2838 73466
rect 2890 73414 5845 73466
rect 5897 73414 5909 73466
rect 5961 73414 5973 73466
rect 6025 73414 6037 73466
rect 6089 73414 6101 73466
rect 6153 73414 9109 73466
rect 9161 73414 9173 73466
rect 9225 73414 9237 73466
rect 9289 73414 9301 73466
rect 9353 73414 9365 73466
rect 9417 73414 10856 73466
rect 1104 73392 10856 73414
rect 2130 73312 2136 73364
rect 2188 73352 2194 73364
rect 2188 73324 2636 73352
rect 2188 73312 2194 73324
rect 2608 73296 2636 73324
rect 2590 73244 2596 73296
rect 2648 73244 2654 73296
rect 2133 73219 2191 73225
rect 2133 73185 2145 73219
rect 2179 73216 2191 73219
rect 2498 73216 2504 73228
rect 2179 73188 2504 73216
rect 2179 73185 2191 73188
rect 2133 73179 2191 73185
rect 2498 73176 2504 73188
rect 2556 73176 2562 73228
rect 6822 73176 6828 73228
rect 6880 73216 6886 73228
rect 7653 73219 7711 73225
rect 7653 73216 7665 73219
rect 6880 73188 7665 73216
rect 6880 73176 6886 73188
rect 7653 73185 7665 73188
rect 7699 73185 7711 73219
rect 7653 73179 7711 73185
rect 9953 73219 10011 73225
rect 9953 73185 9965 73219
rect 9999 73216 10011 73219
rect 10134 73216 10140 73228
rect 9999 73188 10140 73216
rect 9999 73185 10011 73188
rect 9953 73179 10011 73185
rect 10134 73176 10140 73188
rect 10192 73216 10198 73228
rect 11793 73219 11851 73225
rect 11793 73216 11805 73219
rect 10192 73188 11805 73216
rect 10192 73176 10198 73188
rect 11793 73185 11805 73188
rect 11839 73185 11851 73219
rect 11793 73179 11851 73185
rect 1670 73108 1676 73160
rect 1728 73148 1734 73160
rect 1949 73151 2007 73157
rect 1949 73148 1961 73151
rect 1728 73120 1961 73148
rect 1728 73108 1734 73120
rect 1949 73117 1961 73120
rect 1995 73117 2007 73151
rect 2866 73148 2872 73160
rect 2827 73120 2872 73148
rect 1949 73111 2007 73117
rect 2866 73108 2872 73120
rect 2924 73108 2930 73160
rect 9858 73148 9864 73160
rect 7116 73120 9864 73148
rect 6914 73080 6920 73092
rect 1504 73052 6920 73080
rect 1504 73021 1532 73052
rect 6914 73040 6920 73052
rect 6972 73040 6978 73092
rect 1489 73015 1547 73021
rect 1489 72981 1501 73015
rect 1535 72981 1547 73015
rect 1489 72975 1547 72981
rect 1762 72972 1768 73024
rect 1820 73012 1826 73024
rect 1857 73015 1915 73021
rect 1857 73012 1869 73015
rect 1820 72984 1869 73012
rect 1820 72972 1826 72984
rect 1857 72981 1869 72984
rect 1903 73012 1915 73015
rect 2130 73012 2136 73024
rect 1903 72984 2136 73012
rect 1903 72981 1915 72984
rect 1857 72975 1915 72981
rect 2130 72972 2136 72984
rect 2188 72972 2194 73024
rect 2685 73015 2743 73021
rect 2685 72981 2697 73015
rect 2731 73012 2743 73015
rect 7006 73012 7012 73024
rect 2731 72984 7012 73012
rect 2731 72981 2743 72984
rect 2685 72975 2743 72981
rect 7006 72972 7012 72984
rect 7064 72972 7070 73024
rect 7116 73021 7144 73120
rect 9858 73108 9864 73120
rect 9916 73108 9922 73160
rect 10045 73151 10103 73157
rect 10045 73117 10057 73151
rect 10091 73148 10103 73151
rect 10226 73148 10232 73160
rect 10091 73120 10232 73148
rect 10091 73117 10103 73120
rect 10045 73111 10103 73117
rect 10226 73108 10232 73120
rect 10284 73108 10290 73160
rect 7374 73040 7380 73092
rect 7432 73080 7438 73092
rect 7561 73083 7619 73089
rect 7561 73080 7573 73083
rect 7432 73052 7573 73080
rect 7432 73040 7438 73052
rect 7561 73049 7573 73052
rect 7607 73049 7619 73083
rect 9950 73080 9956 73092
rect 9911 73052 9956 73080
rect 7561 73043 7619 73049
rect 9950 73040 9956 73052
rect 10008 73040 10014 73092
rect 7101 73015 7159 73021
rect 7101 72981 7113 73015
rect 7147 72981 7159 73015
rect 7101 72975 7159 72981
rect 7282 72972 7288 73024
rect 7340 73012 7346 73024
rect 7469 73015 7527 73021
rect 7469 73012 7481 73015
rect 7340 72984 7481 73012
rect 7340 72972 7346 72984
rect 7469 72981 7481 72984
rect 7515 72981 7527 73015
rect 7469 72975 7527 72981
rect 8570 72972 8576 73024
rect 8628 73012 8634 73024
rect 9475 73015 9533 73021
rect 9475 73012 9487 73015
rect 8628 72984 9487 73012
rect 8628 72972 8634 72984
rect 9475 72981 9487 72984
rect 9521 72981 9533 73015
rect 9475 72975 9533 72981
rect 1104 72922 10856 72944
rect 1104 72870 4213 72922
rect 4265 72870 4277 72922
rect 4329 72870 4341 72922
rect 4393 72870 4405 72922
rect 4457 72870 4469 72922
rect 4521 72870 7477 72922
rect 7529 72870 7541 72922
rect 7593 72870 7605 72922
rect 7657 72870 7669 72922
rect 7721 72870 7733 72922
rect 7785 72870 10856 72922
rect 1104 72848 10856 72870
rect 1762 72808 1768 72820
rect 1675 72780 1768 72808
rect 1762 72768 1768 72780
rect 1820 72808 1826 72820
rect 2038 72808 2044 72820
rect 1820 72780 2044 72808
rect 1820 72768 1826 72780
rect 2038 72768 2044 72780
rect 2096 72768 2102 72820
rect 2593 72811 2651 72817
rect 2593 72777 2605 72811
rect 2639 72808 2651 72811
rect 8294 72808 8300 72820
rect 2639 72780 8300 72808
rect 2639 72777 2651 72780
rect 2593 72771 2651 72777
rect 8294 72768 8300 72780
rect 8352 72768 8358 72820
rect 2222 72700 2228 72752
rect 2280 72740 2286 72752
rect 2498 72740 2504 72752
rect 2280 72712 2504 72740
rect 2280 72700 2286 72712
rect 2498 72700 2504 72712
rect 2556 72740 2562 72752
rect 2556 72712 3096 72740
rect 2556 72700 2562 72712
rect 934 72632 940 72684
rect 992 72672 998 72684
rect 2958 72672 2964 72684
rect 992 72644 2774 72672
rect 2919 72644 2964 72672
rect 992 72632 998 72644
rect 1854 72604 1860 72616
rect 1815 72576 1860 72604
rect 1854 72564 1860 72576
rect 1912 72564 1918 72616
rect 2041 72607 2099 72613
rect 2041 72573 2053 72607
rect 2087 72604 2099 72607
rect 2222 72604 2228 72616
rect 2087 72576 2228 72604
rect 2087 72573 2099 72576
rect 2041 72567 2099 72573
rect 2222 72564 2228 72576
rect 2280 72564 2286 72616
rect 2746 72604 2774 72644
rect 2958 72632 2964 72644
rect 3016 72632 3022 72684
rect 3068 72672 3096 72712
rect 6914 72700 6920 72752
rect 6972 72740 6978 72752
rect 11057 72743 11115 72749
rect 11057 72740 11069 72743
rect 6972 72712 11069 72740
rect 6972 72700 6978 72712
rect 11057 72709 11069 72712
rect 11103 72709 11115 72743
rect 11057 72703 11115 72709
rect 3068 72644 3188 72672
rect 3160 72613 3188 72644
rect 9030 72632 9036 72684
rect 9088 72672 9094 72684
rect 9125 72675 9183 72681
rect 9125 72672 9137 72675
rect 9088 72644 9137 72672
rect 9088 72632 9094 72644
rect 9125 72641 9137 72644
rect 9171 72641 9183 72675
rect 9125 72635 9183 72641
rect 9861 72675 9919 72681
rect 9861 72641 9873 72675
rect 9907 72672 9919 72675
rect 11609 72675 11667 72681
rect 11609 72672 11621 72675
rect 9907 72644 11621 72672
rect 9907 72641 9919 72644
rect 9861 72635 9919 72641
rect 11609 72641 11621 72644
rect 11655 72641 11667 72675
rect 11609 72635 11667 72641
rect 3053 72607 3111 72613
rect 3053 72604 3065 72607
rect 2746 72576 3065 72604
rect 3053 72573 3065 72576
rect 3099 72573 3111 72607
rect 3053 72567 3111 72573
rect 3145 72607 3203 72613
rect 3145 72573 3157 72607
rect 3191 72573 3203 72607
rect 3145 72567 3203 72573
rect 1397 72539 1455 72545
rect 1397 72505 1409 72539
rect 1443 72536 1455 72539
rect 9306 72536 9312 72548
rect 1443 72508 2544 72536
rect 1443 72505 1455 72508
rect 1397 72499 1455 72505
rect 2516 72468 2544 72508
rect 2746 72508 3004 72536
rect 9267 72508 9312 72536
rect 2746 72468 2774 72508
rect 2516 72440 2774 72468
rect 2976 72468 3004 72508
rect 9306 72496 9312 72508
rect 9364 72496 9370 72548
rect 8478 72468 8484 72480
rect 2976 72440 8484 72468
rect 8478 72428 8484 72440
rect 8536 72428 8542 72480
rect 10045 72471 10103 72477
rect 10045 72437 10057 72471
rect 10091 72468 10103 72471
rect 10134 72468 10140 72480
rect 10091 72440 10140 72468
rect 10091 72437 10103 72440
rect 10045 72431 10103 72437
rect 10134 72428 10140 72440
rect 10192 72428 10198 72480
rect 1104 72378 10856 72400
rect 1104 72326 2582 72378
rect 2634 72326 2646 72378
rect 2698 72326 2710 72378
rect 2762 72326 2774 72378
rect 2826 72326 2838 72378
rect 2890 72326 5845 72378
rect 5897 72326 5909 72378
rect 5961 72326 5973 72378
rect 6025 72326 6037 72378
rect 6089 72326 6101 72378
rect 6153 72326 9109 72378
rect 9161 72326 9173 72378
rect 9225 72326 9237 72378
rect 9289 72326 9301 72378
rect 9353 72326 9365 72378
rect 9417 72326 10856 72378
rect 1104 72304 10856 72326
rect 1397 72199 1455 72205
rect 1397 72165 1409 72199
rect 1443 72196 1455 72199
rect 3142 72196 3148 72208
rect 1443 72168 3148 72196
rect 1443 72165 1455 72168
rect 1397 72159 1455 72165
rect 3142 72156 3148 72168
rect 3200 72156 3206 72208
rect 6178 72196 6184 72208
rect 6139 72168 6184 72196
rect 6178 72156 6184 72168
rect 6236 72156 6242 72208
rect 3694 72088 3700 72140
rect 3752 72128 3758 72140
rect 3752 72100 4200 72128
rect 3752 72088 3758 72100
rect 1578 72060 1584 72072
rect 1539 72032 1584 72060
rect 1578 72020 1584 72032
rect 1636 72020 1642 72072
rect 2222 72060 2228 72072
rect 2183 72032 2228 72060
rect 2222 72020 2228 72032
rect 2280 72020 2286 72072
rect 4062 72060 4068 72072
rect 4023 72032 4068 72060
rect 4062 72020 4068 72032
rect 4120 72020 4126 72072
rect 4172 72069 4200 72100
rect 4157 72063 4215 72069
rect 4157 72029 4169 72063
rect 4203 72029 4215 72063
rect 4157 72023 4215 72029
rect 4341 72063 4399 72069
rect 4341 72029 4353 72063
rect 4387 72060 4399 72063
rect 6733 72063 6791 72069
rect 6733 72060 6745 72063
rect 4387 72032 6745 72060
rect 4387 72029 4399 72032
rect 4341 72023 4399 72029
rect 6733 72029 6745 72032
rect 6779 72029 6791 72063
rect 6733 72023 6791 72029
rect 4798 71992 4804 72004
rect 4759 71964 4804 71992
rect 4798 71952 4804 71964
rect 4856 71952 4862 72004
rect 5718 71952 5724 72004
rect 5776 71992 5782 72004
rect 6362 71992 6368 72004
rect 5776 71964 6368 71992
rect 5776 71952 5782 71964
rect 6362 71952 6368 71964
rect 6420 71992 6426 72004
rect 6457 71995 6515 72001
rect 6457 71992 6469 71995
rect 6420 71964 6469 71992
rect 6420 71952 6426 71964
rect 6457 71961 6469 71964
rect 6503 71961 6515 71995
rect 6638 71992 6644 72004
rect 6599 71964 6644 71992
rect 6457 71955 6515 71961
rect 6638 71952 6644 71964
rect 6696 71952 6702 72004
rect 6748 71992 6776 72023
rect 6822 72020 6828 72072
rect 6880 72060 6886 72072
rect 9125 72063 9183 72069
rect 9125 72060 9137 72063
rect 6880 72032 9137 72060
rect 6880 72020 6886 72032
rect 9125 72029 9137 72032
rect 9171 72029 9183 72063
rect 9125 72023 9183 72029
rect 9769 72063 9827 72069
rect 9769 72029 9781 72063
rect 9815 72060 9827 72063
rect 9861 72063 9919 72069
rect 9861 72060 9873 72063
rect 9815 72032 9873 72060
rect 9815 72029 9827 72032
rect 9769 72023 9827 72029
rect 9861 72029 9873 72032
rect 9907 72060 9919 72063
rect 11333 72063 11391 72069
rect 11333 72060 11345 72063
rect 9907 72032 11345 72060
rect 9907 72029 9919 72032
rect 9861 72023 9919 72029
rect 11333 72029 11345 72032
rect 11379 72029 11391 72063
rect 11333 72023 11391 72029
rect 6914 71992 6920 72004
rect 6748 71964 6920 71992
rect 6914 71952 6920 71964
rect 6972 71952 6978 72004
rect 2038 71924 2044 71936
rect 1999 71896 2044 71924
rect 2038 71884 2044 71896
rect 2096 71884 2102 71936
rect 9306 71924 9312 71936
rect 9267 71896 9312 71924
rect 9306 71884 9312 71896
rect 9364 71884 9370 71936
rect 10042 71924 10048 71936
rect 10003 71896 10048 71924
rect 10042 71884 10048 71896
rect 10100 71884 10106 71936
rect 1104 71834 10856 71856
rect 1104 71782 4213 71834
rect 4265 71782 4277 71834
rect 4329 71782 4341 71834
rect 4393 71782 4405 71834
rect 4457 71782 4469 71834
rect 4521 71782 7477 71834
rect 7529 71782 7541 71834
rect 7593 71782 7605 71834
rect 7657 71782 7669 71834
rect 7721 71782 7733 71834
rect 7785 71782 10856 71834
rect 1104 71760 10856 71782
rect 1486 71544 1492 71596
rect 1544 71584 1550 71596
rect 1581 71587 1639 71593
rect 1581 71584 1593 71587
rect 1544 71556 1593 71584
rect 1544 71544 1550 71556
rect 1581 71553 1593 71556
rect 1627 71553 1639 71587
rect 1581 71547 1639 71553
rect 9861 71587 9919 71593
rect 9861 71553 9873 71587
rect 9907 71584 9919 71587
rect 11057 71587 11115 71593
rect 11057 71584 11069 71587
rect 9907 71556 11069 71584
rect 9907 71553 9919 71556
rect 9861 71547 9919 71553
rect 11057 71553 11069 71556
rect 11103 71553 11115 71587
rect 11057 71547 11115 71553
rect 2130 71476 2136 71528
rect 2188 71516 2194 71528
rect 2314 71516 2320 71528
rect 2188 71488 2320 71516
rect 2188 71476 2194 71488
rect 2314 71476 2320 71488
rect 2372 71476 2378 71528
rect 1397 71383 1455 71389
rect 1397 71349 1409 71383
rect 1443 71380 1455 71383
rect 9766 71380 9772 71392
rect 1443 71352 9772 71380
rect 1443 71349 1455 71352
rect 1397 71343 1455 71349
rect 9766 71340 9772 71352
rect 9824 71340 9830 71392
rect 10045 71383 10103 71389
rect 10045 71349 10057 71383
rect 10091 71380 10103 71383
rect 10134 71380 10140 71392
rect 10091 71352 10140 71380
rect 10091 71349 10103 71352
rect 10045 71343 10103 71349
rect 10134 71340 10140 71352
rect 10192 71340 10198 71392
rect 1104 71290 10856 71312
rect 1104 71238 2582 71290
rect 2634 71238 2646 71290
rect 2698 71238 2710 71290
rect 2762 71238 2774 71290
rect 2826 71238 2838 71290
rect 2890 71238 5845 71290
rect 5897 71238 5909 71290
rect 5961 71238 5973 71290
rect 6025 71238 6037 71290
rect 6089 71238 6101 71290
rect 6153 71238 9109 71290
rect 9161 71238 9173 71290
rect 9225 71238 9237 71290
rect 9289 71238 9301 71290
rect 9353 71238 9365 71290
rect 9417 71238 10856 71290
rect 1104 71216 10856 71238
rect 7098 71108 7104 71120
rect 1688 71080 7104 71108
rect 1688 71049 1716 71080
rect 7098 71068 7104 71080
rect 7156 71068 7162 71120
rect 11149 71111 11207 71117
rect 11149 71077 11161 71111
rect 11195 71108 11207 71111
rect 11425 71111 11483 71117
rect 11425 71108 11437 71111
rect 11195 71080 11437 71108
rect 11195 71077 11207 71080
rect 11149 71071 11207 71077
rect 11425 71077 11437 71080
rect 11471 71077 11483 71111
rect 11425 71071 11483 71077
rect 1673 71043 1731 71049
rect 1673 71009 1685 71043
rect 1719 71009 1731 71043
rect 1673 71003 1731 71009
rect 2130 71000 2136 71052
rect 2188 71040 2194 71052
rect 2590 71040 2596 71052
rect 2188 71012 2596 71040
rect 2188 71000 2194 71012
rect 2590 71000 2596 71012
rect 2648 71040 2654 71052
rect 4433 71043 4491 71049
rect 4433 71040 4445 71043
rect 2648 71012 4445 71040
rect 2648 71000 2654 71012
rect 4433 71009 4445 71012
rect 4479 71040 4491 71043
rect 6914 71040 6920 71052
rect 4479 71012 6920 71040
rect 4479 71009 4491 71012
rect 4433 71003 4491 71009
rect 6914 71000 6920 71012
rect 6972 71040 6978 71052
rect 7926 71040 7932 71052
rect 6972 71012 7932 71040
rect 6972 71000 6978 71012
rect 7926 71000 7932 71012
rect 7984 71000 7990 71052
rect 1394 70972 1400 70984
rect 1355 70944 1400 70972
rect 1394 70932 1400 70944
rect 1452 70932 1458 70984
rect 4157 70975 4215 70981
rect 4157 70941 4169 70975
rect 4203 70972 4215 70975
rect 4614 70972 4620 70984
rect 4203 70944 4620 70972
rect 4203 70941 4215 70944
rect 4157 70935 4215 70941
rect 4614 70932 4620 70944
rect 4672 70932 4678 70984
rect 9861 70975 9919 70981
rect 9861 70941 9873 70975
rect 9907 70972 9919 70975
rect 11149 70975 11207 70981
rect 11149 70972 11161 70975
rect 9907 70944 11161 70972
rect 9907 70941 9919 70944
rect 9861 70935 9919 70941
rect 11149 70941 11161 70944
rect 11195 70941 11207 70975
rect 11149 70935 11207 70941
rect 11241 70907 11299 70913
rect 11241 70904 11253 70907
rect 3804 70876 11253 70904
rect 3804 70845 3832 70876
rect 11241 70873 11253 70876
rect 11287 70873 11299 70907
rect 11241 70867 11299 70873
rect 3789 70839 3847 70845
rect 3789 70805 3801 70839
rect 3835 70805 3847 70839
rect 3789 70799 3847 70805
rect 3878 70796 3884 70848
rect 3936 70836 3942 70848
rect 4249 70839 4307 70845
rect 4249 70836 4261 70839
rect 3936 70808 4261 70836
rect 3936 70796 3942 70808
rect 4249 70805 4261 70808
rect 4295 70805 4307 70839
rect 10042 70836 10048 70848
rect 10003 70808 10048 70836
rect 4249 70799 4307 70805
rect 10042 70796 10048 70808
rect 10100 70796 10106 70848
rect 1104 70746 10856 70768
rect 1104 70694 4213 70746
rect 4265 70694 4277 70746
rect 4329 70694 4341 70746
rect 4393 70694 4405 70746
rect 4457 70694 4469 70746
rect 4521 70694 7477 70746
rect 7529 70694 7541 70746
rect 7593 70694 7605 70746
rect 7657 70694 7669 70746
rect 7721 70694 7733 70746
rect 7785 70694 10856 70746
rect 1104 70672 10856 70694
rect 2498 70592 2504 70644
rect 2556 70592 2562 70644
rect 2516 70564 2544 70592
rect 2424 70536 2544 70564
rect 2222 70496 2228 70508
rect 2183 70468 2228 70496
rect 2222 70456 2228 70468
rect 2280 70456 2286 70508
rect 2317 70499 2375 70505
rect 2317 70465 2329 70499
rect 2363 70496 2375 70499
rect 2424 70496 2452 70536
rect 2363 70468 2452 70496
rect 2501 70499 2559 70505
rect 2363 70465 2375 70468
rect 2317 70459 2375 70465
rect 2501 70465 2513 70499
rect 2547 70496 2559 70499
rect 2590 70496 2596 70508
rect 2547 70468 2596 70496
rect 2547 70465 2559 70468
rect 2501 70459 2559 70465
rect 2590 70456 2596 70468
rect 2648 70456 2654 70508
rect 5074 70496 5080 70508
rect 2884 70468 5080 70496
rect 2240 70428 2268 70456
rect 2884 70428 2912 70468
rect 5074 70456 5080 70468
rect 5132 70456 5138 70508
rect 7282 70456 7288 70508
rect 7340 70496 7346 70508
rect 7469 70499 7527 70505
rect 7469 70496 7481 70499
rect 7340 70468 7481 70496
rect 7340 70456 7346 70468
rect 7469 70465 7481 70468
rect 7515 70465 7527 70499
rect 7469 70459 7527 70465
rect 7653 70499 7711 70505
rect 7653 70465 7665 70499
rect 7699 70496 7711 70499
rect 7926 70496 7932 70508
rect 7699 70468 7932 70496
rect 7699 70465 7711 70468
rect 7653 70459 7711 70465
rect 7926 70456 7932 70468
rect 7984 70456 7990 70508
rect 2240 70400 2912 70428
rect 2961 70431 3019 70437
rect 2961 70397 2973 70431
rect 3007 70428 3019 70431
rect 4890 70428 4896 70440
rect 3007 70400 4896 70428
rect 3007 70397 3019 70400
rect 2961 70391 3019 70397
rect 4890 70388 4896 70400
rect 4948 70388 4954 70440
rect 7374 70428 7380 70440
rect 7335 70400 7380 70428
rect 7374 70388 7380 70400
rect 7432 70388 7438 70440
rect 7834 70388 7840 70440
rect 7892 70428 7898 70440
rect 8113 70431 8171 70437
rect 8113 70428 8125 70431
rect 7892 70400 8125 70428
rect 7892 70388 7898 70400
rect 8113 70397 8125 70400
rect 8159 70397 8171 70431
rect 8113 70391 8171 70397
rect 9309 70431 9367 70437
rect 9309 70397 9321 70431
rect 9355 70428 9367 70431
rect 9858 70428 9864 70440
rect 9355 70400 9864 70428
rect 9355 70397 9367 70400
rect 9309 70391 9367 70397
rect 9858 70388 9864 70400
rect 9916 70428 9922 70440
rect 10229 70431 10287 70437
rect 10229 70428 10241 70431
rect 9916 70400 10241 70428
rect 9916 70388 9922 70400
rect 10229 70397 10241 70400
rect 10275 70397 10287 70431
rect 10229 70391 10287 70397
rect 1104 70202 10856 70224
rect 1104 70150 2582 70202
rect 2634 70150 2646 70202
rect 2698 70150 2710 70202
rect 2762 70150 2774 70202
rect 2826 70150 2838 70202
rect 2890 70150 5845 70202
rect 5897 70150 5909 70202
rect 5961 70150 5973 70202
rect 6025 70150 6037 70202
rect 6089 70150 6101 70202
rect 6153 70150 9109 70202
rect 9161 70150 9173 70202
rect 9225 70150 9237 70202
rect 9289 70150 9301 70202
rect 9353 70150 9365 70202
rect 9417 70150 10856 70202
rect 1104 70128 10856 70150
rect 9030 70048 9036 70100
rect 9088 70088 9094 70100
rect 9401 70091 9459 70097
rect 9401 70088 9413 70091
rect 9088 70060 9413 70088
rect 9088 70048 9094 70060
rect 9401 70057 9413 70060
rect 9447 70057 9459 70091
rect 9401 70051 9459 70057
rect 2869 70023 2927 70029
rect 2869 69989 2881 70023
rect 2915 70020 2927 70023
rect 7190 70020 7196 70032
rect 2915 69992 7196 70020
rect 2915 69989 2927 69992
rect 2869 69983 2927 69989
rect 7190 69980 7196 69992
rect 7248 69980 7254 70032
rect 1854 69952 1860 69964
rect 1688 69924 1860 69952
rect 1118 69844 1124 69896
rect 1176 69884 1182 69896
rect 1688 69893 1716 69924
rect 1854 69912 1860 69924
rect 1912 69912 1918 69964
rect 10045 69955 10103 69961
rect 10045 69921 10057 69955
rect 10091 69952 10103 69955
rect 10226 69952 10232 69964
rect 10091 69924 10232 69952
rect 10091 69921 10103 69924
rect 10045 69915 10103 69921
rect 10226 69912 10232 69924
rect 10284 69912 10290 69964
rect 1673 69887 1731 69893
rect 1673 69884 1685 69887
rect 1176 69856 1685 69884
rect 1176 69844 1182 69856
rect 1673 69853 1685 69856
rect 1719 69853 1731 69887
rect 1673 69847 1731 69853
rect 1762 69844 1768 69896
rect 1820 69884 1826 69896
rect 1949 69887 2007 69893
rect 1820 69856 1865 69884
rect 1820 69844 1826 69856
rect 1949 69853 1961 69887
rect 1995 69884 2007 69887
rect 2130 69884 2136 69896
rect 1995 69856 2136 69884
rect 1995 69853 2007 69856
rect 1949 69847 2007 69853
rect 2130 69844 2136 69856
rect 2188 69844 2194 69896
rect 2866 69844 2872 69896
rect 2924 69884 2930 69896
rect 3053 69887 3111 69893
rect 3053 69884 3065 69887
rect 2924 69856 3065 69884
rect 2924 69844 2930 69856
rect 3053 69853 3065 69856
rect 3099 69853 3111 69887
rect 3970 69884 3976 69896
rect 3931 69856 3976 69884
rect 3053 69847 3111 69853
rect 3970 69844 3976 69856
rect 4028 69844 4034 69896
rect 2409 69819 2467 69825
rect 2409 69785 2421 69819
rect 2455 69816 2467 69819
rect 3510 69816 3516 69828
rect 2455 69788 3516 69816
rect 2455 69785 2467 69788
rect 2409 69779 2467 69785
rect 3510 69776 3516 69788
rect 3568 69776 3574 69828
rect 9769 69819 9827 69825
rect 9769 69816 9781 69819
rect 3804 69788 9781 69816
rect 3804 69757 3832 69788
rect 9769 69785 9781 69788
rect 9815 69816 9827 69819
rect 9950 69816 9956 69828
rect 9815 69788 9956 69816
rect 9815 69785 9827 69788
rect 9769 69779 9827 69785
rect 9950 69776 9956 69788
rect 10008 69776 10014 69828
rect 3789 69751 3847 69757
rect 3789 69717 3801 69751
rect 3835 69717 3847 69751
rect 3789 69711 3847 69717
rect 8846 69708 8852 69760
rect 8904 69748 8910 69760
rect 9217 69751 9275 69757
rect 9217 69748 9229 69751
rect 8904 69720 9229 69748
rect 8904 69708 8910 69720
rect 9217 69717 9229 69720
rect 9263 69717 9275 69751
rect 9858 69748 9864 69760
rect 9819 69720 9864 69748
rect 9217 69711 9275 69717
rect 9858 69708 9864 69720
rect 9916 69708 9922 69760
rect 1104 69658 10856 69680
rect 1104 69606 4213 69658
rect 4265 69606 4277 69658
rect 4329 69606 4341 69658
rect 4393 69606 4405 69658
rect 4457 69606 4469 69658
rect 4521 69606 7477 69658
rect 7529 69606 7541 69658
rect 7593 69606 7605 69658
rect 7657 69606 7669 69658
rect 7721 69606 7733 69658
rect 7785 69606 10856 69658
rect 1104 69584 10856 69606
rect 1489 69547 1547 69553
rect 1489 69513 1501 69547
rect 1535 69513 1547 69547
rect 1489 69507 1547 69513
rect 1857 69547 1915 69553
rect 1857 69513 1869 69547
rect 1903 69544 1915 69547
rect 2038 69544 2044 69556
rect 1903 69516 2044 69544
rect 1903 69513 1915 69516
rect 1857 69507 1915 69513
rect 1504 69476 1532 69507
rect 2038 69504 2044 69516
rect 2096 69504 2102 69556
rect 9217 69547 9275 69553
rect 2746 69516 3556 69544
rect 2746 69476 2774 69516
rect 3326 69476 3332 69488
rect 1504 69448 2774 69476
rect 2884 69448 3332 69476
rect 1210 69368 1216 69420
rect 1268 69408 1274 69420
rect 2884 69408 2912 69448
rect 3326 69436 3332 69448
rect 3384 69436 3390 69488
rect 3528 69476 3556 69516
rect 9217 69513 9229 69547
rect 9263 69544 9275 69547
rect 9582 69544 9588 69556
rect 9263 69516 9588 69544
rect 9263 69513 9275 69516
rect 9217 69507 9275 69513
rect 9582 69504 9588 69516
rect 9640 69504 9646 69556
rect 10410 69544 10416 69556
rect 10371 69516 10416 69544
rect 10410 69504 10416 69516
rect 10468 69504 10474 69556
rect 11057 69547 11115 69553
rect 11057 69513 11069 69547
rect 11103 69544 11115 69547
rect 11241 69547 11299 69553
rect 11241 69544 11253 69547
rect 11103 69516 11253 69544
rect 11103 69513 11115 69516
rect 11057 69507 11115 69513
rect 11241 69513 11253 69516
rect 11287 69513 11299 69547
rect 11241 69507 11299 69513
rect 11701 69479 11759 69485
rect 11701 69476 11713 69479
rect 3528 69448 11713 69476
rect 11701 69445 11713 69448
rect 11747 69445 11759 69479
rect 11701 69439 11759 69445
rect 3050 69408 3056 69420
rect 1268 69380 2912 69408
rect 3011 69380 3056 69408
rect 1268 69368 1274 69380
rect 1949 69343 2007 69349
rect 1949 69309 1961 69343
rect 1995 69309 2007 69343
rect 2130 69340 2136 69352
rect 2091 69312 2136 69340
rect 1949 69303 2007 69309
rect 1964 69204 1992 69303
rect 2130 69300 2136 69312
rect 2188 69300 2194 69352
rect 2884 69340 2912 69380
rect 3050 69368 3056 69380
rect 3108 69368 3114 69420
rect 3237 69411 3295 69417
rect 3237 69377 3249 69411
rect 3283 69377 3295 69411
rect 8386 69408 8392 69420
rect 8347 69380 8392 69408
rect 3237 69371 3295 69377
rect 2961 69343 3019 69349
rect 2961 69340 2973 69343
rect 2884 69312 2973 69340
rect 2961 69309 2973 69312
rect 3007 69309 3019 69343
rect 2961 69303 3019 69309
rect 2148 69272 2176 69300
rect 2498 69272 2504 69284
rect 2148 69244 2504 69272
rect 2498 69232 2504 69244
rect 2556 69272 2562 69284
rect 3252 69272 3280 69371
rect 8386 69368 8392 69380
rect 8444 69368 8450 69420
rect 9030 69408 9036 69420
rect 8991 69380 9036 69408
rect 9030 69368 9036 69380
rect 9088 69368 9094 69420
rect 9766 69408 9772 69420
rect 9727 69380 9772 69408
rect 9766 69368 9772 69380
rect 9824 69368 9830 69420
rect 10229 69411 10287 69417
rect 10229 69377 10241 69411
rect 10275 69408 10287 69411
rect 11057 69411 11115 69417
rect 11057 69408 11069 69411
rect 10275 69380 11069 69408
rect 10275 69377 10287 69380
rect 10229 69371 10287 69377
rect 11057 69377 11069 69380
rect 11103 69377 11115 69411
rect 11057 69371 11115 69377
rect 3697 69343 3755 69349
rect 3697 69309 3709 69343
rect 3743 69340 3755 69343
rect 3786 69340 3792 69352
rect 3743 69312 3792 69340
rect 3743 69309 3755 69312
rect 3697 69303 3755 69309
rect 3786 69300 3792 69312
rect 3844 69300 3850 69352
rect 8846 69300 8852 69352
rect 8904 69340 8910 69352
rect 9861 69343 9919 69349
rect 9861 69340 9873 69343
rect 8904 69312 9873 69340
rect 8904 69300 8910 69312
rect 9861 69309 9873 69312
rect 9907 69309 9919 69343
rect 9861 69303 9919 69309
rect 10045 69343 10103 69349
rect 10045 69309 10057 69343
rect 10091 69340 10103 69343
rect 10134 69340 10140 69352
rect 10091 69312 10140 69340
rect 10091 69309 10103 69312
rect 10045 69303 10103 69309
rect 10134 69300 10140 69312
rect 10192 69300 10198 69352
rect 2556 69244 3280 69272
rect 8573 69275 8631 69281
rect 2556 69232 2562 69244
rect 8573 69241 8585 69275
rect 8619 69272 8631 69275
rect 9490 69272 9496 69284
rect 8619 69244 9496 69272
rect 8619 69241 8631 69244
rect 8573 69235 8631 69241
rect 9490 69232 9496 69244
rect 9548 69232 9554 69284
rect 3418 69204 3424 69216
rect 1964 69176 3424 69204
rect 3418 69164 3424 69176
rect 3476 69164 3482 69216
rect 9401 69207 9459 69213
rect 9401 69173 9413 69207
rect 9447 69204 9459 69207
rect 10965 69207 11023 69213
rect 10965 69204 10977 69207
rect 9447 69176 10977 69204
rect 9447 69173 9459 69176
rect 9401 69167 9459 69173
rect 10965 69173 10977 69176
rect 11011 69173 11023 69207
rect 10965 69167 11023 69173
rect 1104 69114 10856 69136
rect 1104 69062 2582 69114
rect 2634 69062 2646 69114
rect 2698 69062 2710 69114
rect 2762 69062 2774 69114
rect 2826 69062 2838 69114
rect 2890 69062 5845 69114
rect 5897 69062 5909 69114
rect 5961 69062 5973 69114
rect 6025 69062 6037 69114
rect 6089 69062 6101 69114
rect 6153 69062 9109 69114
rect 9161 69062 9173 69114
rect 9225 69062 9237 69114
rect 9289 69062 9301 69114
rect 9353 69062 9365 69114
rect 9417 69062 10856 69114
rect 1104 69040 10856 69062
rect 6822 69000 6828 69012
rect 6783 68972 6828 69000
rect 6822 68960 6828 68972
rect 6880 68960 6886 69012
rect 934 68824 940 68876
rect 992 68864 998 68876
rect 2501 68867 2559 68873
rect 2501 68864 2513 68867
rect 992 68836 2513 68864
rect 992 68824 998 68836
rect 2501 68833 2513 68836
rect 2547 68833 2559 68867
rect 2958 68864 2964 68876
rect 2501 68827 2559 68833
rect 2608 68836 2964 68864
rect 1578 68796 1584 68808
rect 1539 68768 1584 68796
rect 1578 68756 1584 68768
rect 1636 68756 1642 68808
rect 2608 68805 2636 68836
rect 2958 68824 2964 68836
rect 3016 68824 3022 68876
rect 7469 68867 7527 68873
rect 7469 68833 7481 68867
rect 7515 68864 7527 68867
rect 7926 68864 7932 68876
rect 7515 68836 7932 68864
rect 7515 68833 7527 68836
rect 7469 68827 7527 68833
rect 7926 68824 7932 68836
rect 7984 68824 7990 68876
rect 2593 68799 2651 68805
rect 2593 68765 2605 68799
rect 2639 68765 2651 68799
rect 2593 68759 2651 68765
rect 2777 68799 2835 68805
rect 2777 68765 2789 68799
rect 2823 68765 2835 68799
rect 7190 68796 7196 68808
rect 7151 68768 7196 68796
rect 2777 68759 2835 68765
rect 2498 68688 2504 68740
rect 2556 68728 2562 68740
rect 2792 68728 2820 68759
rect 7190 68756 7196 68768
rect 7248 68756 7254 68808
rect 8113 68799 8171 68805
rect 8113 68796 8125 68799
rect 7944 68768 8125 68796
rect 7944 68740 7972 68768
rect 8113 68765 8125 68768
rect 8159 68765 8171 68799
rect 8113 68759 8171 68765
rect 3234 68728 3240 68740
rect 2556 68700 2820 68728
rect 3195 68700 3240 68728
rect 2556 68688 2562 68700
rect 3234 68688 3240 68700
rect 3292 68688 3298 68740
rect 7006 68688 7012 68740
rect 7064 68728 7070 68740
rect 7285 68731 7343 68737
rect 7285 68728 7297 68731
rect 7064 68700 7297 68728
rect 7064 68688 7070 68700
rect 7285 68697 7297 68700
rect 7331 68697 7343 68731
rect 7285 68691 7343 68697
rect 7926 68688 7932 68740
rect 7984 68688 7990 68740
rect 1397 68663 1455 68669
rect 1397 68629 1409 68663
rect 1443 68660 1455 68663
rect 2314 68660 2320 68672
rect 1443 68632 2320 68660
rect 1443 68629 1455 68632
rect 1397 68623 1455 68629
rect 2314 68620 2320 68632
rect 2372 68620 2378 68672
rect 8202 68620 8208 68672
rect 8260 68660 8266 68672
rect 8297 68663 8355 68669
rect 8297 68660 8309 68663
rect 8260 68632 8309 68660
rect 8260 68620 8266 68632
rect 8297 68629 8309 68632
rect 8343 68629 8355 68663
rect 8297 68623 8355 68629
rect 8570 68620 8576 68672
rect 8628 68660 8634 68672
rect 9217 68663 9275 68669
rect 9217 68660 9229 68663
rect 8628 68632 9229 68660
rect 8628 68620 8634 68632
rect 9217 68629 9229 68632
rect 9263 68660 9275 68663
rect 9490 68660 9496 68672
rect 9263 68632 9496 68660
rect 9263 68629 9275 68632
rect 9217 68623 9275 68629
rect 9490 68620 9496 68632
rect 9548 68660 9554 68672
rect 9858 68660 9864 68672
rect 9548 68632 9864 68660
rect 9548 68620 9554 68632
rect 9858 68620 9864 68632
rect 9916 68660 9922 68672
rect 10229 68663 10287 68669
rect 10229 68660 10241 68663
rect 9916 68632 10241 68660
rect 9916 68620 9922 68632
rect 10229 68629 10241 68632
rect 10275 68629 10287 68663
rect 10229 68623 10287 68629
rect 1104 68570 10856 68592
rect 1104 68518 4213 68570
rect 4265 68518 4277 68570
rect 4329 68518 4341 68570
rect 4393 68518 4405 68570
rect 4457 68518 4469 68570
rect 4521 68518 7477 68570
rect 7529 68518 7541 68570
rect 7593 68518 7605 68570
rect 7657 68518 7669 68570
rect 7721 68518 7733 68570
rect 7785 68518 10856 68570
rect 1104 68496 10856 68518
rect 3878 68456 3884 68468
rect 3528 68428 3884 68456
rect 1486 68280 1492 68332
rect 1544 68320 1550 68332
rect 3528 68329 3556 68428
rect 3878 68416 3884 68428
rect 3936 68416 3942 68468
rect 9950 68456 9956 68468
rect 9911 68428 9956 68456
rect 9950 68416 9956 68428
rect 10008 68416 10014 68468
rect 4614 68388 4620 68400
rect 3620 68360 4620 68388
rect 3620 68329 3648 68360
rect 4614 68348 4620 68360
rect 4672 68348 4678 68400
rect 9490 68348 9496 68400
rect 9548 68388 9554 68400
rect 9769 68391 9827 68397
rect 9769 68388 9781 68391
rect 9548 68360 9781 68388
rect 9548 68348 9554 68360
rect 9769 68357 9781 68360
rect 9815 68357 9827 68391
rect 9769 68351 9827 68357
rect 10045 68391 10103 68397
rect 10045 68357 10057 68391
rect 10091 68388 10103 68391
rect 10134 68388 10140 68400
rect 10091 68360 10140 68388
rect 10091 68357 10103 68360
rect 10045 68351 10103 68357
rect 10134 68348 10140 68360
rect 10192 68348 10198 68400
rect 1581 68323 1639 68329
rect 1581 68320 1593 68323
rect 1544 68292 1593 68320
rect 1544 68280 1550 68292
rect 1581 68289 1593 68292
rect 1627 68289 1639 68323
rect 3513 68323 3571 68329
rect 3513 68320 3525 68323
rect 1581 68283 1639 68289
rect 2746 68292 3525 68320
rect 1302 68212 1308 68264
rect 1360 68252 1366 68264
rect 2746 68252 2774 68292
rect 3513 68289 3525 68292
rect 3559 68289 3571 68323
rect 3513 68283 3571 68289
rect 3605 68323 3663 68329
rect 3605 68289 3617 68323
rect 3651 68289 3663 68323
rect 3605 68283 3663 68289
rect 3789 68323 3847 68329
rect 3789 68289 3801 68323
rect 3835 68289 3847 68323
rect 3789 68283 3847 68289
rect 1360 68224 2774 68252
rect 1360 68212 1366 68224
rect 1578 68144 1584 68196
rect 1636 68184 1642 68196
rect 1946 68184 1952 68196
rect 1636 68156 1952 68184
rect 1636 68144 1642 68156
rect 1946 68144 1952 68156
rect 2004 68144 2010 68196
rect 2498 68144 2504 68196
rect 2556 68184 2562 68196
rect 3804 68184 3832 68283
rect 8202 68280 8208 68332
rect 8260 68320 8266 68332
rect 8573 68323 8631 68329
rect 8573 68320 8585 68323
rect 8260 68292 8585 68320
rect 8260 68280 8266 68292
rect 8573 68289 8585 68292
rect 8619 68289 8631 68323
rect 8573 68283 8631 68289
rect 4249 68255 4307 68261
rect 4249 68221 4261 68255
rect 4295 68252 4307 68255
rect 4614 68252 4620 68264
rect 4295 68224 4620 68252
rect 4295 68221 4307 68224
rect 4249 68215 4307 68221
rect 4614 68212 4620 68224
rect 4672 68212 4678 68264
rect 11609 68255 11667 68261
rect 11609 68221 11621 68255
rect 11655 68252 11667 68255
rect 11885 68255 11943 68261
rect 11885 68252 11897 68255
rect 11655 68224 11897 68252
rect 11655 68221 11667 68224
rect 11609 68215 11667 68221
rect 11885 68221 11897 68224
rect 11931 68221 11943 68255
rect 11885 68215 11943 68221
rect 2556 68156 3832 68184
rect 2556 68144 2562 68156
rect 1397 68119 1455 68125
rect 1397 68085 1409 68119
rect 1443 68116 1455 68119
rect 1762 68116 1768 68128
rect 1443 68088 1768 68116
rect 1443 68085 1455 68088
rect 1397 68079 1455 68085
rect 1762 68076 1768 68088
rect 1820 68076 1826 68128
rect 8754 68116 8760 68128
rect 8715 68088 8760 68116
rect 8754 68076 8760 68088
rect 8812 68076 8818 68128
rect 8846 68076 8852 68128
rect 8904 68116 8910 68128
rect 9125 68119 9183 68125
rect 9125 68116 9137 68119
rect 8904 68088 9137 68116
rect 8904 68076 8910 68088
rect 9125 68085 9137 68088
rect 9171 68085 9183 68119
rect 9125 68079 9183 68085
rect 9493 68119 9551 68125
rect 9493 68085 9505 68119
rect 9539 68116 9551 68119
rect 11609 68119 11667 68125
rect 11609 68116 11621 68119
rect 9539 68088 11621 68116
rect 9539 68085 9551 68088
rect 9493 68079 9551 68085
rect 11609 68085 11621 68088
rect 11655 68085 11667 68119
rect 11609 68079 11667 68085
rect 1104 68026 10856 68048
rect 1104 67974 2582 68026
rect 2634 67974 2646 68026
rect 2698 67974 2710 68026
rect 2762 67974 2774 68026
rect 2826 67974 2838 68026
rect 2890 67974 5845 68026
rect 5897 67974 5909 68026
rect 5961 67974 5973 68026
rect 6025 67974 6037 68026
rect 6089 67974 6101 68026
rect 6153 67974 9109 68026
rect 9161 67974 9173 68026
rect 9225 67974 9237 68026
rect 9289 67974 9301 68026
rect 9353 67974 9365 68026
rect 9417 67974 10856 68026
rect 1104 67952 10856 67974
rect 9398 67844 9404 67856
rect 9359 67816 9404 67844
rect 9398 67804 9404 67816
rect 9456 67804 9462 67856
rect 9953 67779 10011 67785
rect 9953 67745 9965 67779
rect 9999 67776 10011 67779
rect 10134 67776 10140 67788
rect 9999 67748 10140 67776
rect 9999 67745 10011 67748
rect 9953 67739 10011 67745
rect 10134 67736 10140 67748
rect 10192 67736 10198 67788
rect 1394 67708 1400 67720
rect 1355 67680 1400 67708
rect 1394 67668 1400 67680
rect 1452 67668 1458 67720
rect 1673 67711 1731 67717
rect 1673 67677 1685 67711
rect 1719 67708 1731 67711
rect 1946 67708 1952 67720
rect 1719 67680 1952 67708
rect 1719 67677 1731 67680
rect 1673 67671 1731 67677
rect 1946 67668 1952 67680
rect 2004 67668 2010 67720
rect 6914 67668 6920 67720
rect 6972 67708 6978 67720
rect 8113 67711 8171 67717
rect 8113 67708 8125 67711
rect 6972 67680 8125 67708
rect 6972 67668 6978 67680
rect 8113 67677 8125 67680
rect 8159 67677 8171 67711
rect 8113 67671 8171 67677
rect 8846 67600 8852 67652
rect 8904 67640 8910 67652
rect 9677 67643 9735 67649
rect 9677 67640 9689 67643
rect 8904 67612 9689 67640
rect 8904 67600 8910 67612
rect 9677 67609 9689 67612
rect 9723 67609 9735 67643
rect 9677 67603 9735 67609
rect 9766 67600 9772 67652
rect 9824 67640 9830 67652
rect 9861 67643 9919 67649
rect 9861 67640 9873 67643
rect 9824 67612 9873 67640
rect 9824 67600 9830 67612
rect 9861 67609 9873 67612
rect 9907 67609 9919 67643
rect 9861 67603 9919 67609
rect 8294 67572 8300 67584
rect 8255 67544 8300 67572
rect 8294 67532 8300 67544
rect 8352 67532 8358 67584
rect 1104 67482 10856 67504
rect 1104 67430 4213 67482
rect 4265 67430 4277 67482
rect 4329 67430 4341 67482
rect 4393 67430 4405 67482
rect 4457 67430 4469 67482
rect 4521 67430 7477 67482
rect 7529 67430 7541 67482
rect 7593 67430 7605 67482
rect 7657 67430 7669 67482
rect 7721 67430 7733 67482
rect 7785 67430 10856 67482
rect 1104 67408 10856 67430
rect 1762 67368 1768 67380
rect 1723 67340 1768 67368
rect 1762 67328 1768 67340
rect 1820 67328 1826 67380
rect 8386 67328 8392 67380
rect 8444 67368 8450 67380
rect 8665 67371 8723 67377
rect 8665 67368 8677 67371
rect 8444 67340 8677 67368
rect 8444 67328 8450 67340
rect 8665 67337 8677 67340
rect 8711 67337 8723 67371
rect 8665 67331 8723 67337
rect 9585 67371 9643 67377
rect 9585 67337 9597 67371
rect 9631 67368 9643 67371
rect 10134 67368 10140 67380
rect 9631 67340 10140 67368
rect 9631 67337 9643 67340
rect 9585 67331 9643 67337
rect 10134 67328 10140 67340
rect 10192 67328 10198 67380
rect 11241 67303 11299 67309
rect 11241 67300 11253 67303
rect 6932 67272 11253 67300
rect 2777 67235 2835 67241
rect 2777 67201 2789 67235
rect 2823 67232 2835 67235
rect 2958 67232 2964 67244
rect 2823 67204 2964 67232
rect 2823 67201 2835 67204
rect 2777 67195 2835 67201
rect 2958 67192 2964 67204
rect 3016 67192 3022 67244
rect 1854 67164 1860 67176
rect 1815 67136 1860 67164
rect 1854 67124 1860 67136
rect 1912 67124 1918 67176
rect 2041 67167 2099 67173
rect 2041 67133 2053 67167
rect 2087 67164 2099 67167
rect 2498 67164 2504 67176
rect 2087 67136 2504 67164
rect 2087 67133 2099 67136
rect 2041 67127 2099 67133
rect 2498 67124 2504 67136
rect 2556 67124 2562 67176
rect 1397 67099 1455 67105
rect 1397 67065 1409 67099
rect 1443 67096 1455 67099
rect 6932 67096 6960 67272
rect 11241 67269 11253 67272
rect 11287 67269 11299 67303
rect 11241 67263 11299 67269
rect 8294 67232 8300 67244
rect 8255 67204 8300 67232
rect 8294 67192 8300 67204
rect 8352 67192 8358 67244
rect 8938 67192 8944 67244
rect 8996 67232 9002 67244
rect 9033 67235 9091 67241
rect 9033 67232 9045 67235
rect 8996 67204 9045 67232
rect 8996 67192 9002 67204
rect 9033 67201 9045 67204
rect 9079 67201 9091 67235
rect 9033 67195 9091 67201
rect 9861 67235 9919 67241
rect 9861 67201 9873 67235
rect 9907 67201 9919 67235
rect 9861 67195 9919 67201
rect 9122 67164 9128 67176
rect 9083 67136 9128 67164
rect 9122 67124 9128 67136
rect 9180 67124 9186 67176
rect 9309 67167 9367 67173
rect 9309 67133 9321 67167
rect 9355 67164 9367 67167
rect 9585 67167 9643 67173
rect 9585 67164 9597 67167
rect 9355 67136 9597 67164
rect 9355 67133 9367 67136
rect 9309 67127 9367 67133
rect 9585 67133 9597 67136
rect 9631 67164 9643 67167
rect 9674 67164 9680 67176
rect 9631 67136 9680 67164
rect 9631 67133 9643 67136
rect 9585 67127 9643 67133
rect 9674 67124 9680 67136
rect 9732 67124 9738 67176
rect 1443 67068 6960 67096
rect 8481 67099 8539 67105
rect 1443 67065 1455 67068
rect 1397 67059 1455 67065
rect 8481 67065 8493 67099
rect 8527 67096 8539 67099
rect 9490 67096 9496 67108
rect 8527 67068 9496 67096
rect 8527 67065 8539 67068
rect 8481 67059 8539 67065
rect 9490 67056 9496 67068
rect 9548 67056 9554 67108
rect 9769 67099 9827 67105
rect 9769 67065 9781 67099
rect 9815 67096 9827 67099
rect 9876 67096 9904 67195
rect 11425 67099 11483 67105
rect 11425 67096 11437 67099
rect 9815 67068 11437 67096
rect 9815 67065 9827 67068
rect 9769 67059 9827 67065
rect 11425 67065 11437 67068
rect 11471 67065 11483 67099
rect 11425 67059 11483 67065
rect 2593 67031 2651 67037
rect 2593 66997 2605 67031
rect 2639 67028 2651 67031
rect 7374 67028 7380 67040
rect 2639 67000 7380 67028
rect 2639 66997 2651 67000
rect 2593 66991 2651 66997
rect 7374 66988 7380 67000
rect 7432 66988 7438 67040
rect 10042 67028 10048 67040
rect 10003 67000 10048 67028
rect 10042 66988 10048 67000
rect 10100 66988 10106 67040
rect 1104 66938 10856 66960
rect 1104 66886 2582 66938
rect 2634 66886 2646 66938
rect 2698 66886 2710 66938
rect 2762 66886 2774 66938
rect 2826 66886 2838 66938
rect 2890 66886 5845 66938
rect 5897 66886 5909 66938
rect 5961 66886 5973 66938
rect 6025 66886 6037 66938
rect 6089 66886 6101 66938
rect 6153 66886 9109 66938
rect 9161 66886 9173 66938
rect 9225 66886 9237 66938
rect 9289 66886 9301 66938
rect 9353 66886 9365 66938
rect 9417 66886 10856 66938
rect 1104 66864 10856 66886
rect 2041 66691 2099 66697
rect 2041 66657 2053 66691
rect 2087 66688 2099 66691
rect 3418 66688 3424 66700
rect 2087 66660 3424 66688
rect 2087 66657 2099 66660
rect 2041 66651 2099 66657
rect 3418 66648 3424 66660
rect 3476 66648 3482 66700
rect 3602 66648 3608 66700
rect 3660 66688 3666 66700
rect 3660 66660 9720 66688
rect 3660 66648 3666 66660
rect 2130 66580 2136 66632
rect 2188 66620 2194 66632
rect 2317 66623 2375 66629
rect 2188 66592 2233 66620
rect 2188 66580 2194 66592
rect 2317 66589 2329 66623
rect 2363 66620 2375 66623
rect 2498 66620 2504 66632
rect 2363 66592 2504 66620
rect 2363 66589 2375 66592
rect 2317 66583 2375 66589
rect 2498 66580 2504 66592
rect 2556 66620 2562 66632
rect 3620 66620 3648 66648
rect 2556 66592 3648 66620
rect 2556 66580 2562 66592
rect 7006 66580 7012 66632
rect 7064 66620 7070 66632
rect 7101 66623 7159 66629
rect 7101 66620 7113 66623
rect 7064 66592 7113 66620
rect 7064 66580 7070 66592
rect 7101 66589 7113 66592
rect 7147 66589 7159 66623
rect 7101 66583 7159 66589
rect 7190 66580 7196 66632
rect 7248 66620 7254 66632
rect 7392 66629 7420 66660
rect 9692 66632 9720 66660
rect 7377 66623 7435 66629
rect 7248 66592 7293 66620
rect 7248 66580 7254 66592
rect 7377 66589 7389 66623
rect 7423 66589 7435 66623
rect 7377 66583 7435 66589
rect 9030 66580 9036 66632
rect 9088 66620 9094 66632
rect 9398 66620 9404 66632
rect 9088 66592 9404 66620
rect 9088 66580 9094 66592
rect 9398 66580 9404 66592
rect 9456 66580 9462 66632
rect 9493 66623 9551 66629
rect 9493 66589 9505 66623
rect 9539 66589 9551 66623
rect 9674 66620 9680 66632
rect 9635 66592 9680 66620
rect 9493 66583 9551 66589
rect 2777 66555 2835 66561
rect 2777 66521 2789 66555
rect 2823 66552 2835 66555
rect 6270 66552 6276 66564
rect 2823 66524 6276 66552
rect 2823 66521 2835 66524
rect 2777 66515 2835 66521
rect 6270 66512 6276 66524
rect 6328 66512 6334 66564
rect 7837 66555 7895 66561
rect 7837 66521 7849 66555
rect 7883 66552 7895 66555
rect 8018 66552 8024 66564
rect 7883 66524 8024 66552
rect 7883 66521 7895 66524
rect 7837 66515 7895 66521
rect 8018 66512 8024 66524
rect 8076 66512 8082 66564
rect 8938 66512 8944 66564
rect 8996 66552 9002 66564
rect 9508 66552 9536 66583
rect 9674 66580 9680 66592
rect 9732 66580 9738 66632
rect 10134 66552 10140 66564
rect 8996 66524 9536 66552
rect 10095 66524 10140 66552
rect 8996 66512 9002 66524
rect 10134 66512 10140 66524
rect 10192 66512 10198 66564
rect 1104 66394 10856 66416
rect 1104 66342 4213 66394
rect 4265 66342 4277 66394
rect 4329 66342 4341 66394
rect 4393 66342 4405 66394
rect 4457 66342 4469 66394
rect 4521 66342 7477 66394
rect 7529 66342 7541 66394
rect 7593 66342 7605 66394
rect 7657 66342 7669 66394
rect 7721 66342 7733 66394
rect 7785 66342 10856 66394
rect 1104 66320 10856 66342
rect 2409 66215 2467 66221
rect 2409 66181 2421 66215
rect 2455 66212 2467 66215
rect 3050 66212 3056 66224
rect 2455 66184 3056 66212
rect 2455 66181 2467 66184
rect 2409 66175 2467 66181
rect 3050 66172 3056 66184
rect 3108 66172 3114 66224
rect 3142 66172 3148 66224
rect 3200 66212 3206 66224
rect 3237 66215 3295 66221
rect 3237 66212 3249 66215
rect 3200 66184 3249 66212
rect 3200 66172 3206 66184
rect 3237 66181 3249 66184
rect 3283 66181 3295 66215
rect 3237 66175 3295 66181
rect 1762 66144 1768 66156
rect 1723 66116 1768 66144
rect 1762 66104 1768 66116
rect 1820 66104 1826 66156
rect 1949 66147 2007 66153
rect 1949 66113 1961 66147
rect 1995 66144 2007 66147
rect 2498 66144 2504 66156
rect 1995 66116 2504 66144
rect 1995 66113 2007 66116
rect 1949 66107 2007 66113
rect 2498 66104 2504 66116
rect 2556 66104 2562 66156
rect 5626 66104 5632 66156
rect 5684 66144 5690 66156
rect 9125 66147 9183 66153
rect 9125 66144 9137 66147
rect 5684 66116 9137 66144
rect 5684 66104 5690 66116
rect 9125 66113 9137 66116
rect 9171 66113 9183 66147
rect 9125 66107 9183 66113
rect 9861 66147 9919 66153
rect 9861 66113 9873 66147
rect 9907 66144 9919 66147
rect 11698 66144 11704 66156
rect 9907 66116 11704 66144
rect 9907 66113 9919 66116
rect 9861 66107 9919 66113
rect 11698 66104 11704 66116
rect 11756 66104 11762 66156
rect 1673 66079 1731 66085
rect 1673 66045 1685 66079
rect 1719 66076 1731 66079
rect 1854 66076 1860 66088
rect 1719 66048 1860 66076
rect 1719 66045 1731 66048
rect 1673 66039 1731 66045
rect 1854 66036 1860 66048
rect 1912 66076 1918 66088
rect 1912 66048 2774 66076
rect 1912 66036 1918 66048
rect 2746 66008 2774 66048
rect 2958 66036 2964 66088
rect 3016 66076 3022 66088
rect 3329 66079 3387 66085
rect 3329 66076 3341 66079
rect 3016 66048 3341 66076
rect 3016 66036 3022 66048
rect 3329 66045 3341 66048
rect 3375 66045 3387 66079
rect 3329 66039 3387 66045
rect 3513 66079 3571 66085
rect 3513 66045 3525 66079
rect 3559 66076 3571 66079
rect 3602 66076 3608 66088
rect 3559 66048 3608 66076
rect 3559 66045 3571 66048
rect 3513 66039 3571 66045
rect 3602 66036 3608 66048
rect 3660 66036 3666 66088
rect 5166 66008 5172 66020
rect 2746 65980 5172 66008
rect 5166 65968 5172 65980
rect 5224 65968 5230 66020
rect 11517 66011 11575 66017
rect 11517 66008 11529 66011
rect 7116 65980 11529 66008
rect 2869 65943 2927 65949
rect 2869 65909 2881 65943
rect 2915 65940 2927 65943
rect 7116 65940 7144 65980
rect 11517 65977 11529 65980
rect 11563 65977 11575 66011
rect 11517 65971 11575 65977
rect 2915 65912 7144 65940
rect 9309 65943 9367 65949
rect 2915 65909 2927 65912
rect 2869 65903 2927 65909
rect 9309 65909 9321 65943
rect 9355 65940 9367 65943
rect 9490 65940 9496 65952
rect 9355 65912 9496 65940
rect 9355 65909 9367 65912
rect 9309 65903 9367 65909
rect 9490 65900 9496 65912
rect 9548 65900 9554 65952
rect 10042 65940 10048 65952
rect 10003 65912 10048 65940
rect 10042 65900 10048 65912
rect 10100 65900 10106 65952
rect 1104 65850 10856 65872
rect 1104 65798 2582 65850
rect 2634 65798 2646 65850
rect 2698 65798 2710 65850
rect 2762 65798 2774 65850
rect 2826 65798 2838 65850
rect 2890 65798 5845 65850
rect 5897 65798 5909 65850
rect 5961 65798 5973 65850
rect 6025 65798 6037 65850
rect 6089 65798 6101 65850
rect 6153 65798 9109 65850
rect 9161 65798 9173 65850
rect 9225 65798 9237 65850
rect 9289 65798 9301 65850
rect 9353 65798 9365 65850
rect 9417 65798 10856 65850
rect 1104 65776 10856 65798
rect 3050 65696 3056 65748
rect 3108 65736 3114 65748
rect 10965 65739 11023 65745
rect 10965 65736 10977 65739
rect 3108 65708 10977 65736
rect 3108 65696 3114 65708
rect 10965 65705 10977 65708
rect 11011 65705 11023 65739
rect 10965 65699 11023 65705
rect 1397 65671 1455 65677
rect 1397 65637 1409 65671
rect 1443 65668 1455 65671
rect 9030 65668 9036 65680
rect 1443 65640 9036 65668
rect 1443 65637 1455 65640
rect 1397 65631 1455 65637
rect 9030 65628 9036 65640
rect 9088 65628 9094 65680
rect 9582 65560 9588 65612
rect 9640 65600 9646 65612
rect 9640 65572 9720 65600
rect 9640 65560 9646 65572
rect 1578 65532 1584 65544
rect 1539 65504 1584 65532
rect 1578 65492 1584 65504
rect 1636 65492 1642 65544
rect 2222 65532 2228 65544
rect 2183 65504 2228 65532
rect 2222 65492 2228 65504
rect 2280 65492 2286 65544
rect 6730 65492 6736 65544
rect 6788 65532 6794 65544
rect 9401 65535 9459 65541
rect 9401 65532 9413 65535
rect 6788 65504 9413 65532
rect 6788 65492 6794 65504
rect 9401 65501 9413 65504
rect 9447 65501 9459 65535
rect 9401 65495 9459 65501
rect 9490 65492 9496 65544
rect 9548 65532 9554 65544
rect 9692 65541 9720 65572
rect 9677 65535 9735 65541
rect 9548 65504 9593 65532
rect 9548 65492 9554 65504
rect 9677 65501 9689 65535
rect 9723 65501 9735 65535
rect 9677 65495 9735 65501
rect 6546 65424 6552 65476
rect 6604 65464 6610 65476
rect 9858 65464 9864 65476
rect 6604 65436 9864 65464
rect 6604 65424 6610 65436
rect 9858 65424 9864 65436
rect 9916 65424 9922 65476
rect 10137 65467 10195 65473
rect 10137 65433 10149 65467
rect 10183 65464 10195 65467
rect 10594 65464 10600 65476
rect 10183 65436 10600 65464
rect 10183 65433 10195 65436
rect 10137 65427 10195 65433
rect 10594 65424 10600 65436
rect 10652 65424 10658 65476
rect 2041 65399 2099 65405
rect 2041 65365 2053 65399
rect 2087 65396 2099 65399
rect 8938 65396 8944 65408
rect 2087 65368 8944 65396
rect 2087 65365 2099 65368
rect 2041 65359 2099 65365
rect 8938 65356 8944 65368
rect 8996 65356 9002 65408
rect 1104 65306 10856 65328
rect 1104 65254 4213 65306
rect 4265 65254 4277 65306
rect 4329 65254 4341 65306
rect 4393 65254 4405 65306
rect 4457 65254 4469 65306
rect 4521 65254 7477 65306
rect 7529 65254 7541 65306
rect 7593 65254 7605 65306
rect 7657 65254 7669 65306
rect 7721 65254 7733 65306
rect 7785 65254 10856 65306
rect 1104 65232 10856 65254
rect 7285 65195 7343 65201
rect 7285 65161 7297 65195
rect 7331 65161 7343 65195
rect 7285 65155 7343 65161
rect 7300 65124 7328 65155
rect 7374 65152 7380 65204
rect 7432 65192 7438 65204
rect 7653 65195 7711 65201
rect 7653 65192 7665 65195
rect 7432 65164 7665 65192
rect 7432 65152 7438 65164
rect 7653 65161 7665 65164
rect 7699 65161 7711 65195
rect 7653 65155 7711 65161
rect 8573 65195 8631 65201
rect 8573 65161 8585 65195
rect 8619 65192 8631 65195
rect 9490 65192 9496 65204
rect 8619 65164 9496 65192
rect 8619 65161 8631 65164
rect 8573 65155 8631 65161
rect 9490 65152 9496 65164
rect 9548 65152 9554 65204
rect 11149 65127 11207 65133
rect 11149 65124 11161 65127
rect 7300 65096 11161 65124
rect 11149 65093 11161 65096
rect 11195 65093 11207 65127
rect 11149 65087 11207 65093
rect 1854 65056 1860 65068
rect 1815 65028 1860 65056
rect 1854 65016 1860 65028
rect 1912 65016 1918 65068
rect 7745 65059 7803 65065
rect 7745 65025 7757 65059
rect 7791 65056 7803 65059
rect 8110 65056 8116 65068
rect 7791 65028 8116 65056
rect 7791 65025 7803 65028
rect 7745 65019 7803 65025
rect 8110 65016 8116 65028
rect 8168 65016 8174 65068
rect 8754 65056 8760 65068
rect 8715 65028 8760 65056
rect 8754 65016 8760 65028
rect 8812 65016 8818 65068
rect 9401 65059 9459 65065
rect 9401 65025 9413 65059
rect 9447 65056 9459 65059
rect 9582 65056 9588 65068
rect 9447 65028 9588 65056
rect 9447 65025 9459 65028
rect 9401 65019 9459 65025
rect 9582 65016 9588 65028
rect 9640 65016 9646 65068
rect 9858 65056 9864 65068
rect 9819 65028 9864 65056
rect 9858 65016 9864 65028
rect 9916 65016 9922 65068
rect 7837 64991 7895 64997
rect 7837 64957 7849 64991
rect 7883 64957 7895 64991
rect 7837 64951 7895 64957
rect 8481 64991 8539 64997
rect 8481 64957 8493 64991
rect 8527 64988 8539 64991
rect 11241 64991 11299 64997
rect 11241 64988 11253 64991
rect 8527 64960 11253 64988
rect 8527 64957 8539 64960
rect 8481 64951 8539 64957
rect 11241 64957 11253 64960
rect 11287 64957 11299 64991
rect 11241 64951 11299 64957
rect 7852 64920 7880 64951
rect 9674 64920 9680 64932
rect 7852 64892 9680 64920
rect 9674 64880 9680 64892
rect 9732 64880 9738 64932
rect 10042 64920 10048 64932
rect 10003 64892 10048 64920
rect 10042 64880 10048 64892
rect 10100 64880 10106 64932
rect 1949 64855 2007 64861
rect 1949 64821 1961 64855
rect 1995 64852 2007 64855
rect 8481 64855 8539 64861
rect 8481 64852 8493 64855
rect 1995 64824 8493 64852
rect 1995 64821 2007 64824
rect 1949 64815 2007 64821
rect 8481 64821 8493 64824
rect 8527 64821 8539 64855
rect 8481 64815 8539 64821
rect 9217 64855 9275 64861
rect 9217 64821 9229 64855
rect 9263 64852 9275 64855
rect 9490 64852 9496 64864
rect 9263 64824 9496 64852
rect 9263 64821 9275 64824
rect 9217 64815 9275 64821
rect 9490 64812 9496 64824
rect 9548 64812 9554 64864
rect 1104 64762 10856 64784
rect 1104 64710 2582 64762
rect 2634 64710 2646 64762
rect 2698 64710 2710 64762
rect 2762 64710 2774 64762
rect 2826 64710 2838 64762
rect 2890 64710 5845 64762
rect 5897 64710 5909 64762
rect 5961 64710 5973 64762
rect 6025 64710 6037 64762
rect 6089 64710 6101 64762
rect 6153 64710 9109 64762
rect 9161 64710 9173 64762
rect 9225 64710 9237 64762
rect 9289 64710 9301 64762
rect 9353 64710 9365 64762
rect 9417 64710 10856 64762
rect 1104 64688 10856 64710
rect 1394 64444 1400 64456
rect 1355 64416 1400 64444
rect 1394 64404 1400 64416
rect 1452 64404 1458 64456
rect 8386 64404 8392 64456
rect 8444 64444 8450 64456
rect 9401 64447 9459 64453
rect 9401 64444 9413 64447
rect 8444 64416 9413 64444
rect 8444 64404 8450 64416
rect 9401 64413 9413 64416
rect 9447 64413 9459 64447
rect 9401 64407 9459 64413
rect 9490 64404 9496 64456
rect 9548 64444 9554 64456
rect 9548 64416 9593 64444
rect 9548 64404 9554 64416
rect 9674 64404 9680 64456
rect 9732 64444 9738 64456
rect 9732 64416 9777 64444
rect 9732 64404 9738 64416
rect 9692 64376 9720 64404
rect 9508 64348 9720 64376
rect 10137 64379 10195 64385
rect 9508 64320 9536 64348
rect 10137 64345 10149 64379
rect 10183 64376 10195 64379
rect 10410 64376 10416 64388
rect 10183 64348 10416 64376
rect 10183 64345 10195 64348
rect 10137 64339 10195 64345
rect 10410 64336 10416 64348
rect 10468 64336 10474 64388
rect 1581 64311 1639 64317
rect 1581 64277 1593 64311
rect 1627 64308 1639 64311
rect 8846 64308 8852 64320
rect 1627 64280 8852 64308
rect 1627 64277 1639 64280
rect 1581 64271 1639 64277
rect 8846 64268 8852 64280
rect 8904 64268 8910 64320
rect 9490 64268 9496 64320
rect 9548 64268 9554 64320
rect 1104 64218 10856 64240
rect 1104 64166 4213 64218
rect 4265 64166 4277 64218
rect 4329 64166 4341 64218
rect 4393 64166 4405 64218
rect 4457 64166 4469 64218
rect 4521 64166 7477 64218
rect 7529 64166 7541 64218
rect 7593 64166 7605 64218
rect 7657 64166 7669 64218
rect 7721 64166 7733 64218
rect 7785 64166 10856 64218
rect 1104 64144 10856 64166
rect 9030 64064 9036 64116
rect 9088 64104 9094 64116
rect 9125 64107 9183 64113
rect 9125 64104 9137 64107
rect 9088 64076 9137 64104
rect 9088 64064 9094 64076
rect 9125 64073 9137 64076
rect 9171 64073 9183 64107
rect 9125 64067 9183 64073
rect 9217 64039 9275 64045
rect 9217 64005 9229 64039
rect 9263 64036 9275 64039
rect 11149 64039 11207 64045
rect 11149 64036 11161 64039
rect 9263 64008 11161 64036
rect 9263 64005 9275 64008
rect 9217 63999 9275 64005
rect 11149 64005 11161 64008
rect 11195 64005 11207 64039
rect 11149 63999 11207 64005
rect 1026 63928 1032 63980
rect 1084 63968 1090 63980
rect 1397 63971 1455 63977
rect 1397 63968 1409 63971
rect 1084 63940 1409 63968
rect 1084 63928 1090 63940
rect 1397 63937 1409 63940
rect 1443 63937 1455 63971
rect 10134 63968 10140 63980
rect 10095 63940 10140 63968
rect 1397 63931 1455 63937
rect 10134 63928 10140 63940
rect 10192 63928 10198 63980
rect 9401 63903 9459 63909
rect 9401 63869 9413 63903
rect 9447 63900 9459 63903
rect 9582 63900 9588 63912
rect 9447 63872 9588 63900
rect 9447 63869 9459 63872
rect 9401 63863 9459 63869
rect 9582 63860 9588 63872
rect 9640 63860 9646 63912
rect 11057 63903 11115 63909
rect 11057 63869 11069 63903
rect 11103 63869 11115 63903
rect 11057 63863 11115 63869
rect 8757 63835 8815 63841
rect 8757 63801 8769 63835
rect 8803 63832 8815 63835
rect 11072 63832 11100 63863
rect 8803 63804 11100 63832
rect 8803 63801 8815 63804
rect 8757 63795 8815 63801
rect 1581 63767 1639 63773
rect 1581 63733 1593 63767
rect 1627 63764 1639 63767
rect 1762 63764 1768 63776
rect 1627 63736 1768 63764
rect 1627 63733 1639 63736
rect 1581 63727 1639 63733
rect 1762 63724 1768 63736
rect 1820 63724 1826 63776
rect 9953 63767 10011 63773
rect 9953 63733 9965 63767
rect 9999 63764 10011 63767
rect 10965 63767 11023 63773
rect 10965 63764 10977 63767
rect 9999 63736 10977 63764
rect 9999 63733 10011 63736
rect 9953 63727 10011 63733
rect 10965 63733 10977 63736
rect 11011 63733 11023 63767
rect 10965 63727 11023 63733
rect 1104 63674 10856 63696
rect 1104 63622 2582 63674
rect 2634 63622 2646 63674
rect 2698 63622 2710 63674
rect 2762 63622 2774 63674
rect 2826 63622 2838 63674
rect 2890 63622 5845 63674
rect 5897 63622 5909 63674
rect 5961 63622 5973 63674
rect 6025 63622 6037 63674
rect 6089 63622 6101 63674
rect 6153 63622 9109 63674
rect 9161 63622 9173 63674
rect 9225 63622 9237 63674
rect 9289 63622 9301 63674
rect 9353 63622 9365 63674
rect 9417 63622 10856 63674
rect 1104 63600 10856 63622
rect 2590 63492 2596 63504
rect 2551 63464 2596 63492
rect 2590 63452 2596 63464
rect 2648 63452 2654 63504
rect 2958 63424 2964 63436
rect 2919 63396 2964 63424
rect 2958 63384 2964 63396
rect 3016 63384 3022 63436
rect 3145 63427 3203 63433
rect 3145 63393 3157 63427
rect 3191 63424 3203 63427
rect 3602 63424 3608 63436
rect 3191 63396 3608 63424
rect 3191 63393 3203 63396
rect 3145 63387 3203 63393
rect 1394 63356 1400 63368
rect 1355 63328 1400 63356
rect 1394 63316 1400 63328
rect 1452 63316 1458 63368
rect 2498 63316 2504 63368
rect 2556 63356 2562 63368
rect 3160 63356 3188 63387
rect 3602 63384 3608 63396
rect 3660 63384 3666 63436
rect 9490 63356 9496 63368
rect 2556 63328 3188 63356
rect 9451 63328 9496 63356
rect 2556 63316 2562 63328
rect 9490 63316 9496 63328
rect 9548 63316 9554 63368
rect 10137 63359 10195 63365
rect 10137 63325 10149 63359
rect 10183 63356 10195 63359
rect 10226 63356 10232 63368
rect 10183 63328 10232 63356
rect 10183 63325 10195 63328
rect 10137 63319 10195 63325
rect 10226 63316 10232 63328
rect 10284 63316 10290 63368
rect 6454 63288 6460 63300
rect 2746 63260 6460 63288
rect 1581 63223 1639 63229
rect 1581 63189 1593 63223
rect 1627 63220 1639 63223
rect 2746 63220 2774 63260
rect 6454 63248 6460 63260
rect 6512 63248 6518 63300
rect 1627 63192 2774 63220
rect 3053 63223 3111 63229
rect 1627 63189 1639 63192
rect 1581 63183 1639 63189
rect 3053 63189 3065 63223
rect 3099 63220 3111 63223
rect 3142 63220 3148 63232
rect 3099 63192 3148 63220
rect 3099 63189 3111 63192
rect 3053 63183 3111 63189
rect 3142 63180 3148 63192
rect 3200 63180 3206 63232
rect 9309 63223 9367 63229
rect 9309 63189 9321 63223
rect 9355 63220 9367 63223
rect 9490 63220 9496 63232
rect 9355 63192 9496 63220
rect 9355 63189 9367 63192
rect 9309 63183 9367 63189
rect 9490 63180 9496 63192
rect 9548 63180 9554 63232
rect 9953 63223 10011 63229
rect 9953 63189 9965 63223
rect 9999 63220 10011 63223
rect 11517 63223 11575 63229
rect 11517 63220 11529 63223
rect 9999 63192 11529 63220
rect 9999 63189 10011 63192
rect 9953 63183 10011 63189
rect 11517 63189 11529 63192
rect 11563 63189 11575 63223
rect 11517 63183 11575 63189
rect 1104 63130 10856 63152
rect 1104 63078 4213 63130
rect 4265 63078 4277 63130
rect 4329 63078 4341 63130
rect 4393 63078 4405 63130
rect 4457 63078 4469 63130
rect 4521 63078 7477 63130
rect 7529 63078 7541 63130
rect 7593 63078 7605 63130
rect 7657 63078 7669 63130
rect 7721 63078 7733 63130
rect 7785 63078 10856 63130
rect 1104 63056 10856 63078
rect 2314 63016 2320 63028
rect 2275 62988 2320 63016
rect 2314 62976 2320 62988
rect 2372 62976 2378 63028
rect 7374 62976 7380 63028
rect 7432 63016 7438 63028
rect 7837 63019 7895 63025
rect 7837 63016 7849 63019
rect 7432 62988 7849 63016
rect 7432 62976 7438 62988
rect 7837 62985 7849 62988
rect 7883 62985 7895 63019
rect 7837 62979 7895 62985
rect 9030 62976 9036 63028
rect 9088 63016 9094 63028
rect 9309 63019 9367 63025
rect 9309 63016 9321 63019
rect 9088 62988 9321 63016
rect 9088 62976 9094 62988
rect 9309 62985 9321 62988
rect 9355 62985 9367 63019
rect 9309 62979 9367 62985
rect 11885 62951 11943 62957
rect 11885 62948 11897 62951
rect 2746 62920 11897 62948
rect 2222 62772 2228 62824
rect 2280 62812 2286 62824
rect 2409 62815 2467 62821
rect 2409 62812 2421 62815
rect 2280 62784 2421 62812
rect 2280 62772 2286 62784
rect 2409 62781 2421 62784
rect 2455 62781 2467 62815
rect 2409 62775 2467 62781
rect 2498 62772 2504 62824
rect 2556 62812 2562 62824
rect 2556 62784 2601 62812
rect 2556 62772 2562 62784
rect 1949 62747 2007 62753
rect 1949 62713 1961 62747
rect 1995 62744 2007 62747
rect 2746 62744 2774 62920
rect 11885 62917 11897 62920
rect 11931 62917 11943 62951
rect 11885 62911 11943 62917
rect 9401 62883 9459 62889
rect 9401 62880 9413 62883
rect 8496 62852 9413 62880
rect 8496 62824 8524 62852
rect 9401 62849 9413 62852
rect 9447 62880 9459 62883
rect 9582 62880 9588 62892
rect 9447 62852 9588 62880
rect 9447 62849 9459 62852
rect 9401 62843 9459 62849
rect 9582 62840 9588 62852
rect 9640 62840 9646 62892
rect 10134 62880 10140 62892
rect 10095 62852 10140 62880
rect 10134 62840 10140 62852
rect 10192 62840 10198 62892
rect 7837 62815 7895 62821
rect 7837 62781 7849 62815
rect 7883 62781 7895 62815
rect 7837 62775 7895 62781
rect 7929 62815 7987 62821
rect 7929 62781 7941 62815
rect 7975 62812 7987 62815
rect 8478 62812 8484 62824
rect 7975 62784 8484 62812
rect 7975 62781 7987 62784
rect 7929 62775 7987 62781
rect 1995 62716 2774 62744
rect 1995 62713 2007 62716
rect 1949 62707 2007 62713
rect 6178 62704 6184 62756
rect 6236 62744 6242 62756
rect 7852 62744 7880 62775
rect 8478 62772 8484 62784
rect 8536 62772 8542 62824
rect 9309 62815 9367 62821
rect 9309 62781 9321 62815
rect 9355 62812 9367 62815
rect 11149 62815 11207 62821
rect 11149 62812 11161 62815
rect 9355 62784 11161 62812
rect 9355 62781 9367 62784
rect 9309 62775 9367 62781
rect 11149 62781 11161 62784
rect 11195 62781 11207 62815
rect 11149 62775 11207 62781
rect 11241 62815 11299 62821
rect 11241 62781 11253 62815
rect 11287 62812 11299 62815
rect 11422 62812 11428 62824
rect 11287 62784 11428 62812
rect 11287 62781 11299 62784
rect 11241 62775 11299 62781
rect 11422 62772 11428 62784
rect 11480 62772 11486 62824
rect 8110 62744 8116 62756
rect 6236 62716 7512 62744
rect 7852 62716 8116 62744
rect 6236 62704 6242 62716
rect 7374 62676 7380 62688
rect 7335 62648 7380 62676
rect 7374 62636 7380 62648
rect 7432 62636 7438 62688
rect 7484 62676 7512 62716
rect 8110 62704 8116 62716
rect 8168 62704 8174 62756
rect 8849 62679 8907 62685
rect 8849 62676 8861 62679
rect 7484 62648 8861 62676
rect 8849 62645 8861 62648
rect 8895 62645 8907 62679
rect 8849 62639 8907 62645
rect 9953 62679 10011 62685
rect 9953 62645 9965 62679
rect 9999 62676 10011 62679
rect 11241 62679 11299 62685
rect 11241 62676 11253 62679
rect 9999 62648 11253 62676
rect 9999 62645 10011 62648
rect 9953 62639 10011 62645
rect 11241 62645 11253 62648
rect 11287 62645 11299 62679
rect 11241 62639 11299 62645
rect 1104 62586 10856 62608
rect 1104 62534 2582 62586
rect 2634 62534 2646 62586
rect 2698 62534 2710 62586
rect 2762 62534 2774 62586
rect 2826 62534 2838 62586
rect 2890 62534 5845 62586
rect 5897 62534 5909 62586
rect 5961 62534 5973 62586
rect 6025 62534 6037 62586
rect 6089 62534 6101 62586
rect 6153 62534 9109 62586
rect 9161 62534 9173 62586
rect 9225 62534 9237 62586
rect 9289 62534 9301 62586
rect 9353 62534 9365 62586
rect 9417 62534 10856 62586
rect 1104 62512 10856 62534
rect 7653 62475 7711 62481
rect 7653 62441 7665 62475
rect 7699 62472 7711 62475
rect 8662 62472 8668 62484
rect 7699 62444 8668 62472
rect 7699 62441 7711 62444
rect 7653 62435 7711 62441
rect 8662 62432 8668 62444
rect 8720 62432 8726 62484
rect 11057 62407 11115 62413
rect 11057 62373 11069 62407
rect 11103 62404 11115 62407
rect 11238 62404 11244 62416
rect 11103 62376 11244 62404
rect 11103 62373 11115 62376
rect 11057 62367 11115 62373
rect 11238 62364 11244 62376
rect 11296 62364 11302 62416
rect 8297 62339 8355 62345
rect 8297 62305 8309 62339
rect 8343 62336 8355 62339
rect 8478 62336 8484 62348
rect 8343 62308 8484 62336
rect 8343 62305 8355 62308
rect 8297 62299 8355 62305
rect 8478 62296 8484 62308
rect 8536 62296 8542 62348
rect 7098 62228 7104 62280
rect 7156 62268 7162 62280
rect 8021 62271 8079 62277
rect 8021 62268 8033 62271
rect 7156 62240 8033 62268
rect 7156 62228 7162 62240
rect 8021 62237 8033 62240
rect 8067 62237 8079 62271
rect 9306 62268 9312 62280
rect 9267 62240 9312 62268
rect 8021 62231 8079 62237
rect 9306 62228 9312 62240
rect 9364 62228 9370 62280
rect 9585 62271 9643 62277
rect 9585 62237 9597 62271
rect 9631 62268 9643 62271
rect 11057 62271 11115 62277
rect 11057 62268 11069 62271
rect 9631 62240 11069 62268
rect 9631 62237 9643 62240
rect 9585 62231 9643 62237
rect 11057 62237 11069 62240
rect 11103 62237 11115 62271
rect 11057 62231 11115 62237
rect 1854 62200 1860 62212
rect 1815 62172 1860 62200
rect 1854 62160 1860 62172
rect 1912 62160 1918 62212
rect 2041 62203 2099 62209
rect 2041 62169 2053 62203
rect 2087 62200 2099 62203
rect 3510 62200 3516 62212
rect 2087 62172 3516 62200
rect 2087 62169 2099 62172
rect 2041 62163 2099 62169
rect 3510 62160 3516 62172
rect 3568 62160 3574 62212
rect 8113 62135 8171 62141
rect 8113 62101 8125 62135
rect 8159 62132 8171 62135
rect 8202 62132 8208 62144
rect 8159 62104 8208 62132
rect 8159 62101 8171 62104
rect 8113 62095 8171 62101
rect 8202 62092 8208 62104
rect 8260 62092 8266 62144
rect 1104 62042 10856 62064
rect 1104 61990 4213 62042
rect 4265 61990 4277 62042
rect 4329 61990 4341 62042
rect 4393 61990 4405 62042
rect 4457 61990 4469 62042
rect 4521 61990 7477 62042
rect 7529 61990 7541 62042
rect 7593 61990 7605 62042
rect 7657 61990 7669 62042
rect 7721 61990 7733 62042
rect 7785 61990 10856 62042
rect 1104 61968 10856 61990
rect 1394 61752 1400 61804
rect 1452 61792 1458 61804
rect 1857 61795 1915 61801
rect 1857 61792 1869 61795
rect 1452 61764 1869 61792
rect 1452 61752 1458 61764
rect 1857 61761 1869 61764
rect 1903 61761 1915 61795
rect 1857 61755 1915 61761
rect 9309 61727 9367 61733
rect 9309 61693 9321 61727
rect 9355 61693 9367 61727
rect 9309 61687 9367 61693
rect 9585 61727 9643 61733
rect 9585 61693 9597 61727
rect 9631 61724 9643 61727
rect 11885 61727 11943 61733
rect 11885 61724 11897 61727
rect 9631 61696 11897 61724
rect 9631 61693 9643 61696
rect 9585 61687 9643 61693
rect 11885 61693 11897 61696
rect 11931 61693 11943 61727
rect 11885 61687 11943 61693
rect 2041 61659 2099 61665
rect 2041 61625 2053 61659
rect 2087 61656 2099 61659
rect 3602 61656 3608 61668
rect 2087 61628 3608 61656
rect 2087 61625 2099 61628
rect 2041 61619 2099 61625
rect 3602 61616 3608 61628
rect 3660 61616 3666 61668
rect 9324 61588 9352 61687
rect 9582 61588 9588 61600
rect 9324 61560 9588 61588
rect 9582 61548 9588 61560
rect 9640 61548 9646 61600
rect 1104 61498 10856 61520
rect 1104 61446 2582 61498
rect 2634 61446 2646 61498
rect 2698 61446 2710 61498
rect 2762 61446 2774 61498
rect 2826 61446 2838 61498
rect 2890 61446 5845 61498
rect 5897 61446 5909 61498
rect 5961 61446 5973 61498
rect 6025 61446 6037 61498
rect 6089 61446 6101 61498
rect 6153 61446 9109 61498
rect 9161 61446 9173 61498
rect 9225 61446 9237 61498
rect 9289 61446 9301 61498
rect 9353 61446 9365 61498
rect 9417 61446 10856 61498
rect 1104 61424 10856 61446
rect 2222 61248 2228 61260
rect 2135 61220 2228 61248
rect 2222 61208 2228 61220
rect 2280 61248 2286 61260
rect 5350 61248 5356 61260
rect 2280 61220 5356 61248
rect 2280 61208 2286 61220
rect 5350 61208 5356 61220
rect 5408 61208 5414 61260
rect 2314 61140 2320 61192
rect 2372 61180 2378 61192
rect 2372 61152 2417 61180
rect 2372 61140 2378 61152
rect 2498 61140 2504 61192
rect 2556 61180 2562 61192
rect 9398 61180 9404 61192
rect 2556 61152 2601 61180
rect 9359 61152 9404 61180
rect 2556 61140 2562 61152
rect 9398 61140 9404 61152
rect 9456 61140 9462 61192
rect 9490 61140 9496 61192
rect 9548 61180 9554 61192
rect 9548 61152 9593 61180
rect 9548 61140 9554 61152
rect 9674 61140 9680 61192
rect 9732 61180 9738 61192
rect 9732 61152 9777 61180
rect 9732 61140 9738 61152
rect 2961 61115 3019 61121
rect 2961 61081 2973 61115
rect 3007 61112 3019 61115
rect 4982 61112 4988 61124
rect 3007 61084 4988 61112
rect 3007 61081 3019 61084
rect 2961 61075 3019 61081
rect 4982 61072 4988 61084
rect 5040 61072 5046 61124
rect 10137 61115 10195 61121
rect 10137 61081 10149 61115
rect 10183 61112 10195 61115
rect 10502 61112 10508 61124
rect 10183 61084 10508 61112
rect 10183 61081 10195 61084
rect 10137 61075 10195 61081
rect 10502 61072 10508 61084
rect 10560 61072 10566 61124
rect 11330 61044 11336 61056
rect 11291 61016 11336 61044
rect 11330 61004 11336 61016
rect 11388 61004 11394 61056
rect 1104 60954 10856 60976
rect 1104 60902 4213 60954
rect 4265 60902 4277 60954
rect 4329 60902 4341 60954
rect 4393 60902 4405 60954
rect 4457 60902 4469 60954
rect 4521 60902 7477 60954
rect 7529 60902 7541 60954
rect 7593 60902 7605 60954
rect 7657 60902 7669 60954
rect 7721 60902 7733 60954
rect 7785 60902 10856 60954
rect 10962 60936 10968 60988
rect 11020 60976 11026 60988
rect 11149 60979 11207 60985
rect 11149 60976 11161 60979
rect 11020 60948 11161 60976
rect 11020 60936 11026 60948
rect 11149 60945 11161 60948
rect 11195 60945 11207 60979
rect 11149 60939 11207 60945
rect 11425 60979 11483 60985
rect 11425 60945 11437 60979
rect 11471 60945 11483 60979
rect 11425 60939 11483 60945
rect 1104 60880 10856 60902
rect 11057 60911 11115 60917
rect 11057 60877 11069 60911
rect 11103 60877 11115 60911
rect 11440 60908 11468 60939
rect 11057 60871 11115 60877
rect 11164 60880 11468 60908
rect 2038 60840 2044 60852
rect 1999 60812 2044 60840
rect 2038 60800 2044 60812
rect 2096 60800 2102 60852
rect 8110 60800 8116 60852
rect 8168 60840 8174 60852
rect 8294 60840 8300 60852
rect 8168 60812 8300 60840
rect 8168 60800 8174 60812
rect 8294 60800 8300 60812
rect 8352 60800 8358 60852
rect 2133 60775 2191 60781
rect 2133 60741 2145 60775
rect 2179 60772 2191 60775
rect 2498 60772 2504 60784
rect 2179 60744 2504 60772
rect 2179 60741 2191 60744
rect 2133 60735 2191 60741
rect 2498 60732 2504 60744
rect 2556 60732 2562 60784
rect 8662 60772 8668 60784
rect 8623 60744 8668 60772
rect 8662 60732 8668 60744
rect 8720 60732 8726 60784
rect 2774 60664 2780 60716
rect 2832 60704 2838 60716
rect 9306 60704 9312 60716
rect 2832 60676 2877 60704
rect 9267 60676 9312 60704
rect 2832 60664 2838 60676
rect 9306 60664 9312 60676
rect 9364 60664 9370 60716
rect 11072 60704 11100 60871
rect 11164 60849 11192 60880
rect 11149 60843 11207 60849
rect 11149 60809 11161 60843
rect 11195 60809 11207 60843
rect 11422 60840 11428 60852
rect 11383 60812 11428 60840
rect 11149 60803 11207 60809
rect 11422 60800 11428 60812
rect 11480 60800 11486 60852
rect 11609 60843 11667 60849
rect 11609 60809 11621 60843
rect 11655 60809 11667 60843
rect 11790 60840 11796 60852
rect 11751 60812 11796 60840
rect 11609 60803 11667 60809
rect 11238 60732 11244 60784
rect 11296 60772 11302 60784
rect 11624 60772 11652 60803
rect 11790 60800 11796 60812
rect 11848 60800 11854 60852
rect 11296 60744 11341 60772
rect 11624 60744 11836 60772
rect 11296 60732 11302 60744
rect 11808 60713 11836 60744
rect 11609 60707 11667 60713
rect 11609 60704 11621 60707
rect 11072 60676 11621 60704
rect 11609 60673 11621 60676
rect 11655 60673 11667 60707
rect 11609 60667 11667 60673
rect 11793 60707 11851 60713
rect 11793 60673 11805 60707
rect 11839 60673 11851 60707
rect 11793 60667 11851 60673
rect 1670 60596 1676 60648
rect 1728 60636 1734 60648
rect 2038 60636 2044 60648
rect 1728 60608 2044 60636
rect 1728 60596 1734 60608
rect 2038 60596 2044 60608
rect 2096 60596 2102 60648
rect 9585 60639 9643 60645
rect 9585 60605 9597 60639
rect 9631 60636 9643 60639
rect 10226 60636 10232 60648
rect 9631 60608 10232 60636
rect 9631 60605 9643 60608
rect 9585 60599 9643 60605
rect 10226 60596 10232 60608
rect 10284 60596 10290 60648
rect 10962 60596 10968 60648
rect 11020 60636 11026 60648
rect 11057 60639 11115 60645
rect 11057 60636 11069 60639
rect 11020 60608 11069 60636
rect 11020 60596 11026 60608
rect 11057 60605 11069 60608
rect 11103 60605 11115 60639
rect 11057 60599 11115 60605
rect 2961 60571 3019 60577
rect 2961 60537 2973 60571
rect 3007 60568 3019 60571
rect 3970 60568 3976 60580
rect 3007 60540 3976 60568
rect 3007 60537 3019 60540
rect 2961 60531 3019 60537
rect 3970 60528 3976 60540
rect 4028 60528 4034 60580
rect 1578 60500 1584 60512
rect 1539 60472 1584 60500
rect 1578 60460 1584 60472
rect 1636 60460 1642 60512
rect 8754 60500 8760 60512
rect 8715 60472 8760 60500
rect 8754 60460 8760 60472
rect 8812 60460 8818 60512
rect 1104 60410 10856 60432
rect 1104 60358 2582 60410
rect 2634 60358 2646 60410
rect 2698 60358 2710 60410
rect 2762 60358 2774 60410
rect 2826 60358 2838 60410
rect 2890 60358 5845 60410
rect 5897 60358 5909 60410
rect 5961 60358 5973 60410
rect 6025 60358 6037 60410
rect 6089 60358 6101 60410
rect 6153 60358 9109 60410
rect 9161 60358 9173 60410
rect 9225 60358 9237 60410
rect 9289 60358 9301 60410
rect 9353 60358 9365 60410
rect 9417 60358 10856 60410
rect 1104 60336 10856 60358
rect 11514 60296 11520 60308
rect 11475 60268 11520 60296
rect 11514 60256 11520 60268
rect 11572 60256 11578 60308
rect 7098 60188 7104 60240
rect 7156 60228 7162 60240
rect 7745 60231 7803 60237
rect 7745 60228 7757 60231
rect 7156 60200 7757 60228
rect 7156 60188 7162 60200
rect 7745 60197 7757 60200
rect 7791 60197 7803 60231
rect 7745 60191 7803 60197
rect 8202 60160 8208 60172
rect 8163 60132 8208 60160
rect 8202 60120 8208 60132
rect 8260 60120 8266 60172
rect 8297 60163 8355 60169
rect 8297 60129 8309 60163
rect 8343 60160 8355 60163
rect 8478 60160 8484 60172
rect 8343 60132 8484 60160
rect 8343 60129 8355 60132
rect 8297 60123 8355 60129
rect 8478 60120 8484 60132
rect 8536 60120 8542 60172
rect 11149 60163 11207 60169
rect 11149 60129 11161 60163
rect 11195 60160 11207 60163
rect 11517 60163 11575 60169
rect 11517 60160 11529 60163
rect 11195 60132 11529 60160
rect 11195 60129 11207 60132
rect 11149 60123 11207 60129
rect 11517 60129 11529 60132
rect 11563 60129 11575 60163
rect 11517 60123 11575 60129
rect 9953 60095 10011 60101
rect 9953 60061 9965 60095
rect 9999 60092 10011 60095
rect 10042 60092 10048 60104
rect 9999 60064 10048 60092
rect 9999 60061 10011 60064
rect 9953 60055 10011 60061
rect 10042 60052 10048 60064
rect 10100 60052 10106 60104
rect 1854 60024 1860 60036
rect 1815 59996 1860 60024
rect 1854 59984 1860 59996
rect 1912 59984 1918 60036
rect 10137 60027 10195 60033
rect 10137 59993 10149 60027
rect 10183 60024 10195 60027
rect 11149 60027 11207 60033
rect 11149 60024 11161 60027
rect 10183 59996 11161 60024
rect 10183 59993 10195 59996
rect 10137 59987 10195 59993
rect 11149 59993 11161 59996
rect 11195 59993 11207 60027
rect 11149 59987 11207 59993
rect 842 59916 848 59968
rect 900 59956 906 59968
rect 1949 59959 2007 59965
rect 1949 59956 1961 59959
rect 900 59928 1961 59956
rect 900 59916 906 59928
rect 1949 59925 1961 59928
rect 1995 59925 2007 59959
rect 1949 59919 2007 59925
rect 7190 59916 7196 59968
rect 7248 59956 7254 59968
rect 8205 59959 8263 59965
rect 8205 59956 8217 59959
rect 7248 59928 8217 59956
rect 7248 59916 7254 59928
rect 8205 59925 8217 59928
rect 8251 59925 8263 59959
rect 8205 59919 8263 59925
rect 1104 59866 10856 59888
rect 1104 59814 4213 59866
rect 4265 59814 4277 59866
rect 4329 59814 4341 59866
rect 4393 59814 4405 59866
rect 4457 59814 4469 59866
rect 4521 59814 7477 59866
rect 7529 59814 7541 59866
rect 7593 59814 7605 59866
rect 7657 59814 7669 59866
rect 7721 59814 7733 59866
rect 7785 59814 10856 59866
rect 1104 59792 10856 59814
rect 7190 59712 7196 59764
rect 7248 59752 7254 59764
rect 8202 59752 8208 59764
rect 7248 59724 8208 59752
rect 7248 59712 7254 59724
rect 8202 59712 8208 59724
rect 8260 59712 8266 59764
rect 9214 59684 9220 59696
rect 9175 59656 9220 59684
rect 9214 59644 9220 59656
rect 9272 59644 9278 59696
rect 1854 59616 1860 59628
rect 1815 59588 1860 59616
rect 1854 59576 1860 59588
rect 1912 59576 1918 59628
rect 9950 59616 9956 59628
rect 9911 59588 9956 59616
rect 9950 59576 9956 59588
rect 10008 59576 10014 59628
rect 10137 59483 10195 59489
rect 10137 59449 10149 59483
rect 10183 59480 10195 59483
rect 10778 59480 10784 59492
rect 10183 59452 10784 59480
rect 10183 59449 10195 59452
rect 10137 59443 10195 59449
rect 10778 59440 10784 59452
rect 10836 59440 10842 59492
rect 658 59372 664 59424
rect 716 59412 722 59424
rect 1949 59415 2007 59421
rect 1949 59412 1961 59415
rect 716 59384 1961 59412
rect 716 59372 722 59384
rect 1949 59381 1961 59384
rect 1995 59381 2007 59415
rect 1949 59375 2007 59381
rect 8478 59372 8484 59424
rect 8536 59412 8542 59424
rect 9309 59415 9367 59421
rect 9309 59412 9321 59415
rect 8536 59384 9321 59412
rect 8536 59372 8542 59384
rect 9309 59381 9321 59384
rect 9355 59381 9367 59415
rect 9309 59375 9367 59381
rect 1104 59322 10856 59344
rect 1104 59270 2582 59322
rect 2634 59270 2646 59322
rect 2698 59270 2710 59322
rect 2762 59270 2774 59322
rect 2826 59270 2838 59322
rect 2890 59270 5845 59322
rect 5897 59270 5909 59322
rect 5961 59270 5973 59322
rect 6025 59270 6037 59322
rect 6089 59270 6101 59322
rect 6153 59270 9109 59322
rect 9161 59270 9173 59322
rect 9225 59270 9237 59322
rect 9289 59270 9301 59322
rect 9353 59270 9365 59322
rect 9417 59270 10856 59322
rect 1104 59248 10856 59270
rect 11333 59143 11391 59149
rect 11333 59109 11345 59143
rect 11379 59140 11391 59143
rect 11701 59143 11759 59149
rect 11701 59140 11713 59143
rect 11379 59112 11713 59140
rect 11379 59109 11391 59112
rect 11333 59103 11391 59109
rect 11701 59109 11713 59112
rect 11747 59109 11759 59143
rect 11701 59103 11759 59109
rect 10137 59007 10195 59013
rect 10137 58973 10149 59007
rect 10183 59004 10195 59007
rect 11333 59007 11391 59013
rect 11333 59004 11345 59007
rect 10183 58976 11345 59004
rect 10183 58973 10195 58976
rect 10137 58967 10195 58973
rect 11333 58973 11345 58976
rect 11379 58973 11391 59007
rect 11333 58967 11391 58973
rect 9953 58939 10011 58945
rect 9953 58905 9965 58939
rect 9999 58936 10011 58939
rect 10226 58936 10232 58948
rect 9999 58908 10232 58936
rect 9999 58905 10011 58908
rect 9953 58899 10011 58905
rect 10226 58896 10232 58908
rect 10284 58896 10290 58948
rect 1104 58778 10856 58800
rect 1104 58726 4213 58778
rect 4265 58726 4277 58778
rect 4329 58726 4341 58778
rect 4393 58726 4405 58778
rect 4457 58726 4469 58778
rect 4521 58726 7477 58778
rect 7529 58726 7541 58778
rect 7593 58726 7605 58778
rect 7657 58726 7669 58778
rect 7721 58726 7733 58778
rect 7785 58726 10856 58778
rect 1104 58704 10856 58726
rect 3602 58624 3608 58676
rect 3660 58664 3666 58676
rect 3878 58664 3884 58676
rect 3660 58636 3884 58664
rect 3660 58624 3666 58636
rect 3878 58624 3884 58636
rect 3936 58624 3942 58676
rect 8294 58624 8300 58676
rect 8352 58664 8358 58676
rect 8846 58664 8852 58676
rect 8352 58636 8852 58664
rect 8352 58624 8358 58636
rect 8846 58624 8852 58636
rect 8904 58624 8910 58676
rect 1397 58531 1455 58537
rect 1397 58497 1409 58531
rect 1443 58528 1455 58531
rect 8846 58528 8852 58540
rect 1443 58500 8852 58528
rect 1443 58497 1455 58500
rect 1397 58491 1455 58497
rect 8846 58488 8852 58500
rect 8904 58488 8910 58540
rect 9950 58528 9956 58540
rect 9911 58500 9956 58528
rect 9950 58488 9956 58500
rect 10008 58488 10014 58540
rect 1578 58392 1584 58404
rect 1539 58364 1584 58392
rect 1578 58352 1584 58364
rect 1636 58352 1642 58404
rect 10137 58395 10195 58401
rect 10137 58361 10149 58395
rect 10183 58392 10195 58395
rect 11882 58392 11888 58404
rect 10183 58364 11888 58392
rect 10183 58361 10195 58364
rect 10137 58355 10195 58361
rect 11882 58352 11888 58364
rect 11940 58352 11946 58404
rect 1104 58234 10856 58256
rect 1104 58182 2582 58234
rect 2634 58182 2646 58234
rect 2698 58182 2710 58234
rect 2762 58182 2774 58234
rect 2826 58182 2838 58234
rect 2890 58182 5845 58234
rect 5897 58182 5909 58234
rect 5961 58182 5973 58234
rect 6025 58182 6037 58234
rect 6089 58182 6101 58234
rect 6153 58182 9109 58234
rect 9161 58182 9173 58234
rect 9225 58182 9237 58234
rect 9289 58182 9301 58234
rect 9353 58182 9365 58234
rect 9417 58182 10856 58234
rect 1104 58160 10856 58182
rect 1397 57919 1455 57925
rect 1397 57885 1409 57919
rect 1443 57916 1455 57919
rect 8662 57916 8668 57928
rect 1443 57888 8668 57916
rect 1443 57885 1455 57888
rect 1397 57879 1455 57885
rect 8662 57876 8668 57888
rect 8720 57876 8726 57928
rect 11698 57916 11704 57928
rect 9646 57888 11704 57916
rect 5258 57808 5264 57860
rect 5316 57848 5322 57860
rect 9646 57848 9674 57888
rect 11698 57876 11704 57888
rect 11756 57876 11762 57928
rect 5316 57820 9674 57848
rect 9953 57851 10011 57857
rect 5316 57808 5322 57820
rect 9953 57817 9965 57851
rect 9999 57848 10011 57851
rect 10318 57848 10324 57860
rect 9999 57820 10324 57848
rect 9999 57817 10011 57820
rect 9953 57811 10011 57817
rect 10318 57808 10324 57820
rect 10376 57808 10382 57860
rect 1578 57780 1584 57792
rect 1539 57752 1584 57780
rect 1578 57740 1584 57752
rect 1636 57740 1642 57792
rect 9769 57783 9827 57789
rect 9769 57749 9781 57783
rect 9815 57780 9827 57783
rect 10045 57783 10103 57789
rect 10045 57780 10057 57783
rect 9815 57752 10057 57780
rect 9815 57749 9827 57752
rect 9769 57743 9827 57749
rect 10045 57749 10057 57752
rect 10091 57780 10103 57783
rect 11238 57780 11244 57792
rect 10091 57752 11244 57780
rect 10091 57749 10103 57752
rect 10045 57743 10103 57749
rect 11238 57740 11244 57752
rect 11296 57740 11302 57792
rect 1104 57690 10856 57712
rect 1104 57638 4213 57690
rect 4265 57638 4277 57690
rect 4329 57638 4341 57690
rect 4393 57638 4405 57690
rect 4457 57638 4469 57690
rect 4521 57638 7477 57690
rect 7529 57638 7541 57690
rect 7593 57638 7605 57690
rect 7657 57638 7669 57690
rect 7721 57638 7733 57690
rect 7785 57638 10856 57690
rect 1104 57616 10856 57638
rect 1670 57468 1676 57520
rect 1728 57508 1734 57520
rect 11330 57508 11336 57520
rect 1728 57480 11336 57508
rect 1728 57468 1734 57480
rect 11330 57468 11336 57480
rect 11388 57468 11394 57520
rect 1397 57443 1455 57449
rect 1397 57409 1409 57443
rect 1443 57440 1455 57443
rect 9030 57440 9036 57452
rect 1443 57412 9036 57440
rect 1443 57409 1455 57412
rect 1397 57403 1455 57409
rect 9030 57400 9036 57412
rect 9088 57400 9094 57452
rect 9214 57440 9220 57452
rect 9175 57412 9220 57440
rect 9214 57400 9220 57412
rect 9272 57400 9278 57452
rect 9582 57400 9588 57452
rect 9640 57440 9646 57452
rect 9861 57443 9919 57449
rect 9861 57440 9873 57443
rect 9640 57412 9873 57440
rect 9640 57400 9646 57412
rect 9861 57409 9873 57412
rect 9907 57409 9919 57443
rect 9861 57403 9919 57409
rect 1854 57332 1860 57384
rect 1912 57372 1918 57384
rect 5718 57372 5724 57384
rect 1912 57344 5724 57372
rect 1912 57332 1918 57344
rect 5718 57332 5724 57344
rect 5776 57332 5782 57384
rect 1578 57236 1584 57248
rect 1539 57208 1584 57236
rect 1578 57196 1584 57208
rect 1636 57196 1642 57248
rect 5718 57196 5724 57248
rect 5776 57236 5782 57248
rect 9309 57239 9367 57245
rect 9309 57236 9321 57239
rect 5776 57208 9321 57236
rect 5776 57196 5782 57208
rect 9309 57205 9321 57208
rect 9355 57205 9367 57239
rect 9309 57199 9367 57205
rect 10045 57239 10103 57245
rect 10045 57205 10057 57239
rect 10091 57236 10103 57239
rect 11146 57236 11152 57248
rect 10091 57208 11152 57236
rect 10091 57205 10103 57208
rect 10045 57199 10103 57205
rect 11146 57196 11152 57208
rect 11204 57196 11210 57248
rect 1104 57146 10856 57168
rect 1104 57094 2582 57146
rect 2634 57094 2646 57146
rect 2698 57094 2710 57146
rect 2762 57094 2774 57146
rect 2826 57094 2838 57146
rect 2890 57094 5845 57146
rect 5897 57094 5909 57146
rect 5961 57094 5973 57146
rect 6025 57094 6037 57146
rect 6089 57094 6101 57146
rect 6153 57094 9109 57146
rect 9161 57094 9173 57146
rect 9225 57094 9237 57146
rect 9289 57094 9301 57146
rect 9353 57094 9365 57146
rect 9417 57094 10856 57146
rect 1104 57072 10856 57094
rect 1026 56992 1032 57044
rect 1084 57032 1090 57044
rect 5718 57032 5724 57044
rect 1084 57004 5724 57032
rect 1084 56992 1090 57004
rect 5718 56992 5724 57004
rect 5776 56992 5782 57044
rect 3234 56924 3240 56976
rect 3292 56964 3298 56976
rect 3602 56964 3608 56976
rect 3292 56936 3608 56964
rect 3292 56924 3298 56936
rect 3602 56924 3608 56936
rect 3660 56924 3666 56976
rect 5442 56924 5448 56976
rect 5500 56964 5506 56976
rect 9493 56967 9551 56973
rect 9493 56964 9505 56967
rect 5500 56936 9505 56964
rect 5500 56924 5506 56936
rect 9493 56933 9505 56936
rect 9539 56933 9551 56967
rect 11698 56964 11704 56976
rect 11659 56936 11704 56964
rect 9493 56927 9551 56933
rect 11698 56924 11704 56936
rect 11756 56924 11762 56976
rect 9953 56899 10011 56905
rect 9953 56865 9965 56899
rect 9999 56896 10011 56899
rect 10226 56896 10232 56908
rect 9999 56868 10232 56896
rect 9999 56865 10011 56868
rect 9953 56859 10011 56865
rect 10226 56856 10232 56868
rect 10284 56856 10290 56908
rect 1397 56831 1455 56837
rect 1397 56797 1409 56831
rect 1443 56828 1455 56831
rect 3786 56828 3792 56840
rect 1443 56800 3792 56828
rect 1443 56797 1455 56800
rect 1397 56791 1455 56797
rect 3786 56788 3792 56800
rect 3844 56788 3850 56840
rect 6638 56788 6644 56840
rect 6696 56828 6702 56840
rect 11790 56828 11796 56840
rect 6696 56800 11796 56828
rect 6696 56788 6702 56800
rect 11790 56788 11796 56800
rect 11848 56788 11854 56840
rect 10042 56760 10048 56772
rect 10003 56732 10048 56760
rect 10042 56720 10048 56732
rect 10100 56720 10106 56772
rect 1578 56692 1584 56704
rect 1539 56664 1584 56692
rect 1578 56652 1584 56664
rect 1636 56652 1642 56704
rect 9953 56695 10011 56701
rect 9953 56661 9965 56695
rect 9999 56692 10011 56695
rect 10965 56695 11023 56701
rect 10965 56692 10977 56695
rect 9999 56664 10977 56692
rect 9999 56661 10011 56664
rect 9953 56655 10011 56661
rect 10965 56661 10977 56664
rect 11011 56661 11023 56695
rect 10965 56655 11023 56661
rect 1104 56602 10856 56624
rect 1104 56550 4213 56602
rect 4265 56550 4277 56602
rect 4329 56550 4341 56602
rect 4393 56550 4405 56602
rect 4457 56550 4469 56602
rect 4521 56550 7477 56602
rect 7529 56550 7541 56602
rect 7593 56550 7605 56602
rect 7657 56550 7669 56602
rect 7721 56550 7733 56602
rect 7785 56550 10856 56602
rect 1104 56528 10856 56550
rect 1397 56355 1455 56361
rect 1397 56321 1409 56355
rect 1443 56352 1455 56355
rect 2958 56352 2964 56364
rect 1443 56324 2964 56352
rect 1443 56321 1455 56324
rect 1397 56315 1455 56321
rect 2958 56312 2964 56324
rect 3016 56312 3022 56364
rect 9858 56352 9864 56364
rect 9819 56324 9864 56352
rect 9858 56312 9864 56324
rect 9916 56312 9922 56364
rect 1578 56148 1584 56160
rect 1539 56120 1584 56148
rect 1578 56108 1584 56120
rect 1636 56108 1642 56160
rect 7742 56108 7748 56160
rect 7800 56148 7806 56160
rect 8018 56148 8024 56160
rect 7800 56120 8024 56148
rect 7800 56108 7806 56120
rect 8018 56108 8024 56120
rect 8076 56108 8082 56160
rect 10045 56151 10103 56157
rect 10045 56117 10057 56151
rect 10091 56148 10103 56151
rect 10686 56148 10692 56160
rect 10091 56120 10692 56148
rect 10091 56117 10103 56120
rect 10045 56111 10103 56117
rect 10686 56108 10692 56120
rect 10744 56108 10750 56160
rect 1104 56058 10856 56080
rect 1104 56006 2582 56058
rect 2634 56006 2646 56058
rect 2698 56006 2710 56058
rect 2762 56006 2774 56058
rect 2826 56006 2838 56058
rect 2890 56006 5845 56058
rect 5897 56006 5909 56058
rect 5961 56006 5973 56058
rect 6025 56006 6037 56058
rect 6089 56006 6101 56058
rect 6153 56006 9109 56058
rect 9161 56006 9173 56058
rect 9225 56006 9237 56058
rect 9289 56006 9301 56058
rect 9353 56006 9365 56058
rect 9417 56006 10856 56058
rect 10962 56040 10968 56092
rect 11020 56080 11026 56092
rect 11517 56083 11575 56089
rect 11517 56080 11529 56083
rect 11020 56052 11529 56080
rect 11020 56040 11026 56052
rect 11517 56049 11529 56052
rect 11563 56049 11575 56083
rect 11517 56043 11575 56049
rect 1104 55984 10856 56006
rect 11609 55879 11667 55885
rect 11609 55845 11621 55879
rect 11655 55845 11667 55879
rect 11790 55876 11796 55888
rect 11751 55848 11796 55876
rect 11609 55839 11667 55845
rect 1397 55743 1455 55749
rect 1397 55709 1409 55743
rect 1443 55740 1455 55743
rect 5534 55740 5540 55752
rect 1443 55712 5540 55740
rect 1443 55709 1455 55712
rect 1397 55703 1455 55709
rect 5534 55700 5540 55712
rect 5592 55700 5598 55752
rect 9858 55740 9864 55752
rect 9819 55712 9864 55740
rect 9858 55700 9864 55712
rect 9916 55700 9922 55752
rect 11624 55740 11652 55839
rect 11790 55836 11796 55848
rect 11848 55836 11854 55888
rect 11701 55743 11759 55749
rect 11701 55740 11713 55743
rect 11624 55712 11713 55740
rect 11701 55709 11713 55712
rect 11747 55709 11759 55743
rect 11701 55703 11759 55709
rect 1578 55604 1584 55616
rect 1539 55576 1584 55604
rect 1578 55564 1584 55576
rect 1636 55564 1642 55616
rect 9769 55607 9827 55613
rect 9769 55573 9781 55607
rect 9815 55604 9827 55607
rect 10045 55607 10103 55613
rect 10045 55604 10057 55607
rect 9815 55576 10057 55604
rect 9815 55573 9827 55576
rect 9769 55567 9827 55573
rect 10045 55573 10057 55576
rect 10091 55604 10103 55607
rect 11517 55607 11575 55613
rect 11517 55604 11529 55607
rect 10091 55576 11529 55604
rect 10091 55573 10103 55576
rect 10045 55567 10103 55573
rect 11517 55573 11529 55576
rect 11563 55573 11575 55607
rect 11517 55567 11575 55573
rect 1104 55514 10856 55536
rect 1104 55462 4213 55514
rect 4265 55462 4277 55514
rect 4329 55462 4341 55514
rect 4393 55462 4405 55514
rect 4457 55462 4469 55514
rect 4521 55462 7477 55514
rect 7529 55462 7541 55514
rect 7593 55462 7605 55514
rect 7657 55462 7669 55514
rect 7721 55462 7733 55514
rect 7785 55462 10856 55514
rect 1104 55440 10856 55462
rect 1397 55267 1455 55273
rect 1397 55233 1409 55267
rect 1443 55264 1455 55267
rect 2222 55264 2228 55276
rect 1443 55236 2228 55264
rect 1443 55233 1455 55236
rect 1397 55227 1455 55233
rect 2222 55224 2228 55236
rect 2280 55224 2286 55276
rect 9858 55264 9864 55276
rect 9819 55236 9864 55264
rect 9858 55224 9864 55236
rect 9916 55224 9922 55276
rect 10870 55156 10876 55208
rect 10928 55196 10934 55208
rect 11149 55199 11207 55205
rect 11149 55196 11161 55199
rect 10928 55168 11161 55196
rect 10928 55156 10934 55168
rect 11149 55165 11161 55168
rect 11195 55165 11207 55199
rect 11149 55159 11207 55165
rect 1578 55060 1584 55072
rect 1539 55032 1584 55060
rect 1578 55020 1584 55032
rect 1636 55020 1642 55072
rect 10045 55063 10103 55069
rect 10045 55029 10057 55063
rect 10091 55060 10103 55063
rect 11149 55063 11207 55069
rect 11149 55060 11161 55063
rect 10091 55032 11161 55060
rect 10091 55029 10103 55032
rect 10045 55023 10103 55029
rect 11149 55029 11161 55032
rect 11195 55029 11207 55063
rect 11149 55023 11207 55029
rect 1104 54970 10856 54992
rect 1104 54918 2582 54970
rect 2634 54918 2646 54970
rect 2698 54918 2710 54970
rect 2762 54918 2774 54970
rect 2826 54918 2838 54970
rect 2890 54918 5845 54970
rect 5897 54918 5909 54970
rect 5961 54918 5973 54970
rect 6025 54918 6037 54970
rect 6089 54918 6101 54970
rect 6153 54918 9109 54970
rect 9161 54918 9173 54970
rect 9225 54918 9237 54970
rect 9289 54918 9301 54970
rect 9353 54918 9365 54970
rect 9417 54918 10856 54970
rect 1104 54896 10856 54918
rect 1670 54856 1676 54868
rect 1631 54828 1676 54856
rect 1670 54816 1676 54828
rect 1728 54816 1734 54868
rect 1946 54680 1952 54732
rect 2004 54720 2010 54732
rect 2130 54720 2136 54732
rect 2004 54692 2136 54720
rect 2004 54680 2010 54692
rect 2130 54680 2136 54692
rect 2188 54680 2194 54732
rect 2225 54587 2283 54593
rect 2225 54553 2237 54587
rect 2271 54584 2283 54587
rect 2314 54584 2320 54596
rect 2271 54556 2320 54584
rect 2271 54553 2283 54556
rect 2225 54547 2283 54553
rect 2314 54544 2320 54556
rect 2372 54584 2378 54596
rect 2498 54584 2504 54596
rect 2372 54556 2504 54584
rect 2372 54544 2378 54556
rect 2498 54544 2504 54556
rect 2556 54544 2562 54596
rect 9950 54584 9956 54596
rect 9911 54556 9956 54584
rect 9950 54544 9956 54556
rect 10008 54544 10014 54596
rect 10137 54587 10195 54593
rect 10137 54553 10149 54587
rect 10183 54584 10195 54587
rect 11609 54587 11667 54593
rect 11609 54584 11621 54587
rect 10183 54556 11621 54584
rect 10183 54553 10195 54556
rect 10137 54547 10195 54553
rect 11609 54553 11621 54556
rect 11655 54553 11667 54587
rect 11609 54547 11667 54553
rect 1670 54476 1676 54528
rect 1728 54516 1734 54528
rect 2133 54519 2191 54525
rect 2133 54516 2145 54519
rect 1728 54488 2145 54516
rect 1728 54476 1734 54488
rect 2133 54485 2145 54488
rect 2179 54485 2191 54519
rect 2133 54479 2191 54485
rect 1104 54426 10856 54448
rect 1104 54374 4213 54426
rect 4265 54374 4277 54426
rect 4329 54374 4341 54426
rect 4393 54374 4405 54426
rect 4457 54374 4469 54426
rect 4521 54374 7477 54426
rect 7529 54374 7541 54426
rect 7593 54374 7605 54426
rect 7657 54374 7669 54426
rect 7721 54374 7733 54426
rect 7785 54374 10856 54426
rect 1104 54352 10856 54374
rect 2406 54312 2412 54324
rect 2367 54284 2412 54312
rect 2406 54272 2412 54284
rect 2464 54272 2470 54324
rect 1486 54136 1492 54188
rect 1544 54176 1550 54188
rect 1946 54176 1952 54188
rect 1544 54148 1952 54176
rect 1544 54136 1550 54148
rect 1946 54136 1952 54148
rect 2004 54176 2010 54188
rect 2225 54179 2283 54185
rect 2225 54176 2237 54179
rect 2004 54148 2237 54176
rect 2004 54136 2010 54148
rect 2225 54145 2237 54148
rect 2271 54145 2283 54179
rect 2225 54139 2283 54145
rect 9125 54179 9183 54185
rect 9125 54145 9137 54179
rect 9171 54176 9183 54179
rect 9490 54176 9496 54188
rect 9171 54148 9496 54176
rect 9171 54145 9183 54148
rect 9125 54139 9183 54145
rect 9490 54136 9496 54148
rect 9548 54136 9554 54188
rect 9861 54179 9919 54185
rect 9861 54145 9873 54179
rect 9907 54176 9919 54179
rect 9950 54176 9956 54188
rect 9907 54148 9956 54176
rect 9907 54145 9919 54148
rect 9861 54139 9919 54145
rect 9950 54136 9956 54148
rect 10008 54136 10014 54188
rect 2406 54068 2412 54120
rect 2464 54108 2470 54120
rect 2501 54111 2559 54117
rect 2501 54108 2513 54111
rect 2464 54080 2513 54108
rect 2464 54068 2470 54080
rect 2501 54077 2513 54080
rect 2547 54077 2559 54111
rect 2501 54071 2559 54077
rect 9769 54043 9827 54049
rect 9769 54009 9781 54043
rect 9815 54040 9827 54043
rect 10045 54043 10103 54049
rect 10045 54040 10057 54043
rect 9815 54012 10057 54040
rect 9815 54009 9827 54012
rect 9769 54003 9827 54009
rect 10045 54009 10057 54012
rect 10091 54040 10103 54043
rect 11793 54043 11851 54049
rect 11793 54040 11805 54043
rect 10091 54012 11805 54040
rect 10091 54009 10103 54012
rect 10045 54003 10103 54009
rect 11793 54009 11805 54012
rect 11839 54009 11851 54043
rect 11793 54003 11851 54009
rect 382 53932 388 53984
rect 440 53972 446 53984
rect 1949 53975 2007 53981
rect 1949 53972 1961 53975
rect 440 53944 1961 53972
rect 440 53932 446 53944
rect 1949 53941 1961 53944
rect 1995 53941 2007 53975
rect 1949 53935 2007 53941
rect 3050 53932 3056 53984
rect 3108 53972 3114 53984
rect 6546 53972 6552 53984
rect 3108 53944 6552 53972
rect 3108 53932 3114 53944
rect 6546 53932 6552 53944
rect 6604 53932 6610 53984
rect 8662 53932 8668 53984
rect 8720 53972 8726 53984
rect 9309 53975 9367 53981
rect 9309 53972 9321 53975
rect 8720 53944 9321 53972
rect 8720 53932 8726 53944
rect 9309 53941 9321 53944
rect 9355 53941 9367 53975
rect 9309 53935 9367 53941
rect 10226 53932 10232 53984
rect 10284 53972 10290 53984
rect 10410 53972 10416 53984
rect 10284 53944 10416 53972
rect 10284 53932 10290 53944
rect 10410 53932 10416 53944
rect 10468 53932 10474 53984
rect 1104 53882 10856 53904
rect 1104 53830 2582 53882
rect 2634 53830 2646 53882
rect 2698 53830 2710 53882
rect 2762 53830 2774 53882
rect 2826 53830 2838 53882
rect 2890 53830 5845 53882
rect 5897 53830 5909 53882
rect 5961 53830 5973 53882
rect 6025 53830 6037 53882
rect 6089 53830 6101 53882
rect 6153 53830 9109 53882
rect 9161 53830 9173 53882
rect 9225 53830 9237 53882
rect 9289 53830 9301 53882
rect 9353 53830 9365 53882
rect 9417 53830 10856 53882
rect 1104 53808 10856 53830
rect 1578 53768 1584 53780
rect 1539 53740 1584 53768
rect 1578 53728 1584 53740
rect 1636 53728 1642 53780
rect 10134 53592 10140 53644
rect 10192 53592 10198 53644
rect 1397 53567 1455 53573
rect 1397 53533 1409 53567
rect 1443 53564 1455 53567
rect 1486 53564 1492 53576
rect 1443 53536 1492 53564
rect 1443 53533 1455 53536
rect 1397 53527 1455 53533
rect 1486 53524 1492 53536
rect 1544 53524 1550 53576
rect 9125 53567 9183 53573
rect 9125 53533 9137 53567
rect 9171 53564 9183 53567
rect 9582 53564 9588 53576
rect 9171 53536 9588 53564
rect 9171 53533 9183 53536
rect 9125 53527 9183 53533
rect 9582 53524 9588 53536
rect 9640 53524 9646 53576
rect 9858 53564 9864 53576
rect 9819 53536 9864 53564
rect 9858 53524 9864 53536
rect 9916 53524 9922 53576
rect 10152 53440 10180 53592
rect 8570 53388 8576 53440
rect 8628 53428 8634 53440
rect 9309 53431 9367 53437
rect 9309 53428 9321 53431
rect 8628 53400 9321 53428
rect 8628 53388 8634 53400
rect 9309 53397 9321 53400
rect 9355 53397 9367 53431
rect 9309 53391 9367 53397
rect 9769 53431 9827 53437
rect 9769 53397 9781 53431
rect 9815 53428 9827 53431
rect 10042 53428 10048 53440
rect 9815 53400 10048 53428
rect 9815 53397 9827 53400
rect 9769 53391 9827 53397
rect 10042 53388 10048 53400
rect 10100 53388 10106 53440
rect 10134 53388 10140 53440
rect 10192 53388 10198 53440
rect 1104 53338 10856 53360
rect 1104 53286 4213 53338
rect 4265 53286 4277 53338
rect 4329 53286 4341 53338
rect 4393 53286 4405 53338
rect 4457 53286 4469 53338
rect 4521 53286 7477 53338
rect 7529 53286 7541 53338
rect 7593 53286 7605 53338
rect 7657 53286 7669 53338
rect 7721 53286 7733 53338
rect 7785 53286 10856 53338
rect 1104 53264 10856 53286
rect 1578 53224 1584 53236
rect 1539 53196 1584 53224
rect 1578 53184 1584 53196
rect 1636 53184 1642 53236
rect 9953 53227 10011 53233
rect 9953 53193 9965 53227
rect 9999 53224 10011 53227
rect 11514 53224 11520 53236
rect 9999 53196 11520 53224
rect 9999 53193 10011 53196
rect 9953 53187 10011 53193
rect 11514 53184 11520 53196
rect 11572 53184 11578 53236
rect 10962 53116 10968 53168
rect 11020 53156 11026 53168
rect 11885 53159 11943 53165
rect 11885 53156 11897 53159
rect 11020 53128 11897 53156
rect 11020 53116 11026 53128
rect 11885 53125 11897 53128
rect 11931 53125 11943 53159
rect 11885 53119 11943 53125
rect 1397 53091 1455 53097
rect 1397 53057 1409 53091
rect 1443 53088 1455 53091
rect 2498 53088 2504 53100
rect 1443 53060 2504 53088
rect 1443 53057 1455 53060
rect 1397 53051 1455 53057
rect 2498 53048 2504 53060
rect 2556 53048 2562 53100
rect 9766 53088 9772 53100
rect 9727 53060 9772 53088
rect 9766 53048 9772 53060
rect 9824 53048 9830 53100
rect 11425 53091 11483 53097
rect 11425 53057 11437 53091
rect 11471 53088 11483 53091
rect 11514 53088 11520 53100
rect 11471 53060 11520 53088
rect 11471 53057 11483 53060
rect 11425 53051 11483 53057
rect 11514 53048 11520 53060
rect 11572 53048 11578 53100
rect 10045 53023 10103 53029
rect 10045 52989 10057 53023
rect 10091 53020 10103 53023
rect 10226 53020 10232 53032
rect 10091 52992 10232 53020
rect 10091 52989 10103 52992
rect 10045 52983 10103 52989
rect 10226 52980 10232 52992
rect 10284 52980 10290 53032
rect 11882 53020 11888 53032
rect 11843 52992 11888 53020
rect 11882 52980 11888 52992
rect 11940 52980 11946 53032
rect 9493 52887 9551 52893
rect 9493 52853 9505 52887
rect 9539 52884 9551 52887
rect 11238 52884 11244 52896
rect 9539 52856 11244 52884
rect 9539 52853 9551 52856
rect 9493 52847 9551 52853
rect 11238 52844 11244 52856
rect 11296 52844 11302 52896
rect 1104 52794 10856 52816
rect 1104 52742 2582 52794
rect 2634 52742 2646 52794
rect 2698 52742 2710 52794
rect 2762 52742 2774 52794
rect 2826 52742 2838 52794
rect 2890 52742 5845 52794
rect 5897 52742 5909 52794
rect 5961 52742 5973 52794
rect 6025 52742 6037 52794
rect 6089 52742 6101 52794
rect 6153 52742 9109 52794
rect 9161 52742 9173 52794
rect 9225 52742 9237 52794
rect 9289 52742 9301 52794
rect 9353 52742 9365 52794
rect 9417 52742 10856 52794
rect 1104 52720 10856 52742
rect 1673 52683 1731 52689
rect 1673 52649 1685 52683
rect 1719 52680 1731 52683
rect 11422 52680 11428 52692
rect 1719 52652 11428 52680
rect 1719 52649 1731 52652
rect 1673 52643 1731 52649
rect 11422 52640 11428 52652
rect 11480 52640 11486 52692
rect 2774 52572 2780 52624
rect 2832 52612 2838 52624
rect 2832 52584 2877 52612
rect 2832 52572 2838 52584
rect 4706 52572 4712 52624
rect 4764 52612 4770 52624
rect 9309 52615 9367 52621
rect 9309 52612 9321 52615
rect 4764 52584 9321 52612
rect 4764 52572 4770 52584
rect 9309 52581 9321 52584
rect 9355 52581 9367 52615
rect 9309 52575 9367 52581
rect 1670 52436 1676 52488
rect 1728 52476 1734 52488
rect 1949 52479 2007 52485
rect 1949 52476 1961 52479
rect 1728 52448 1961 52476
rect 1728 52436 1734 52448
rect 1949 52445 1961 52448
rect 1995 52445 2007 52479
rect 1949 52439 2007 52445
rect 2225 52479 2283 52485
rect 2225 52445 2237 52479
rect 2271 52476 2283 52479
rect 2406 52476 2412 52488
rect 2271 52448 2412 52476
rect 2271 52445 2283 52448
rect 2225 52439 2283 52445
rect 2406 52436 2412 52448
rect 2464 52436 2470 52488
rect 2958 52476 2964 52488
rect 2919 52448 2964 52476
rect 2958 52436 2964 52448
rect 3016 52436 3022 52488
rect 9122 52476 9128 52488
rect 9083 52448 9128 52476
rect 9122 52436 9128 52448
rect 9180 52436 9186 52488
rect 9861 52479 9919 52485
rect 9861 52445 9873 52479
rect 9907 52476 9919 52479
rect 10965 52479 11023 52485
rect 10965 52476 10977 52479
rect 9907 52448 10977 52476
rect 9907 52445 9919 52448
rect 9861 52439 9919 52445
rect 10965 52445 10977 52448
rect 11011 52445 11023 52479
rect 10965 52439 11023 52445
rect 2130 52408 2136 52420
rect 2091 52380 2136 52408
rect 2130 52368 2136 52380
rect 2188 52368 2194 52420
rect 9769 52343 9827 52349
rect 9769 52309 9781 52343
rect 9815 52340 9827 52343
rect 10045 52343 10103 52349
rect 10045 52340 10057 52343
rect 9815 52312 10057 52340
rect 9815 52309 9827 52312
rect 9769 52303 9827 52309
rect 10045 52309 10057 52312
rect 10091 52340 10103 52343
rect 10686 52340 10692 52352
rect 10091 52312 10692 52340
rect 10091 52309 10103 52312
rect 10045 52303 10103 52309
rect 10686 52300 10692 52312
rect 10744 52300 10750 52352
rect 1104 52250 10856 52272
rect 1104 52198 4213 52250
rect 4265 52198 4277 52250
rect 4329 52198 4341 52250
rect 4393 52198 4405 52250
rect 4457 52198 4469 52250
rect 4521 52198 7477 52250
rect 7529 52198 7541 52250
rect 7593 52198 7605 52250
rect 7657 52198 7669 52250
rect 7721 52198 7733 52250
rect 7785 52198 10856 52250
rect 1104 52176 10856 52198
rect 1854 52096 1860 52148
rect 1912 52136 1918 52148
rect 1949 52139 2007 52145
rect 1949 52136 1961 52139
rect 1912 52108 1961 52136
rect 1912 52096 1918 52108
rect 1949 52105 1961 52108
rect 1995 52105 2007 52139
rect 1949 52099 2007 52105
rect 1854 52000 1860 52012
rect 1815 51972 1860 52000
rect 1854 51960 1860 51972
rect 1912 51960 1918 52012
rect 9125 52003 9183 52009
rect 9125 51969 9137 52003
rect 9171 52000 9183 52003
rect 9490 52000 9496 52012
rect 9171 51972 9496 52000
rect 9171 51969 9183 51972
rect 9125 51963 9183 51969
rect 9490 51960 9496 51972
rect 9548 51960 9554 52012
rect 9858 52000 9864 52012
rect 9819 51972 9864 52000
rect 9858 51960 9864 51972
rect 9916 51960 9922 52012
rect 6822 51756 6828 51808
rect 6880 51796 6886 51808
rect 9309 51799 9367 51805
rect 9309 51796 9321 51799
rect 6880 51768 9321 51796
rect 6880 51756 6886 51768
rect 9309 51765 9321 51768
rect 9355 51765 9367 51799
rect 10042 51796 10048 51808
rect 10003 51768 10048 51796
rect 9309 51759 9367 51765
rect 10042 51756 10048 51768
rect 10100 51756 10106 51808
rect 1104 51706 10856 51728
rect 1104 51654 2582 51706
rect 2634 51654 2646 51706
rect 2698 51654 2710 51706
rect 2762 51654 2774 51706
rect 2826 51654 2838 51706
rect 2890 51654 5845 51706
rect 5897 51654 5909 51706
rect 5961 51654 5973 51706
rect 6025 51654 6037 51706
rect 6089 51654 6101 51706
rect 6153 51654 9109 51706
rect 9161 51654 9173 51706
rect 9225 51654 9237 51706
rect 9289 51654 9301 51706
rect 9353 51654 9365 51706
rect 9417 51654 10856 51706
rect 1104 51632 10856 51654
rect 1581 51595 1639 51601
rect 1581 51561 1593 51595
rect 1627 51592 1639 51595
rect 6638 51592 6644 51604
rect 1627 51564 6644 51592
rect 1627 51561 1639 51564
rect 1581 51555 1639 51561
rect 6638 51552 6644 51564
rect 6696 51552 6702 51604
rect 8846 51552 8852 51604
rect 8904 51592 8910 51604
rect 8941 51595 8999 51601
rect 8941 51592 8953 51595
rect 8904 51564 8953 51592
rect 8904 51552 8910 51564
rect 8941 51561 8953 51564
rect 8987 51561 8999 51595
rect 10870 51592 10876 51604
rect 10831 51564 10876 51592
rect 8941 51555 8999 51561
rect 10870 51552 10876 51564
rect 10928 51552 10934 51604
rect 2590 51484 2596 51536
rect 2648 51524 2654 51536
rect 9582 51524 9588 51536
rect 2648 51496 9588 51524
rect 2648 51484 2654 51496
rect 9582 51484 9588 51496
rect 9640 51484 9646 51536
rect 11241 51527 11299 51533
rect 11241 51493 11253 51527
rect 11287 51493 11299 51527
rect 11241 51487 11299 51493
rect 2406 51416 2412 51468
rect 2464 51456 2470 51468
rect 9493 51459 9551 51465
rect 9493 51456 9505 51459
rect 2464 51428 9505 51456
rect 2464 51416 2470 51428
rect 9493 51425 9505 51428
rect 9539 51456 9551 51459
rect 10226 51456 10232 51468
rect 9539 51428 10232 51456
rect 9539 51425 9551 51428
rect 9493 51419 9551 51425
rect 10226 51416 10232 51428
rect 10284 51416 10290 51468
rect 10870 51416 10876 51468
rect 10928 51456 10934 51468
rect 11149 51459 11207 51465
rect 11149 51456 11161 51459
rect 10928 51428 11161 51456
rect 10928 51416 10934 51428
rect 11149 51425 11161 51428
rect 11195 51425 11207 51459
rect 11149 51419 11207 51425
rect 1394 51388 1400 51400
rect 1355 51360 1400 51388
rect 1394 51348 1400 51360
rect 1452 51348 1458 51400
rect 10962 51388 10968 51400
rect 10923 51360 10968 51388
rect 10962 51348 10968 51360
rect 11020 51348 11026 51400
rect 11054 51348 11060 51400
rect 11112 51388 11118 51400
rect 11112 51360 11157 51388
rect 11112 51348 11118 51360
rect 9309 51323 9367 51329
rect 9309 51289 9321 51323
rect 9355 51320 9367 51323
rect 9490 51320 9496 51332
rect 9355 51292 9496 51320
rect 9355 51289 9367 51292
rect 9309 51283 9367 51289
rect 9490 51280 9496 51292
rect 9548 51280 9554 51332
rect 6638 51212 6644 51264
rect 6696 51252 6702 51264
rect 8202 51252 8208 51264
rect 6696 51224 8208 51252
rect 6696 51212 6702 51224
rect 8202 51212 8208 51224
rect 8260 51212 8266 51264
rect 9401 51255 9459 51261
rect 9401 51221 9413 51255
rect 9447 51252 9459 51255
rect 9674 51252 9680 51264
rect 9447 51224 9680 51252
rect 9447 51221 9459 51224
rect 9401 51215 9459 51221
rect 9674 51212 9680 51224
rect 9732 51212 9738 51264
rect 10778 51212 10784 51264
rect 10836 51252 10842 51264
rect 10836 51224 10916 51252
rect 10836 51212 10842 51224
rect 1104 51162 10856 51184
rect 1104 51110 4213 51162
rect 4265 51110 4277 51162
rect 4329 51110 4341 51162
rect 4393 51110 4405 51162
rect 4457 51110 4469 51162
rect 4521 51110 7477 51162
rect 7529 51110 7541 51162
rect 7593 51110 7605 51162
rect 7657 51110 7669 51162
rect 7721 51110 7733 51162
rect 7785 51110 10856 51162
rect 1104 51088 10856 51110
rect 10888 51116 10916 51224
rect 10962 51144 10968 51196
rect 11020 51184 11026 51196
rect 11256 51184 11284 51487
rect 11330 51416 11336 51468
rect 11388 51456 11394 51468
rect 11425 51459 11483 51465
rect 11425 51456 11437 51459
rect 11388 51428 11437 51456
rect 11388 51416 11394 51428
rect 11425 51425 11437 51428
rect 11471 51425 11483 51459
rect 11425 51419 11483 51425
rect 11790 51388 11796 51400
rect 11751 51360 11796 51388
rect 11790 51348 11796 51360
rect 11848 51348 11854 51400
rect 11517 51323 11575 51329
rect 11517 51289 11529 51323
rect 11563 51289 11575 51323
rect 11517 51283 11575 51289
rect 11609 51323 11667 51329
rect 11609 51289 11621 51323
rect 11655 51289 11667 51323
rect 11609 51283 11667 51289
rect 11532 51193 11560 51283
rect 11624 51193 11652 51283
rect 11020 51156 11284 51184
rect 11517 51187 11575 51193
rect 11020 51144 11026 51156
rect 11517 51153 11529 51187
rect 11563 51153 11575 51187
rect 11517 51147 11575 51153
rect 11609 51187 11667 51193
rect 11609 51153 11621 51187
rect 11655 51153 11667 51187
rect 11609 51147 11667 51153
rect 11330 51116 11336 51128
rect 10888 51088 11336 51116
rect 11330 51076 11336 51088
rect 11388 51076 11394 51128
rect 934 51008 940 51060
rect 992 51048 998 51060
rect 1949 51051 2007 51057
rect 1949 51048 1961 51051
rect 992 51020 1961 51048
rect 992 51008 998 51020
rect 1949 51017 1961 51020
rect 1995 51017 2007 51051
rect 2498 51048 2504 51060
rect 2459 51020 2504 51048
rect 1949 51011 2007 51017
rect 2498 51008 2504 51020
rect 2556 51008 2562 51060
rect 3142 51008 3148 51060
rect 3200 51008 3206 51060
rect 7006 51008 7012 51060
rect 7064 51048 7070 51060
rect 7064 51020 7236 51048
rect 7064 51008 7070 51020
rect 1854 50912 1860 50924
rect 1815 50884 1860 50912
rect 1854 50872 1860 50884
rect 1912 50872 1918 50924
rect 2685 50915 2743 50921
rect 2685 50881 2697 50915
rect 2731 50881 2743 50915
rect 2685 50875 2743 50881
rect 474 50804 480 50856
rect 532 50844 538 50856
rect 2700 50844 2728 50875
rect 532 50816 2728 50844
rect 3160 50844 3188 51008
rect 7208 50856 7236 51020
rect 7282 51008 7288 51060
rect 7340 51008 7346 51060
rect 7374 51008 7380 51060
rect 7432 51008 7438 51060
rect 8294 51008 8300 51060
rect 8352 51048 8358 51060
rect 8757 51051 8815 51057
rect 8757 51048 8769 51051
rect 8352 51020 8769 51048
rect 8352 51008 8358 51020
rect 8757 51017 8769 51020
rect 8803 51017 8815 51051
rect 8757 51011 8815 51017
rect 10962 51008 10968 51060
rect 11020 51048 11026 51060
rect 11057 51051 11115 51057
rect 11057 51048 11069 51051
rect 11020 51020 11069 51048
rect 11020 51008 11026 51020
rect 11057 51017 11069 51020
rect 11103 51017 11115 51051
rect 11057 51011 11115 51017
rect 11425 51051 11483 51057
rect 11425 51017 11437 51051
rect 11471 51017 11483 51051
rect 11425 51011 11483 51017
rect 7300 50856 7328 51008
rect 7392 50856 7420 51008
rect 9766 50980 9772 50992
rect 8312 50952 9772 50980
rect 8312 50924 8340 50952
rect 9766 50940 9772 50952
rect 9824 50940 9830 50992
rect 10686 50940 10692 50992
rect 10744 50980 10750 50992
rect 11333 50983 11391 50989
rect 11333 50980 11345 50983
rect 10744 50952 11345 50980
rect 10744 50940 10750 50952
rect 11333 50949 11345 50952
rect 11379 50949 11391 50983
rect 11333 50943 11391 50949
rect 8294 50872 8300 50924
rect 8352 50872 8358 50924
rect 8938 50872 8944 50924
rect 8996 50912 9002 50924
rect 9125 50915 9183 50921
rect 9125 50912 9137 50915
rect 8996 50884 9137 50912
rect 8996 50872 9002 50884
rect 9125 50881 9137 50884
rect 9171 50881 9183 50915
rect 9125 50875 9183 50881
rect 10137 50915 10195 50921
rect 10137 50881 10149 50915
rect 10183 50912 10195 50915
rect 10965 50915 11023 50921
rect 10965 50912 10977 50915
rect 10183 50884 10977 50912
rect 10183 50881 10195 50884
rect 10137 50875 10195 50881
rect 10965 50881 10977 50884
rect 11011 50881 11023 50915
rect 11440 50912 11468 51011
rect 11698 50940 11704 50992
rect 11756 50980 11762 50992
rect 11756 50952 11801 50980
rect 11756 50940 11762 50952
rect 11440 50884 11836 50912
rect 10965 50875 11023 50881
rect 3602 50844 3608 50856
rect 3160 50816 3608 50844
rect 532 50804 538 50816
rect 3602 50804 3608 50816
rect 3660 50804 3666 50856
rect 7190 50804 7196 50856
rect 7248 50804 7254 50856
rect 7282 50804 7288 50856
rect 7340 50804 7346 50856
rect 7374 50804 7380 50856
rect 7432 50804 7438 50856
rect 8846 50804 8852 50856
rect 8904 50844 8910 50856
rect 9217 50847 9275 50853
rect 9217 50844 9229 50847
rect 8904 50816 9229 50844
rect 8904 50804 8910 50816
rect 9217 50813 9229 50816
rect 9263 50813 9275 50847
rect 9217 50807 9275 50813
rect 9401 50847 9459 50853
rect 9401 50813 9413 50847
rect 9447 50844 9459 50847
rect 10226 50844 10232 50856
rect 9447 50816 10232 50844
rect 9447 50813 9459 50816
rect 9401 50807 9459 50813
rect 9508 50720 9536 50816
rect 10226 50804 10232 50816
rect 10284 50804 10290 50856
rect 11146 50804 11152 50856
rect 11204 50804 11210 50856
rect 11164 50776 11192 50804
rect 10796 50748 11192 50776
rect 11609 50779 11667 50785
rect 10796 50720 10824 50748
rect 11609 50745 11621 50779
rect 11655 50776 11667 50779
rect 11655 50748 11744 50776
rect 11655 50745 11667 50748
rect 11609 50739 11667 50745
rect 9490 50668 9496 50720
rect 9548 50668 9554 50720
rect 9582 50668 9588 50720
rect 9640 50708 9646 50720
rect 9953 50711 10011 50717
rect 9953 50708 9965 50711
rect 9640 50680 9965 50708
rect 9640 50668 9646 50680
rect 9953 50677 9965 50680
rect 9999 50677 10011 50711
rect 9953 50671 10011 50677
rect 10778 50668 10784 50720
rect 10836 50668 10842 50720
rect 10873 50711 10931 50717
rect 10873 50677 10885 50711
rect 10919 50677 10931 50711
rect 10873 50671 10931 50677
rect 11149 50711 11207 50717
rect 11149 50677 11161 50711
rect 11195 50708 11207 50711
rect 11422 50708 11428 50720
rect 11195 50680 11428 50708
rect 11195 50677 11207 50680
rect 11149 50671 11207 50677
rect 10888 50640 10916 50671
rect 11422 50668 11428 50680
rect 11480 50668 11486 50720
rect 11241 50643 11299 50649
rect 11241 50640 11253 50643
rect 1104 50618 10856 50640
rect 1104 50566 2582 50618
rect 2634 50566 2646 50618
rect 2698 50566 2710 50618
rect 2762 50566 2774 50618
rect 2826 50566 2838 50618
rect 2890 50566 5845 50618
rect 5897 50566 5909 50618
rect 5961 50566 5973 50618
rect 6025 50566 6037 50618
rect 6089 50566 6101 50618
rect 6153 50566 9109 50618
rect 9161 50566 9173 50618
rect 9225 50566 9237 50618
rect 9289 50566 9301 50618
rect 9353 50566 9365 50618
rect 9417 50566 10856 50618
rect 10888 50612 11253 50640
rect 11241 50609 11253 50612
rect 11287 50609 11299 50643
rect 11241 50603 11299 50609
rect 11330 50600 11336 50652
rect 11388 50640 11394 50652
rect 11609 50643 11667 50649
rect 11609 50640 11621 50643
rect 11388 50612 11621 50640
rect 11388 50600 11394 50612
rect 11609 50609 11621 50612
rect 11655 50609 11667 50643
rect 11716 50640 11744 50748
rect 11808 50717 11836 50884
rect 11793 50711 11851 50717
rect 11793 50677 11805 50711
rect 11839 50677 11851 50711
rect 11793 50671 11851 50677
rect 11716 50612 11836 50640
rect 11609 50603 11667 50609
rect 1104 50544 10856 50566
rect 1210 50464 1216 50516
rect 1268 50504 1274 50516
rect 1949 50507 2007 50513
rect 1949 50504 1961 50507
rect 1268 50476 1961 50504
rect 1268 50464 1274 50476
rect 1949 50473 1961 50476
rect 1995 50473 2007 50507
rect 1949 50467 2007 50473
rect 9030 50464 9036 50516
rect 9088 50504 9094 50516
rect 9125 50507 9183 50513
rect 9125 50504 9137 50507
rect 9088 50476 9137 50504
rect 9088 50464 9094 50476
rect 9125 50473 9137 50476
rect 9171 50473 9183 50507
rect 9125 50467 9183 50473
rect 11517 50507 11575 50513
rect 11517 50473 11529 50507
rect 11563 50504 11575 50507
rect 11808 50504 11836 50612
rect 11563 50476 11836 50504
rect 11563 50473 11575 50476
rect 11517 50467 11575 50473
rect 9950 50396 9956 50448
rect 10008 50436 10014 50448
rect 11882 50436 11888 50448
rect 10008 50408 11888 50436
rect 10008 50396 10014 50408
rect 11882 50396 11888 50408
rect 11940 50396 11946 50448
rect 9490 50328 9496 50380
rect 9548 50368 9554 50380
rect 9769 50371 9827 50377
rect 9769 50368 9781 50371
rect 9548 50340 9781 50368
rect 9548 50328 9554 50340
rect 9769 50337 9781 50340
rect 9815 50368 9827 50371
rect 9858 50368 9864 50380
rect 9815 50340 9864 50368
rect 9815 50337 9827 50340
rect 9769 50331 9827 50337
rect 9858 50328 9864 50340
rect 9916 50328 9922 50380
rect 11701 50371 11759 50377
rect 11701 50337 11713 50371
rect 11747 50368 11759 50371
rect 11790 50368 11796 50380
rect 11747 50340 11796 50368
rect 11747 50337 11759 50340
rect 11701 50331 11759 50337
rect 11790 50328 11796 50340
rect 11848 50328 11854 50380
rect 8110 50300 8116 50312
rect 8071 50272 8116 50300
rect 8110 50260 8116 50272
rect 8168 50260 8174 50312
rect 1854 50232 1860 50244
rect 1815 50204 1860 50232
rect 1854 50192 1860 50204
rect 1912 50192 1918 50244
rect 3050 50192 3056 50244
rect 3108 50232 3114 50244
rect 5258 50232 5264 50244
rect 3108 50204 5264 50232
rect 3108 50192 3114 50204
rect 5258 50192 5264 50204
rect 5316 50192 5322 50244
rect 8297 50167 8355 50173
rect 8297 50133 8309 50167
rect 8343 50164 8355 50167
rect 8386 50164 8392 50176
rect 8343 50136 8392 50164
rect 8343 50133 8355 50136
rect 8297 50127 8355 50133
rect 8386 50124 8392 50136
rect 8444 50124 8450 50176
rect 8754 50124 8760 50176
rect 8812 50164 8818 50176
rect 9030 50164 9036 50176
rect 8812 50136 9036 50164
rect 8812 50124 8818 50136
rect 9030 50124 9036 50136
rect 9088 50124 9094 50176
rect 9490 50164 9496 50176
rect 9451 50136 9496 50164
rect 9490 50124 9496 50136
rect 9548 50124 9554 50176
rect 9585 50167 9643 50173
rect 9585 50133 9597 50167
rect 9631 50164 9643 50167
rect 9674 50164 9680 50176
rect 9631 50136 9680 50164
rect 9631 50133 9643 50136
rect 9585 50127 9643 50133
rect 9674 50124 9680 50136
rect 9732 50124 9738 50176
rect 1104 50074 10856 50096
rect 1104 50022 4213 50074
rect 4265 50022 4277 50074
rect 4329 50022 4341 50074
rect 4393 50022 4405 50074
rect 4457 50022 4469 50074
rect 4521 50022 7477 50074
rect 7529 50022 7541 50074
rect 7593 50022 7605 50074
rect 7657 50022 7669 50074
rect 7721 50022 7733 50074
rect 7785 50022 10856 50074
rect 1104 50000 10856 50022
rect 5258 49920 5264 49972
rect 5316 49960 5322 49972
rect 8849 49963 8907 49969
rect 8849 49960 8861 49963
rect 5316 49932 8861 49960
rect 5316 49920 5322 49932
rect 8849 49929 8861 49932
rect 8895 49929 8907 49963
rect 9950 49960 9956 49972
rect 9911 49932 9956 49960
rect 8849 49923 8907 49929
rect 9950 49920 9956 49932
rect 10008 49920 10014 49972
rect 6546 49852 6552 49904
rect 6604 49892 6610 49904
rect 6822 49892 6828 49904
rect 6604 49864 6828 49892
rect 6604 49852 6610 49864
rect 6822 49852 6828 49864
rect 6880 49852 6886 49904
rect 8662 49824 8668 49836
rect 8623 49796 8668 49824
rect 8662 49784 8668 49796
rect 8720 49784 8726 49836
rect 9858 49784 9864 49836
rect 9916 49824 9922 49836
rect 10045 49827 10103 49833
rect 10045 49824 10057 49827
rect 9916 49796 10057 49824
rect 9916 49784 9922 49796
rect 10045 49793 10057 49796
rect 10091 49793 10103 49827
rect 10045 49787 10103 49793
rect 11149 49827 11207 49833
rect 11149 49793 11161 49827
rect 11195 49824 11207 49827
rect 11238 49824 11244 49836
rect 11195 49796 11244 49824
rect 11195 49793 11207 49796
rect 11149 49787 11207 49793
rect 11238 49784 11244 49796
rect 11296 49784 11302 49836
rect 3602 49716 3608 49768
rect 3660 49756 3666 49768
rect 4154 49756 4160 49768
rect 3660 49728 4160 49756
rect 3660 49716 3666 49728
rect 4154 49716 4160 49728
rect 4212 49716 4218 49768
rect 6822 49716 6828 49768
rect 6880 49756 6886 49768
rect 9953 49759 10011 49765
rect 6880 49728 9536 49756
rect 6880 49716 6886 49728
rect 2406 49648 2412 49700
rect 2464 49688 2470 49700
rect 7006 49688 7012 49700
rect 2464 49660 7012 49688
rect 2464 49648 2470 49660
rect 7006 49648 7012 49660
rect 7064 49648 7070 49700
rect 8662 49648 8668 49700
rect 8720 49688 8726 49700
rect 9122 49688 9128 49700
rect 8720 49660 9128 49688
rect 8720 49648 8726 49660
rect 9122 49648 9128 49660
rect 9180 49648 9186 49700
rect 9508 49697 9536 49728
rect 9953 49725 9965 49759
rect 9999 49756 10011 49759
rect 11790 49756 11796 49768
rect 9999 49728 11796 49756
rect 9999 49725 10011 49728
rect 9953 49719 10011 49725
rect 11790 49716 11796 49728
rect 11848 49716 11854 49768
rect 9493 49691 9551 49697
rect 9493 49657 9505 49691
rect 9539 49657 9551 49691
rect 9493 49651 9551 49657
rect 2314 49580 2320 49632
rect 2372 49620 2378 49632
rect 7190 49620 7196 49632
rect 2372 49592 7196 49620
rect 2372 49580 2378 49592
rect 7190 49580 7196 49592
rect 7248 49580 7254 49632
rect 1104 49530 10856 49552
rect 1104 49478 2582 49530
rect 2634 49478 2646 49530
rect 2698 49478 2710 49530
rect 2762 49478 2774 49530
rect 2826 49478 2838 49530
rect 2890 49478 5845 49530
rect 5897 49478 5909 49530
rect 5961 49478 5973 49530
rect 6025 49478 6037 49530
rect 6089 49478 6101 49530
rect 6153 49478 9109 49530
rect 9161 49478 9173 49530
rect 9225 49478 9237 49530
rect 9289 49478 9301 49530
rect 9353 49478 9365 49530
rect 9417 49478 10856 49530
rect 1104 49456 10856 49478
rect 3786 49376 3792 49428
rect 3844 49416 3850 49428
rect 6638 49416 6644 49428
rect 3844 49388 6644 49416
rect 3844 49376 3850 49388
rect 6638 49376 6644 49388
rect 6696 49376 6702 49428
rect 8205 49419 8263 49425
rect 8205 49385 8217 49419
rect 8251 49416 8263 49419
rect 8938 49416 8944 49428
rect 8251 49388 8944 49416
rect 8251 49385 8263 49388
rect 8205 49379 8263 49385
rect 8938 49376 8944 49388
rect 8996 49376 9002 49428
rect 2041 49351 2099 49357
rect 2041 49317 2053 49351
rect 2087 49348 2099 49351
rect 4062 49348 4068 49360
rect 2087 49320 4068 49348
rect 2087 49317 2099 49320
rect 2041 49311 2099 49317
rect 4062 49308 4068 49320
rect 4120 49308 4126 49360
rect 9766 49348 9772 49360
rect 9232 49320 9772 49348
rect 7190 49240 7196 49292
rect 7248 49280 7254 49292
rect 9232 49289 9260 49320
rect 9766 49308 9772 49320
rect 9824 49308 9830 49360
rect 10962 49348 10968 49360
rect 10923 49320 10968 49348
rect 10962 49308 10968 49320
rect 11020 49308 11026 49360
rect 9217 49283 9275 49289
rect 9217 49280 9229 49283
rect 7248 49252 9229 49280
rect 7248 49240 7254 49252
rect 9217 49249 9229 49252
rect 9263 49249 9275 49283
rect 9582 49280 9588 49292
rect 9217 49243 9275 49249
rect 9324 49252 9588 49280
rect 1854 49212 1860 49224
rect 1815 49184 1860 49212
rect 1854 49172 1860 49184
rect 1912 49172 1918 49224
rect 8202 49172 8208 49224
rect 8260 49212 8266 49224
rect 9324 49221 9352 49252
rect 9582 49240 9588 49252
rect 9640 49240 9646 49292
rect 8389 49215 8447 49221
rect 8389 49212 8401 49215
rect 8260 49184 8401 49212
rect 8260 49172 8266 49184
rect 8389 49181 8401 49184
rect 8435 49181 8447 49215
rect 8389 49175 8447 49181
rect 9309 49215 9367 49221
rect 9309 49181 9321 49215
rect 9355 49181 9367 49215
rect 9309 49175 9367 49181
rect 9398 49172 9404 49224
rect 9456 49212 9462 49224
rect 9493 49215 9551 49221
rect 9493 49212 9505 49215
rect 9456 49184 9505 49212
rect 9456 49172 9462 49184
rect 9493 49181 9505 49184
rect 9539 49181 9551 49215
rect 9493 49175 9551 49181
rect 9953 49147 10011 49153
rect 9953 49113 9965 49147
rect 9999 49144 10011 49147
rect 10965 49147 11023 49153
rect 10965 49144 10977 49147
rect 9999 49116 10977 49144
rect 9999 49113 10011 49116
rect 9953 49107 10011 49113
rect 10965 49113 10977 49116
rect 11011 49113 11023 49147
rect 10965 49107 11023 49113
rect 566 49036 572 49088
rect 624 49076 630 49088
rect 11146 49076 11152 49088
rect 624 49048 11152 49076
rect 624 49036 630 49048
rect 11146 49036 11152 49048
rect 11204 49036 11210 49088
rect 1104 48986 10856 49008
rect 1104 48934 4213 48986
rect 4265 48934 4277 48986
rect 4329 48934 4341 48986
rect 4393 48934 4405 48986
rect 4457 48934 4469 48986
rect 4521 48934 7477 48986
rect 7529 48934 7541 48986
rect 7593 48934 7605 48986
rect 7657 48934 7669 48986
rect 7721 48934 7733 48986
rect 7785 48934 10856 48986
rect 1104 48912 10856 48934
rect 8113 48875 8171 48881
rect 8113 48841 8125 48875
rect 8159 48872 8171 48875
rect 9490 48872 9496 48884
rect 8159 48844 9496 48872
rect 8159 48841 8171 48844
rect 8113 48835 8171 48841
rect 9490 48832 9496 48844
rect 9548 48832 9554 48884
rect 2041 48807 2099 48813
rect 2041 48773 2053 48807
rect 2087 48804 2099 48807
rect 5074 48804 5080 48816
rect 2087 48776 5080 48804
rect 2087 48773 2099 48776
rect 2041 48767 2099 48773
rect 5074 48764 5080 48776
rect 5132 48764 5138 48816
rect 1854 48736 1860 48748
rect 1815 48708 1860 48736
rect 1854 48696 1860 48708
rect 1912 48696 1918 48748
rect 8202 48696 8208 48748
rect 8260 48736 8266 48748
rect 8297 48739 8355 48745
rect 8297 48736 8309 48739
rect 8260 48708 8309 48736
rect 8260 48696 8266 48708
rect 8297 48705 8309 48708
rect 8343 48705 8355 48739
rect 8297 48699 8355 48705
rect 8938 48696 8944 48748
rect 8996 48736 9002 48748
rect 9125 48739 9183 48745
rect 9125 48736 9137 48739
rect 8996 48708 9137 48736
rect 8996 48696 9002 48708
rect 9125 48705 9137 48708
rect 9171 48705 9183 48739
rect 9125 48699 9183 48705
rect 9309 48739 9367 48745
rect 9309 48705 9321 48739
rect 9355 48736 9367 48739
rect 9398 48736 9404 48748
rect 9355 48708 9404 48736
rect 9355 48705 9367 48708
rect 9309 48699 9367 48705
rect 9398 48696 9404 48708
rect 9456 48736 9462 48748
rect 9950 48736 9956 48748
rect 9456 48708 9956 48736
rect 9456 48696 9462 48708
rect 9950 48696 9956 48708
rect 10008 48696 10014 48748
rect 1578 48628 1584 48680
rect 1636 48668 1642 48680
rect 8846 48668 8852 48680
rect 1636 48640 8852 48668
rect 1636 48628 1642 48640
rect 8846 48628 8852 48640
rect 8904 48668 8910 48680
rect 9033 48671 9091 48677
rect 9033 48668 9045 48671
rect 8904 48640 9045 48668
rect 8904 48628 8910 48640
rect 9033 48637 9045 48640
rect 9079 48637 9091 48671
rect 9033 48631 9091 48637
rect 9769 48671 9827 48677
rect 9769 48637 9781 48671
rect 9815 48668 9827 48671
rect 10778 48668 10784 48680
rect 9815 48640 10784 48668
rect 9815 48637 9827 48640
rect 9769 48631 9827 48637
rect 10778 48628 10784 48640
rect 10836 48628 10842 48680
rect 1104 48442 10856 48464
rect 1104 48390 2582 48442
rect 2634 48390 2646 48442
rect 2698 48390 2710 48442
rect 2762 48390 2774 48442
rect 2826 48390 2838 48442
rect 2890 48390 5845 48442
rect 5897 48390 5909 48442
rect 5961 48390 5973 48442
rect 6025 48390 6037 48442
rect 6089 48390 6101 48442
rect 6153 48390 9109 48442
rect 9161 48390 9173 48442
rect 9225 48390 9237 48442
rect 9289 48390 9301 48442
rect 9353 48390 9365 48442
rect 9417 48390 10856 48442
rect 1104 48368 10856 48390
rect 5350 48288 5356 48340
rect 5408 48288 5414 48340
rect 8846 48288 8852 48340
rect 8904 48328 8910 48340
rect 9030 48328 9036 48340
rect 8904 48300 9036 48328
rect 8904 48288 8910 48300
rect 9030 48288 9036 48300
rect 9088 48288 9094 48340
rect 2038 48260 2044 48272
rect 1999 48232 2044 48260
rect 2038 48220 2044 48232
rect 2096 48220 2102 48272
rect 2130 48220 2136 48272
rect 2188 48260 2194 48272
rect 5368 48260 5396 48288
rect 9582 48260 9588 48272
rect 2188 48232 5396 48260
rect 9324 48232 9588 48260
rect 2188 48220 2194 48232
rect 4706 48152 4712 48204
rect 4764 48152 4770 48204
rect 8754 48152 8760 48204
rect 8812 48192 8818 48204
rect 9030 48192 9036 48204
rect 8812 48164 9036 48192
rect 8812 48152 8818 48164
rect 9030 48152 9036 48164
rect 9088 48152 9094 48204
rect 4724 48124 4752 48152
rect 5258 48124 5264 48136
rect 4724 48096 5264 48124
rect 5258 48084 5264 48096
rect 5316 48084 5322 48136
rect 8202 48084 8208 48136
rect 8260 48124 8266 48136
rect 8389 48127 8447 48133
rect 8389 48124 8401 48127
rect 8260 48096 8401 48124
rect 8260 48084 8266 48096
rect 8389 48093 8401 48096
rect 8435 48093 8447 48127
rect 8389 48087 8447 48093
rect 8846 48084 8852 48136
rect 8904 48124 8910 48136
rect 9324 48133 9352 48232
rect 9582 48220 9588 48232
rect 9640 48220 9646 48272
rect 9309 48127 9367 48133
rect 9309 48124 9321 48127
rect 8904 48096 9321 48124
rect 8904 48084 8910 48096
rect 9309 48093 9321 48096
rect 9355 48093 9367 48127
rect 9309 48087 9367 48093
rect 9401 48127 9459 48133
rect 9401 48093 9413 48127
rect 9447 48124 9459 48127
rect 9490 48124 9496 48136
rect 9447 48096 9496 48124
rect 9447 48093 9459 48096
rect 9401 48087 9459 48093
rect 9490 48084 9496 48096
rect 9548 48084 9554 48136
rect 9585 48127 9643 48133
rect 9585 48093 9597 48127
rect 9631 48124 9643 48127
rect 9950 48124 9956 48136
rect 9631 48096 9956 48124
rect 9631 48093 9643 48096
rect 9585 48087 9643 48093
rect 9950 48084 9956 48096
rect 10008 48084 10014 48136
rect 11238 48084 11244 48136
rect 11296 48124 11302 48136
rect 11606 48124 11612 48136
rect 11296 48096 11612 48124
rect 11296 48084 11302 48096
rect 11606 48084 11612 48096
rect 11664 48084 11670 48136
rect 1854 48056 1860 48068
rect 1815 48028 1860 48056
rect 1854 48016 1860 48028
rect 1912 48016 1918 48068
rect 4706 48016 4712 48068
rect 4764 48056 4770 48068
rect 10045 48059 10103 48065
rect 10045 48056 10057 48059
rect 4764 48028 10057 48056
rect 4764 48016 4770 48028
rect 10045 48025 10057 48028
rect 10091 48025 10103 48059
rect 10045 48019 10103 48025
rect 8205 47991 8263 47997
rect 8205 47957 8217 47991
rect 8251 47988 8263 47991
rect 9674 47988 9680 48000
rect 8251 47960 9680 47988
rect 8251 47957 8263 47960
rect 8205 47951 8263 47957
rect 9674 47948 9680 47960
rect 9732 47948 9738 48000
rect 11606 47988 11612 48000
rect 11567 47960 11612 47988
rect 11606 47948 11612 47960
rect 11664 47948 11670 48000
rect 1104 47898 10856 47920
rect 1104 47846 4213 47898
rect 4265 47846 4277 47898
rect 4329 47846 4341 47898
rect 4393 47846 4405 47898
rect 4457 47846 4469 47898
rect 4521 47846 7477 47898
rect 7529 47846 7541 47898
rect 7593 47846 7605 47898
rect 7657 47846 7669 47898
rect 7721 47846 7733 47898
rect 7785 47846 10856 47898
rect 1104 47824 10856 47846
rect 11425 47855 11483 47861
rect 11425 47821 11437 47855
rect 11471 47852 11483 47855
rect 11609 47855 11667 47861
rect 11609 47852 11621 47855
rect 11471 47824 11621 47852
rect 11471 47821 11483 47824
rect 11425 47815 11483 47821
rect 11609 47821 11621 47824
rect 11655 47821 11667 47855
rect 11609 47815 11667 47821
rect 1946 47784 1952 47796
rect 1907 47756 1952 47784
rect 1946 47744 1952 47756
rect 2004 47744 2010 47796
rect 2222 47744 2228 47796
rect 2280 47784 2286 47796
rect 4709 47787 4767 47793
rect 4709 47784 4721 47787
rect 2280 47756 4721 47784
rect 2280 47744 2286 47756
rect 4709 47753 4721 47756
rect 4755 47753 4767 47787
rect 5074 47784 5080 47796
rect 4987 47756 5080 47784
rect 4709 47747 4767 47753
rect 5074 47744 5080 47756
rect 5132 47784 5138 47796
rect 9033 47787 9091 47793
rect 9033 47784 9045 47787
rect 5132 47756 9045 47784
rect 5132 47744 5138 47756
rect 9033 47753 9045 47756
rect 9079 47753 9091 47787
rect 9033 47747 9091 47753
rect 9214 47744 9220 47796
rect 9272 47784 9278 47796
rect 10042 47784 10048 47796
rect 9272 47756 10048 47784
rect 9272 47744 9278 47756
rect 10042 47744 10048 47756
rect 10100 47744 10106 47796
rect 3602 47676 3608 47728
rect 3660 47716 3666 47728
rect 9674 47716 9680 47728
rect 3660 47688 5672 47716
rect 9587 47688 9680 47716
rect 3660 47676 3666 47688
rect 1854 47648 1860 47660
rect 1815 47620 1860 47648
rect 1854 47608 1860 47620
rect 1912 47608 1918 47660
rect 750 47540 756 47592
rect 808 47580 814 47592
rect 4706 47580 4712 47592
rect 808 47552 4712 47580
rect 808 47540 814 47552
rect 4706 47540 4712 47552
rect 4764 47540 4770 47592
rect 5169 47583 5227 47589
rect 5169 47549 5181 47583
rect 5215 47549 5227 47583
rect 5169 47543 5227 47549
rect 5353 47583 5411 47589
rect 5353 47549 5365 47583
rect 5399 47580 5411 47583
rect 5399 47552 5580 47580
rect 5399 47549 5411 47552
rect 5353 47543 5411 47549
rect 2866 47472 2872 47524
rect 2924 47512 2930 47524
rect 3602 47512 3608 47524
rect 2924 47484 3608 47512
rect 2924 47472 2930 47484
rect 3602 47472 3608 47484
rect 3660 47472 3666 47524
rect 4706 47404 4712 47456
rect 4764 47444 4770 47456
rect 5184 47444 5212 47543
rect 4764 47416 5212 47444
rect 5552 47444 5580 47552
rect 5644 47512 5672 47688
rect 9674 47676 9680 47688
rect 9732 47716 9738 47728
rect 11425 47719 11483 47725
rect 11425 47716 11437 47719
rect 9732 47688 11437 47716
rect 9732 47676 9738 47688
rect 11425 47685 11437 47688
rect 11471 47685 11483 47719
rect 11425 47679 11483 47685
rect 8849 47651 8907 47657
rect 8849 47617 8861 47651
rect 8895 47617 8907 47651
rect 8849 47611 8907 47617
rect 9217 47651 9275 47657
rect 9217 47617 9229 47651
rect 9263 47648 9275 47651
rect 9582 47648 9588 47660
rect 9263 47620 9588 47648
rect 9263 47617 9275 47620
rect 9217 47611 9275 47617
rect 8864 47580 8892 47611
rect 9582 47608 9588 47620
rect 9640 47608 9646 47660
rect 9769 47651 9827 47657
rect 9769 47617 9781 47651
rect 9815 47648 9827 47651
rect 9858 47648 9864 47660
rect 9815 47620 9864 47648
rect 9815 47617 9827 47620
rect 9769 47611 9827 47617
rect 9858 47608 9864 47620
rect 9916 47608 9922 47660
rect 10226 47608 10232 47660
rect 10284 47648 10290 47660
rect 10321 47651 10379 47657
rect 10321 47648 10333 47651
rect 10284 47620 10333 47648
rect 10284 47608 10290 47620
rect 10321 47617 10333 47620
rect 10367 47617 10379 47651
rect 10321 47611 10379 47617
rect 9490 47580 9496 47592
rect 8864 47552 9496 47580
rect 9490 47540 9496 47552
rect 9548 47540 9554 47592
rect 9950 47580 9956 47592
rect 9911 47552 9956 47580
rect 9950 47540 9956 47552
rect 10008 47540 10014 47592
rect 9309 47515 9367 47521
rect 9309 47512 9321 47515
rect 5644 47484 9321 47512
rect 9309 47481 9321 47484
rect 9355 47481 9367 47515
rect 9309 47475 9367 47481
rect 5718 47444 5724 47456
rect 5552 47416 5724 47444
rect 4764 47404 4770 47416
rect 5718 47404 5724 47416
rect 5776 47404 5782 47456
rect 8662 47444 8668 47456
rect 8623 47416 8668 47444
rect 8662 47404 8668 47416
rect 8720 47404 8726 47456
rect 10042 47404 10048 47456
rect 10100 47444 10106 47456
rect 10137 47447 10195 47453
rect 10137 47444 10149 47447
rect 10100 47416 10149 47444
rect 10100 47404 10106 47416
rect 10137 47413 10149 47416
rect 10183 47413 10195 47447
rect 10137 47407 10195 47413
rect 1104 47354 10856 47376
rect 1104 47302 2582 47354
rect 2634 47302 2646 47354
rect 2698 47302 2710 47354
rect 2762 47302 2774 47354
rect 2826 47302 2838 47354
rect 2890 47302 5845 47354
rect 5897 47302 5909 47354
rect 5961 47302 5973 47354
rect 6025 47302 6037 47354
rect 6089 47302 6101 47354
rect 6153 47302 9109 47354
rect 9161 47302 9173 47354
rect 9225 47302 9237 47354
rect 9289 47302 9301 47354
rect 9353 47302 9365 47354
rect 9417 47302 10856 47354
rect 1104 47280 10856 47302
rect 1118 47200 1124 47252
rect 1176 47240 1182 47252
rect 1949 47243 2007 47249
rect 1949 47240 1961 47243
rect 1176 47212 1961 47240
rect 1176 47200 1182 47212
rect 1949 47209 1961 47212
rect 1995 47209 2007 47243
rect 1949 47203 2007 47209
rect 4062 47200 4068 47252
rect 4120 47240 4126 47252
rect 9401 47243 9459 47249
rect 9401 47240 9413 47243
rect 4120 47212 9413 47240
rect 4120 47200 4126 47212
rect 9401 47209 9413 47212
rect 9447 47209 9459 47243
rect 9401 47203 9459 47209
rect 10870 47200 10876 47252
rect 10928 47240 10934 47252
rect 10965 47243 11023 47249
rect 10965 47240 10977 47243
rect 10928 47212 10977 47240
rect 10928 47200 10934 47212
rect 10965 47209 10977 47212
rect 11011 47209 11023 47243
rect 10965 47203 11023 47209
rect 8205 47175 8263 47181
rect 8205 47141 8217 47175
rect 8251 47172 8263 47175
rect 9766 47172 9772 47184
rect 8251 47144 9772 47172
rect 8251 47141 8263 47144
rect 8205 47135 8263 47141
rect 9766 47132 9772 47144
rect 9824 47132 9830 47184
rect 6638 47064 6644 47116
rect 6696 47104 6702 47116
rect 8846 47104 8852 47116
rect 6696 47076 8852 47104
rect 6696 47064 6702 47076
rect 8846 47064 8852 47076
rect 8904 47064 8910 47116
rect 9398 47064 9404 47116
rect 9456 47104 9462 47116
rect 9950 47104 9956 47116
rect 9456 47076 9956 47104
rect 9456 47064 9462 47076
rect 9950 47064 9956 47076
rect 10008 47064 10014 47116
rect 10965 47107 11023 47113
rect 10965 47073 10977 47107
rect 11011 47104 11023 47107
rect 11149 47107 11207 47113
rect 11149 47104 11161 47107
rect 11011 47076 11161 47104
rect 11011 47073 11023 47076
rect 10965 47067 11023 47073
rect 11149 47073 11161 47076
rect 11195 47073 11207 47107
rect 11149 47067 11207 47073
rect 8202 46996 8208 47048
rect 8260 47036 8266 47048
rect 8389 47039 8447 47045
rect 8389 47036 8401 47039
rect 8260 47008 8401 47036
rect 8260 46996 8266 47008
rect 8389 47005 8401 47008
rect 8435 47005 8447 47039
rect 8389 46999 8447 47005
rect 1854 46968 1860 46980
rect 1815 46940 1860 46968
rect 1854 46928 1860 46940
rect 1912 46928 1918 46980
rect 8662 46928 8668 46980
rect 8720 46968 8726 46980
rect 9769 46971 9827 46977
rect 9769 46968 9781 46971
rect 8720 46940 9781 46968
rect 8720 46928 8726 46940
rect 9769 46937 9781 46940
rect 9815 46968 9827 46971
rect 11149 46971 11207 46977
rect 11149 46968 11161 46971
rect 9815 46940 11161 46968
rect 9815 46937 9827 46940
rect 9769 46931 9827 46937
rect 11149 46937 11161 46940
rect 11195 46937 11207 46971
rect 11149 46931 11207 46937
rect 9674 46860 9680 46912
rect 9732 46900 9738 46912
rect 9861 46903 9919 46909
rect 9861 46900 9873 46903
rect 9732 46872 9873 46900
rect 9732 46860 9738 46872
rect 9861 46869 9873 46872
rect 9907 46869 9919 46903
rect 9861 46863 9919 46869
rect 1104 46810 10856 46832
rect 1104 46758 4213 46810
rect 4265 46758 4277 46810
rect 4329 46758 4341 46810
rect 4393 46758 4405 46810
rect 4457 46758 4469 46810
rect 4521 46758 7477 46810
rect 7529 46758 7541 46810
rect 7593 46758 7605 46810
rect 7657 46758 7669 46810
rect 7721 46758 7733 46810
rect 7785 46758 10856 46810
rect 1104 46736 10856 46758
rect 5534 46656 5540 46708
rect 5592 46696 5598 46708
rect 9401 46699 9459 46705
rect 9401 46696 9413 46699
rect 5592 46668 9413 46696
rect 5592 46656 5598 46668
rect 9401 46665 9413 46668
rect 9447 46665 9459 46699
rect 9766 46696 9772 46708
rect 9727 46668 9772 46696
rect 9401 46659 9459 46665
rect 9766 46656 9772 46668
rect 9824 46656 9830 46708
rect 4062 46588 4068 46640
rect 4120 46628 4126 46640
rect 5718 46628 5724 46640
rect 4120 46600 5724 46628
rect 4120 46588 4126 46600
rect 5074 46560 5080 46572
rect 5035 46532 5080 46560
rect 5074 46520 5080 46532
rect 5132 46520 5138 46572
rect 5276 46569 5304 46600
rect 5718 46588 5724 46600
rect 5776 46588 5782 46640
rect 8110 46588 8116 46640
rect 8168 46628 8174 46640
rect 8665 46631 8723 46637
rect 8665 46628 8677 46631
rect 8168 46600 8677 46628
rect 8168 46588 8174 46600
rect 8665 46597 8677 46600
rect 8711 46597 8723 46631
rect 8665 46591 8723 46597
rect 9508 46600 9674 46628
rect 5261 46563 5319 46569
rect 5261 46529 5273 46563
rect 5307 46529 5319 46563
rect 5261 46523 5319 46529
rect 8481 46563 8539 46569
rect 8481 46529 8493 46563
rect 8527 46560 8539 46563
rect 9508 46560 9536 46600
rect 8527 46532 9536 46560
rect 9646 46560 9674 46600
rect 11238 46560 11244 46572
rect 9646 46532 11244 46560
rect 8527 46529 8539 46532
rect 8481 46523 8539 46529
rect 11238 46520 11244 46532
rect 11296 46520 11302 46572
rect 4706 46452 4712 46504
rect 4764 46492 4770 46504
rect 4985 46495 5043 46501
rect 4985 46492 4997 46495
rect 4764 46464 4997 46492
rect 4764 46452 4770 46464
rect 4985 46461 4997 46464
rect 5031 46461 5043 46495
rect 5718 46492 5724 46504
rect 5679 46464 5724 46492
rect 4985 46455 5043 46461
rect 5000 46356 5028 46455
rect 5718 46452 5724 46464
rect 5776 46452 5782 46504
rect 8757 46495 8815 46501
rect 8757 46461 8769 46495
rect 8803 46492 8815 46495
rect 9398 46492 9404 46504
rect 8803 46464 9404 46492
rect 8803 46461 8815 46464
rect 8757 46455 8815 46461
rect 9398 46452 9404 46464
rect 9456 46452 9462 46504
rect 9490 46452 9496 46504
rect 9548 46492 9554 46504
rect 9861 46495 9919 46501
rect 9861 46492 9873 46495
rect 9548 46464 9873 46492
rect 9548 46452 9554 46464
rect 9861 46461 9873 46464
rect 9907 46461 9919 46495
rect 9861 46455 9919 46461
rect 9953 46495 10011 46501
rect 9953 46461 9965 46495
rect 9999 46461 10011 46495
rect 9953 46455 10011 46461
rect 8018 46384 8024 46436
rect 8076 46424 8082 46436
rect 8205 46427 8263 46433
rect 8205 46424 8217 46427
rect 8076 46396 8217 46424
rect 8076 46384 8082 46396
rect 8205 46393 8217 46396
rect 8251 46393 8263 46427
rect 8205 46387 8263 46393
rect 8570 46384 8576 46436
rect 8628 46424 8634 46436
rect 8846 46424 8852 46436
rect 8628 46396 8852 46424
rect 8628 46384 8634 46396
rect 8846 46384 8852 46396
rect 8904 46384 8910 46436
rect 9416 46424 9444 46452
rect 9582 46424 9588 46436
rect 9416 46396 9588 46424
rect 9582 46384 9588 46396
rect 9640 46424 9646 46436
rect 9968 46424 9996 46455
rect 9640 46396 9996 46424
rect 9640 46384 9646 46396
rect 9950 46356 9956 46368
rect 5000 46328 9956 46356
rect 9950 46316 9956 46328
rect 10008 46316 10014 46368
rect 1104 46266 10856 46288
rect 1104 46214 2582 46266
rect 2634 46214 2646 46266
rect 2698 46214 2710 46266
rect 2762 46214 2774 46266
rect 2826 46214 2838 46266
rect 2890 46214 5845 46266
rect 5897 46214 5909 46266
rect 5961 46214 5973 46266
rect 6025 46214 6037 46266
rect 6089 46214 6101 46266
rect 6153 46214 9109 46266
rect 9161 46214 9173 46266
rect 9225 46214 9237 46266
rect 9289 46214 9301 46266
rect 9353 46214 9365 46266
rect 9417 46214 10856 46266
rect 1104 46192 10856 46214
rect 1302 46112 1308 46164
rect 1360 46152 1366 46164
rect 1949 46155 2007 46161
rect 1949 46152 1961 46155
rect 1360 46124 1961 46152
rect 1360 46112 1366 46124
rect 1949 46121 1961 46124
rect 1995 46121 2007 46155
rect 1949 46115 2007 46121
rect 7006 46112 7012 46164
rect 7064 46112 7070 46164
rect 10226 46112 10232 46164
rect 10284 46152 10290 46164
rect 10410 46152 10416 46164
rect 10284 46124 10416 46152
rect 10284 46112 10290 46124
rect 10410 46112 10416 46124
rect 10468 46112 10474 46164
rect 7024 46016 7052 46112
rect 8662 46044 8668 46096
rect 8720 46084 8726 46096
rect 9493 46087 9551 46093
rect 9493 46084 9505 46087
rect 8720 46056 9505 46084
rect 8720 46044 8726 46056
rect 9493 46053 9505 46056
rect 9539 46053 9551 46087
rect 9493 46047 9551 46053
rect 6932 45988 7052 46016
rect 6932 45960 6960 45988
rect 9582 45976 9588 46028
rect 9640 46016 9646 46028
rect 9640 45988 10088 46016
rect 9640 45976 9646 45988
rect 1854 45948 1860 45960
rect 1815 45920 1860 45948
rect 1854 45908 1860 45920
rect 1912 45908 1918 45960
rect 6914 45908 6920 45960
rect 6972 45908 6978 45960
rect 7006 45908 7012 45960
rect 7064 45948 7070 45960
rect 8202 45948 8208 45960
rect 7064 45920 8208 45948
rect 7064 45908 7070 45920
rect 8202 45908 8208 45920
rect 8260 45908 8266 45960
rect 9582 45840 9588 45892
rect 9640 45880 9646 45892
rect 10060 45889 10088 45988
rect 9769 45883 9827 45889
rect 9769 45880 9781 45883
rect 9640 45852 9781 45880
rect 9640 45840 9646 45852
rect 9769 45849 9781 45852
rect 9815 45849 9827 45883
rect 9769 45843 9827 45849
rect 10045 45883 10103 45889
rect 10045 45849 10057 45883
rect 10091 45880 10103 45883
rect 10410 45880 10416 45892
rect 10091 45852 10416 45880
rect 10091 45849 10103 45852
rect 10045 45843 10103 45849
rect 10410 45840 10416 45852
rect 10468 45840 10474 45892
rect 9950 45812 9956 45824
rect 9911 45784 9956 45812
rect 9950 45772 9956 45784
rect 10008 45772 10014 45824
rect 1104 45722 10856 45744
rect 1104 45670 4213 45722
rect 4265 45670 4277 45722
rect 4329 45670 4341 45722
rect 4393 45670 4405 45722
rect 4457 45670 4469 45722
rect 4521 45670 7477 45722
rect 7529 45670 7541 45722
rect 7593 45670 7605 45722
rect 7657 45670 7669 45722
rect 7721 45670 7733 45722
rect 7785 45670 10856 45722
rect 1104 45648 10856 45670
rect 3878 45568 3884 45620
rect 3936 45608 3942 45620
rect 5166 45608 5172 45620
rect 3936 45580 5172 45608
rect 3936 45568 3942 45580
rect 5166 45568 5172 45580
rect 5224 45568 5230 45620
rect 9950 45568 9956 45620
rect 10008 45608 10014 45620
rect 10321 45611 10379 45617
rect 10321 45608 10333 45611
rect 10008 45580 10333 45608
rect 10008 45568 10014 45580
rect 10321 45577 10333 45580
rect 10367 45608 10379 45611
rect 11698 45608 11704 45620
rect 10367 45580 11704 45608
rect 10367 45577 10379 45580
rect 10321 45571 10379 45577
rect 11698 45568 11704 45580
rect 11756 45568 11762 45620
rect 1946 45500 1952 45552
rect 2004 45540 2010 45552
rect 2314 45540 2320 45552
rect 2004 45512 2320 45540
rect 2004 45500 2010 45512
rect 2314 45500 2320 45512
rect 2372 45500 2378 45552
rect 3329 45543 3387 45549
rect 3329 45509 3341 45543
rect 3375 45540 3387 45543
rect 4706 45540 4712 45552
rect 3375 45512 4712 45540
rect 3375 45509 3387 45512
rect 3329 45503 3387 45509
rect 4706 45500 4712 45512
rect 4764 45540 4770 45552
rect 10042 45540 10048 45552
rect 4764 45512 10048 45540
rect 4764 45500 4770 45512
rect 10042 45500 10048 45512
rect 10100 45500 10106 45552
rect 1394 45472 1400 45484
rect 1355 45444 1400 45472
rect 1394 45432 1400 45444
rect 1452 45432 1458 45484
rect 3421 45475 3479 45481
rect 3421 45441 3433 45475
rect 3467 45472 3479 45475
rect 4062 45472 4068 45484
rect 3467 45444 4068 45472
rect 3467 45441 3479 45444
rect 3421 45435 3479 45441
rect 4062 45432 4068 45444
rect 4120 45432 4126 45484
rect 8202 45432 8208 45484
rect 8260 45472 8266 45484
rect 8665 45475 8723 45481
rect 8665 45472 8677 45475
rect 8260 45444 8677 45472
rect 8260 45432 8266 45444
rect 8665 45441 8677 45444
rect 8711 45441 8723 45475
rect 8665 45435 8723 45441
rect 10962 45432 10968 45484
rect 11020 45472 11026 45484
rect 11698 45472 11704 45484
rect 11020 45444 11704 45472
rect 11020 45432 11026 45444
rect 11698 45432 11704 45444
rect 11756 45432 11762 45484
rect 1762 45364 1768 45416
rect 1820 45404 1826 45416
rect 2222 45404 2228 45416
rect 1820 45376 2228 45404
rect 1820 45364 1826 45376
rect 2222 45364 2228 45376
rect 2280 45364 2286 45416
rect 3605 45407 3663 45413
rect 3605 45373 3617 45407
rect 3651 45404 3663 45407
rect 4154 45404 4160 45416
rect 3651 45376 4160 45404
rect 3651 45373 3663 45376
rect 3605 45367 3663 45373
rect 4154 45364 4160 45376
rect 4212 45364 4218 45416
rect 1486 45296 1492 45348
rect 1544 45336 1550 45348
rect 2961 45339 3019 45345
rect 2961 45336 2973 45339
rect 1544 45308 2973 45336
rect 1544 45296 1550 45308
rect 2961 45305 2973 45308
rect 3007 45305 3019 45339
rect 2961 45299 3019 45305
rect 8754 45296 8760 45348
rect 8812 45336 8818 45348
rect 9217 45339 9275 45345
rect 9217 45336 9229 45339
rect 8812 45308 9229 45336
rect 8812 45296 8818 45308
rect 9217 45305 9229 45308
rect 9263 45336 9275 45339
rect 9582 45336 9588 45348
rect 9263 45308 9588 45336
rect 9263 45305 9275 45308
rect 9217 45299 9275 45305
rect 9582 45296 9588 45308
rect 9640 45296 9646 45348
rect 1581 45271 1639 45277
rect 1581 45237 1593 45271
rect 1627 45268 1639 45271
rect 7282 45268 7288 45280
rect 1627 45240 7288 45268
rect 1627 45237 1639 45240
rect 1581 45231 1639 45237
rect 7282 45228 7288 45240
rect 7340 45228 7346 45280
rect 8849 45271 8907 45277
rect 8849 45237 8861 45271
rect 8895 45268 8907 45271
rect 11238 45268 11244 45280
rect 8895 45240 11244 45268
rect 8895 45237 8907 45240
rect 8849 45231 8907 45237
rect 11238 45228 11244 45240
rect 11296 45228 11302 45280
rect 1104 45178 10856 45200
rect 1104 45126 2582 45178
rect 2634 45126 2646 45178
rect 2698 45126 2710 45178
rect 2762 45126 2774 45178
rect 2826 45126 2838 45178
rect 2890 45126 5845 45178
rect 5897 45126 5909 45178
rect 5961 45126 5973 45178
rect 6025 45126 6037 45178
rect 6089 45126 6101 45178
rect 6153 45126 9109 45178
rect 9161 45126 9173 45178
rect 9225 45126 9237 45178
rect 9289 45126 9301 45178
rect 9353 45126 9365 45178
rect 9417 45126 10856 45178
rect 1104 45104 10856 45126
rect 1578 45024 1584 45076
rect 1636 45064 1642 45076
rect 1762 45064 1768 45076
rect 1636 45036 1768 45064
rect 1636 45024 1642 45036
rect 1762 45024 1768 45036
rect 1820 45024 1826 45076
rect 9582 45024 9588 45076
rect 9640 45064 9646 45076
rect 9858 45064 9864 45076
rect 9640 45036 9864 45064
rect 9640 45024 9646 45036
rect 9858 45024 9864 45036
rect 9916 45024 9922 45076
rect 2041 44999 2099 45005
rect 2041 44965 2053 44999
rect 2087 44996 2099 44999
rect 3326 44996 3332 45008
rect 2087 44968 3332 44996
rect 2087 44965 2099 44968
rect 2041 44959 2099 44965
rect 3326 44956 3332 44968
rect 3384 44956 3390 45008
rect 9766 44928 9772 44940
rect 9508 44900 9772 44928
rect 3326 44820 3332 44872
rect 3384 44860 3390 44872
rect 4154 44860 4160 44872
rect 3384 44832 4160 44860
rect 3384 44820 3390 44832
rect 4154 44820 4160 44832
rect 4212 44820 4218 44872
rect 9398 44860 9404 44872
rect 9359 44832 9404 44860
rect 9398 44820 9404 44832
rect 9456 44820 9462 44872
rect 9508 44869 9536 44900
rect 9766 44888 9772 44900
rect 9824 44888 9830 44940
rect 9493 44863 9551 44869
rect 9493 44829 9505 44863
rect 9539 44829 9551 44863
rect 9493 44823 9551 44829
rect 9677 44863 9735 44869
rect 9677 44829 9689 44863
rect 9723 44860 9735 44863
rect 9950 44860 9956 44872
rect 9723 44832 9956 44860
rect 9723 44829 9735 44832
rect 9677 44823 9735 44829
rect 9950 44820 9956 44832
rect 10008 44860 10014 44872
rect 10410 44860 10416 44872
rect 10008 44832 10416 44860
rect 10008 44820 10014 44832
rect 10410 44820 10416 44832
rect 10468 44820 10474 44872
rect 1854 44792 1860 44804
rect 1815 44764 1860 44792
rect 1854 44752 1860 44764
rect 1912 44752 1918 44804
rect 10134 44792 10140 44804
rect 10095 44764 10140 44792
rect 10134 44752 10140 44764
rect 10192 44752 10198 44804
rect 5626 44684 5632 44736
rect 5684 44724 5690 44736
rect 6362 44724 6368 44736
rect 5684 44696 6368 44724
rect 5684 44684 5690 44696
rect 6362 44684 6368 44696
rect 6420 44684 6426 44736
rect 7282 44684 7288 44736
rect 7340 44724 7346 44736
rect 8386 44724 8392 44736
rect 7340 44696 8392 44724
rect 7340 44684 7346 44696
rect 8386 44684 8392 44696
rect 8444 44684 8450 44736
rect 1104 44634 10856 44656
rect 1104 44582 4213 44634
rect 4265 44582 4277 44634
rect 4329 44582 4341 44634
rect 4393 44582 4405 44634
rect 4457 44582 4469 44634
rect 4521 44582 7477 44634
rect 7529 44582 7541 44634
rect 7593 44582 7605 44634
rect 7657 44582 7669 44634
rect 7721 44582 7733 44634
rect 7785 44582 10856 44634
rect 1104 44560 10856 44582
rect 9582 44480 9588 44532
rect 9640 44520 9646 44532
rect 10134 44520 10140 44532
rect 9640 44492 10140 44520
rect 9640 44480 9646 44492
rect 10134 44480 10140 44492
rect 10192 44480 10198 44532
rect 2041 44455 2099 44461
rect 2041 44421 2053 44455
rect 2087 44452 2099 44455
rect 3234 44452 3240 44464
rect 2087 44424 3240 44452
rect 2087 44421 2099 44424
rect 2041 44415 2099 44421
rect 3234 44412 3240 44424
rect 3292 44412 3298 44464
rect 8202 44412 8208 44464
rect 8260 44452 8266 44464
rect 11425 44455 11483 44461
rect 11425 44452 11437 44455
rect 8260 44412 8294 44452
rect 1854 44384 1860 44396
rect 1815 44356 1860 44384
rect 1854 44344 1860 44356
rect 1912 44344 1918 44396
rect 1578 44276 1584 44328
rect 1636 44316 1642 44328
rect 2498 44316 2504 44328
rect 1636 44288 2504 44316
rect 1636 44276 1642 44288
rect 2498 44276 2504 44288
rect 2556 44276 2562 44328
rect 2038 44208 2044 44260
rect 2096 44248 2102 44260
rect 5074 44248 5080 44260
rect 2096 44220 5080 44248
rect 2096 44208 2102 44220
rect 5074 44208 5080 44220
rect 5132 44208 5138 44260
rect 8266 44248 8294 44412
rect 9508 44424 11437 44452
rect 8389 44387 8447 44393
rect 8389 44353 8401 44387
rect 8435 44384 8447 44387
rect 9214 44384 9220 44396
rect 8435 44356 9220 44384
rect 8435 44353 8447 44356
rect 8389 44347 8447 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 9508 44393 9536 44424
rect 11425 44421 11437 44424
rect 11471 44421 11483 44455
rect 11425 44415 11483 44421
rect 9493 44387 9551 44393
rect 9493 44353 9505 44387
rect 9539 44353 9551 44387
rect 9493 44347 9551 44353
rect 9677 44387 9735 44393
rect 9677 44353 9689 44387
rect 9723 44384 9735 44387
rect 9950 44384 9956 44396
rect 9723 44356 9956 44384
rect 9723 44353 9735 44356
rect 9677 44347 9735 44353
rect 9398 44276 9404 44328
rect 9456 44316 9462 44328
rect 9692 44316 9720 44347
rect 9950 44344 9956 44356
rect 10008 44344 10014 44396
rect 9456 44288 9501 44316
rect 9600 44288 9720 44316
rect 9456 44276 9462 44288
rect 9600 44248 9628 44288
rect 10042 44276 10048 44328
rect 10100 44316 10106 44328
rect 10137 44319 10195 44325
rect 10137 44316 10149 44319
rect 10100 44288 10149 44316
rect 10100 44276 10106 44288
rect 10137 44285 10149 44288
rect 10183 44285 10195 44319
rect 10137 44279 10195 44285
rect 8266 44220 9628 44248
rect 2314 44140 2320 44192
rect 2372 44180 2378 44192
rect 3970 44180 3976 44192
rect 2372 44152 3976 44180
rect 2372 44140 2378 44152
rect 3970 44140 3976 44152
rect 4028 44140 4034 44192
rect 8386 44140 8392 44192
rect 8444 44180 8450 44192
rect 8573 44183 8631 44189
rect 8573 44180 8585 44183
rect 8444 44152 8585 44180
rect 8444 44140 8450 44152
rect 8573 44149 8585 44152
rect 8619 44149 8631 44183
rect 8573 44143 8631 44149
rect 1104 44090 10856 44112
rect 1104 44038 2582 44090
rect 2634 44038 2646 44090
rect 2698 44038 2710 44090
rect 2762 44038 2774 44090
rect 2826 44038 2838 44090
rect 2890 44038 5845 44090
rect 5897 44038 5909 44090
rect 5961 44038 5973 44090
rect 6025 44038 6037 44090
rect 6089 44038 6101 44090
rect 6153 44038 9109 44090
rect 9161 44038 9173 44090
rect 9225 44038 9237 44090
rect 9289 44038 9301 44090
rect 9353 44038 9365 44090
rect 9417 44038 10856 44090
rect 1104 44016 10856 44038
rect 382 43936 388 43988
rect 440 43976 446 43988
rect 1486 43976 1492 43988
rect 440 43948 1492 43976
rect 440 43936 446 43948
rect 1486 43936 1492 43948
rect 1544 43936 1550 43988
rect 7558 43936 7564 43988
rect 7616 43976 7622 43988
rect 10873 43979 10931 43985
rect 10873 43976 10885 43979
rect 7616 43948 10885 43976
rect 7616 43936 7622 43948
rect 10873 43945 10885 43948
rect 10919 43945 10931 43979
rect 10873 43939 10931 43945
rect 11146 43936 11152 43988
rect 11204 43936 11210 43988
rect 842 43868 848 43920
rect 900 43908 906 43920
rect 2498 43908 2504 43920
rect 900 43880 2504 43908
rect 900 43868 906 43880
rect 2498 43868 2504 43880
rect 2556 43868 2562 43920
rect 8941 43911 8999 43917
rect 8941 43877 8953 43911
rect 8987 43908 8999 43911
rect 11164 43908 11192 43936
rect 8987 43880 11192 43908
rect 8987 43877 8999 43880
rect 8941 43871 8999 43877
rect 4706 43840 4712 43852
rect 4172 43812 4712 43840
rect 4062 43772 4068 43784
rect 4023 43744 4068 43772
rect 4062 43732 4068 43744
rect 4120 43732 4126 43784
rect 4172 43781 4200 43812
rect 4706 43800 4712 43812
rect 4764 43800 4770 43852
rect 8202 43840 8208 43852
rect 5092 43812 8208 43840
rect 5092 43784 5120 43812
rect 8202 43800 8208 43812
rect 8260 43840 8266 43852
rect 11149 43843 11207 43849
rect 11149 43840 11161 43843
rect 8260 43812 9720 43840
rect 8260 43800 8266 43812
rect 4157 43775 4215 43781
rect 4157 43741 4169 43775
rect 4203 43741 4215 43775
rect 4157 43735 4215 43741
rect 4341 43775 4399 43781
rect 4341 43741 4353 43775
rect 4387 43772 4399 43775
rect 5074 43772 5080 43784
rect 4387 43744 5080 43772
rect 4387 43741 4399 43744
rect 4341 43735 4399 43741
rect 5074 43732 5080 43744
rect 5132 43732 5138 43784
rect 8021 43775 8079 43781
rect 8021 43741 8033 43775
rect 8067 43772 8079 43775
rect 8110 43772 8116 43784
rect 8067 43744 8116 43772
rect 8067 43741 8079 43744
rect 8021 43735 8079 43741
rect 8110 43732 8116 43744
rect 8168 43732 8174 43784
rect 9692 43781 9720 43812
rect 9968 43812 11161 43840
rect 9401 43775 9459 43781
rect 9401 43741 9413 43775
rect 9447 43741 9459 43775
rect 9401 43735 9459 43741
rect 9493 43775 9551 43781
rect 9493 43741 9505 43775
rect 9539 43741 9551 43775
rect 9493 43735 9551 43741
rect 9677 43775 9735 43781
rect 9677 43741 9689 43775
rect 9723 43741 9735 43775
rect 9677 43735 9735 43741
rect 1210 43664 1216 43716
rect 1268 43704 1274 43716
rect 4801 43707 4859 43713
rect 4801 43704 4813 43707
rect 1268 43676 4813 43704
rect 1268 43664 1274 43676
rect 4801 43673 4813 43676
rect 4847 43673 4859 43707
rect 4801 43667 4859 43673
rect 4706 43596 4712 43648
rect 4764 43636 4770 43648
rect 5350 43636 5356 43648
rect 4764 43608 5356 43636
rect 4764 43596 4770 43608
rect 5350 43596 5356 43608
rect 5408 43596 5414 43648
rect 7282 43596 7288 43648
rect 7340 43636 7346 43648
rect 7653 43639 7711 43645
rect 7653 43636 7665 43639
rect 7340 43608 7665 43636
rect 7340 43596 7346 43608
rect 7653 43605 7665 43608
rect 7699 43605 7711 43639
rect 7653 43599 7711 43605
rect 8113 43639 8171 43645
rect 8113 43605 8125 43639
rect 8159 43636 8171 43639
rect 8941 43639 8999 43645
rect 8941 43636 8953 43639
rect 8159 43608 8953 43636
rect 8159 43605 8171 43608
rect 8113 43599 8171 43605
rect 8941 43605 8953 43608
rect 8987 43605 8999 43639
rect 9416 43636 9444 43735
rect 9508 43704 9536 43735
rect 9968 43704 9996 43812
rect 11149 43809 11161 43812
rect 11195 43809 11207 43843
rect 11149 43803 11207 43809
rect 11425 43775 11483 43781
rect 11425 43741 11437 43775
rect 11471 43772 11483 43775
rect 11606 43772 11612 43784
rect 11471 43744 11612 43772
rect 11471 43741 11483 43744
rect 11425 43735 11483 43741
rect 11606 43732 11612 43744
rect 11664 43732 11670 43784
rect 10134 43704 10140 43716
rect 9508 43676 9996 43704
rect 10095 43676 10140 43704
rect 10134 43664 10140 43676
rect 10192 43664 10198 43716
rect 11149 43707 11207 43713
rect 11149 43673 11161 43707
rect 11195 43704 11207 43707
rect 11330 43704 11336 43716
rect 11195 43676 11336 43704
rect 11195 43673 11207 43676
rect 11149 43667 11207 43673
rect 11330 43664 11336 43676
rect 11388 43664 11394 43716
rect 9674 43636 9680 43648
rect 9416 43608 9680 43636
rect 8941 43599 8999 43605
rect 9674 43596 9680 43608
rect 9732 43636 9738 43648
rect 10410 43636 10416 43648
rect 9732 43608 10416 43636
rect 9732 43596 9738 43608
rect 10410 43596 10416 43608
rect 10468 43596 10474 43648
rect 10873 43639 10931 43645
rect 10873 43605 10885 43639
rect 10919 43636 10931 43639
rect 11606 43636 11612 43648
rect 10919 43608 11612 43636
rect 10919 43605 10931 43608
rect 10873 43599 10931 43605
rect 11606 43596 11612 43608
rect 11664 43596 11670 43648
rect 1104 43546 10856 43568
rect 1104 43494 4213 43546
rect 4265 43494 4277 43546
rect 4329 43494 4341 43546
rect 4393 43494 4405 43546
rect 4457 43494 4469 43546
rect 4521 43494 7477 43546
rect 7529 43494 7541 43546
rect 7593 43494 7605 43546
rect 7657 43494 7669 43546
rect 7721 43494 7733 43546
rect 7785 43494 10856 43546
rect 1104 43472 10856 43494
rect 1949 43435 2007 43441
rect 1949 43401 1961 43435
rect 1995 43432 2007 43435
rect 6914 43432 6920 43444
rect 1995 43404 6920 43432
rect 1995 43401 2007 43404
rect 1949 43395 2007 43401
rect 6914 43392 6920 43404
rect 6972 43392 6978 43444
rect 8294 43392 8300 43444
rect 8352 43432 8358 43444
rect 9309 43435 9367 43441
rect 9309 43432 9321 43435
rect 8352 43404 9321 43432
rect 8352 43392 8358 43404
rect 9309 43401 9321 43404
rect 9355 43401 9367 43435
rect 9309 43395 9367 43401
rect 9674 43392 9680 43444
rect 9732 43432 9738 43444
rect 9858 43432 9864 43444
rect 9732 43404 9864 43432
rect 9732 43392 9738 43404
rect 9858 43392 9864 43404
rect 9916 43392 9922 43444
rect 3602 43324 3608 43376
rect 3660 43364 3666 43376
rect 3970 43364 3976 43376
rect 3660 43336 3976 43364
rect 3660 43324 3666 43336
rect 3970 43324 3976 43336
rect 4028 43324 4034 43376
rect 5350 43324 5356 43376
rect 5408 43364 5414 43376
rect 6638 43364 6644 43376
rect 5408 43336 6644 43364
rect 5408 43324 5414 43336
rect 6638 43324 6644 43336
rect 6696 43324 6702 43376
rect 8570 43364 8576 43376
rect 6748 43336 8576 43364
rect 1854 43296 1860 43308
rect 1815 43268 1860 43296
rect 1854 43256 1860 43268
rect 1912 43256 1918 43308
rect 6362 43256 6368 43308
rect 6420 43296 6426 43308
rect 6748 43296 6776 43336
rect 8570 43324 8576 43336
rect 8628 43324 8634 43376
rect 6420 43268 6776 43296
rect 8389 43299 8447 43305
rect 6420 43256 6426 43268
rect 8389 43265 8401 43299
rect 8435 43265 8447 43299
rect 9122 43296 9128 43308
rect 9083 43268 9128 43296
rect 8389 43259 8447 43265
rect 8404 43228 8432 43259
rect 9122 43256 9128 43268
rect 9180 43256 9186 43308
rect 9858 43296 9864 43308
rect 9819 43268 9864 43296
rect 9858 43256 9864 43268
rect 9916 43256 9922 43308
rect 9950 43256 9956 43308
rect 10008 43296 10014 43308
rect 10686 43296 10692 43308
rect 10008 43268 10692 43296
rect 10008 43256 10014 43268
rect 10686 43256 10692 43268
rect 10744 43256 10750 43308
rect 10962 43228 10968 43240
rect 8404 43200 10968 43228
rect 10962 43188 10968 43200
rect 11020 43188 11026 43240
rect 11054 43188 11060 43240
rect 11112 43228 11118 43240
rect 11330 43228 11336 43240
rect 11112 43200 11336 43228
rect 11112 43188 11118 43200
rect 11330 43188 11336 43200
rect 11388 43188 11394 43240
rect 1118 43120 1124 43172
rect 1176 43160 1182 43172
rect 10134 43160 10140 43172
rect 1176 43132 10140 43160
rect 1176 43120 1182 43132
rect 10134 43120 10140 43132
rect 10192 43120 10198 43172
rect 8570 43092 8576 43104
rect 8531 43064 8576 43092
rect 8570 43052 8576 43064
rect 8628 43052 8634 43104
rect 9769 43095 9827 43101
rect 9769 43061 9781 43095
rect 9815 43092 9827 43095
rect 10045 43095 10103 43101
rect 10045 43092 10057 43095
rect 9815 43064 10057 43092
rect 9815 43061 9827 43064
rect 9769 43055 9827 43061
rect 10045 43061 10057 43064
rect 10091 43092 10103 43095
rect 11054 43092 11060 43104
rect 10091 43064 11060 43092
rect 10091 43061 10103 43064
rect 10045 43055 10103 43061
rect 11054 43052 11060 43064
rect 11112 43052 11118 43104
rect 1104 43002 10856 43024
rect 1104 42950 2582 43002
rect 2634 42950 2646 43002
rect 2698 42950 2710 43002
rect 2762 42950 2774 43002
rect 2826 42950 2838 43002
rect 2890 42950 5845 43002
rect 5897 42950 5909 43002
rect 5961 42950 5973 43002
rect 6025 42950 6037 43002
rect 6089 42950 6101 43002
rect 6153 42950 9109 43002
rect 9161 42950 9173 43002
rect 9225 42950 9237 43002
rect 9289 42950 9301 43002
rect 9353 42950 9365 43002
rect 9417 42950 10856 43002
rect 1104 42928 10856 42950
rect 4062 42848 4068 42900
rect 4120 42888 4126 42900
rect 4120 42860 6684 42888
rect 4120 42848 4126 42860
rect 6549 42823 6607 42829
rect 6549 42789 6561 42823
rect 6595 42789 6607 42823
rect 6656 42820 6684 42860
rect 6822 42848 6828 42900
rect 6880 42888 6886 42900
rect 10686 42888 10692 42900
rect 6880 42860 10692 42888
rect 6880 42848 6886 42860
rect 10686 42848 10692 42860
rect 10744 42848 10750 42900
rect 10134 42820 10140 42832
rect 6656 42792 10140 42820
rect 6549 42783 6607 42789
rect 6362 42752 6368 42764
rect 2746 42724 6368 42752
rect 1394 42684 1400 42696
rect 1355 42656 1400 42684
rect 1394 42644 1400 42656
rect 1452 42644 1458 42696
rect 1581 42551 1639 42557
rect 1581 42517 1593 42551
rect 1627 42548 1639 42551
rect 2746 42548 2774 42724
rect 6362 42712 6368 42724
rect 6420 42712 6426 42764
rect 6564 42752 6592 42783
rect 10134 42780 10140 42792
rect 10192 42780 10198 42832
rect 6822 42752 6828 42764
rect 6564 42724 6828 42752
rect 6822 42712 6828 42724
rect 6880 42712 6886 42764
rect 6914 42712 6920 42764
rect 6972 42752 6978 42764
rect 7101 42755 7159 42761
rect 7101 42752 7113 42755
rect 6972 42724 7113 42752
rect 6972 42712 6978 42724
rect 7101 42721 7113 42724
rect 7147 42752 7159 42755
rect 9953 42755 10011 42761
rect 7147 42724 9628 42752
rect 7147 42721 7159 42724
rect 7101 42715 7159 42721
rect 3602 42644 3608 42696
rect 3660 42684 3666 42696
rect 9475 42687 9533 42693
rect 9475 42684 9487 42687
rect 3660 42656 9487 42684
rect 3660 42644 3666 42656
rect 9475 42653 9487 42656
rect 9521 42653 9533 42687
rect 9600 42684 9628 42724
rect 9953 42721 9965 42755
rect 9999 42752 10011 42755
rect 9999 42724 10364 42752
rect 9999 42721 10011 42724
rect 9953 42715 10011 42721
rect 10045 42687 10103 42693
rect 10045 42684 10057 42687
rect 9600 42656 10057 42684
rect 9475 42647 9533 42653
rect 10045 42653 10057 42656
rect 10091 42653 10103 42687
rect 10045 42647 10103 42653
rect 3970 42576 3976 42628
rect 4028 42616 4034 42628
rect 6546 42616 6552 42628
rect 4028 42588 6552 42616
rect 4028 42576 4034 42588
rect 6546 42576 6552 42588
rect 6604 42576 6610 42628
rect 6825 42619 6883 42625
rect 6825 42585 6837 42619
rect 6871 42585 6883 42619
rect 6825 42579 6883 42585
rect 1627 42520 2774 42548
rect 1627 42517 1639 42520
rect 1581 42511 1639 42517
rect 3510 42508 3516 42560
rect 3568 42548 3574 42560
rect 6362 42548 6368 42560
rect 3568 42520 6368 42548
rect 3568 42508 3574 42520
rect 6362 42508 6368 42520
rect 6420 42548 6426 42560
rect 6840 42548 6868 42579
rect 8202 42576 8208 42628
rect 8260 42616 8266 42628
rect 8570 42616 8576 42628
rect 8260 42588 8576 42616
rect 8260 42576 8266 42588
rect 8570 42576 8576 42588
rect 8628 42576 8634 42628
rect 9125 42619 9183 42625
rect 9125 42585 9137 42619
rect 9171 42616 9183 42619
rect 9309 42619 9367 42625
rect 9309 42616 9321 42619
rect 9171 42588 9321 42616
rect 9171 42585 9183 42588
rect 9125 42579 9183 42585
rect 9309 42585 9321 42588
rect 9355 42616 9367 42619
rect 9950 42616 9956 42628
rect 9355 42588 9956 42616
rect 9355 42585 9367 42588
rect 9309 42579 9367 42585
rect 9950 42576 9956 42588
rect 10008 42576 10014 42628
rect 6420 42520 6868 42548
rect 6420 42508 6426 42520
rect 6914 42508 6920 42560
rect 6972 42548 6978 42560
rect 10336 42557 10364 42724
rect 11146 42712 11152 42764
rect 11204 42752 11210 42764
rect 11698 42752 11704 42764
rect 11204 42724 11704 42752
rect 11204 42712 11210 42724
rect 11698 42712 11704 42724
rect 11756 42712 11762 42764
rect 7009 42551 7067 42557
rect 7009 42548 7021 42551
rect 6972 42520 7021 42548
rect 6972 42508 6978 42520
rect 7009 42517 7021 42520
rect 7055 42517 7067 42551
rect 7009 42511 7067 42517
rect 10321 42551 10379 42557
rect 10321 42517 10333 42551
rect 10367 42548 10379 42551
rect 11698 42548 11704 42560
rect 10367 42520 11704 42548
rect 10367 42517 10379 42520
rect 10321 42511 10379 42517
rect 11698 42508 11704 42520
rect 11756 42508 11762 42560
rect 1104 42458 10856 42480
rect 1104 42406 4213 42458
rect 4265 42406 4277 42458
rect 4329 42406 4341 42458
rect 4393 42406 4405 42458
rect 4457 42406 4469 42458
rect 4521 42406 7477 42458
rect 7529 42406 7541 42458
rect 7593 42406 7605 42458
rect 7657 42406 7669 42458
rect 7721 42406 7733 42458
rect 7785 42406 10856 42458
rect 1104 42384 10856 42406
rect 1578 42344 1584 42356
rect 1539 42316 1584 42344
rect 1578 42304 1584 42316
rect 1636 42304 1642 42356
rect 5074 42236 5080 42288
rect 5132 42276 5138 42288
rect 5261 42279 5319 42285
rect 5261 42276 5273 42279
rect 5132 42248 5273 42276
rect 5132 42236 5138 42248
rect 5261 42245 5273 42248
rect 5307 42245 5319 42279
rect 5261 42239 5319 42245
rect 6362 42236 6368 42288
rect 6420 42276 6426 42288
rect 6546 42276 6552 42288
rect 6420 42248 6552 42276
rect 6420 42236 6426 42248
rect 6546 42236 6552 42248
rect 6604 42236 6610 42288
rect 6914 42236 6920 42288
rect 6972 42276 6978 42288
rect 11146 42276 11152 42288
rect 6972 42248 11152 42276
rect 6972 42236 6978 42248
rect 11146 42236 11152 42248
rect 11204 42236 11210 42288
rect 1394 42208 1400 42220
rect 1355 42180 1400 42208
rect 1394 42168 1400 42180
rect 1452 42168 1458 42220
rect 3234 42168 3240 42220
rect 3292 42208 3298 42220
rect 5353 42211 5411 42217
rect 5353 42208 5365 42211
rect 3292 42180 5365 42208
rect 3292 42168 3298 42180
rect 5353 42177 5365 42180
rect 5399 42208 5411 42211
rect 6086 42208 6092 42220
rect 5399 42180 6092 42208
rect 5399 42177 5411 42180
rect 5353 42171 5411 42177
rect 6086 42168 6092 42180
rect 6144 42168 6150 42220
rect 9122 42208 9128 42220
rect 9083 42180 9128 42208
rect 9122 42168 9128 42180
rect 9180 42168 9186 42220
rect 9950 42208 9956 42220
rect 9911 42180 9956 42208
rect 9950 42168 9956 42180
rect 10008 42168 10014 42220
rect 10134 42168 10140 42220
rect 10192 42168 10198 42220
rect 5166 42140 5172 42152
rect 5127 42112 5172 42140
rect 5166 42100 5172 42112
rect 5224 42100 5230 42152
rect 10152 42140 10180 42168
rect 8128 42112 10180 42140
rect 4801 42075 4859 42081
rect 4801 42041 4813 42075
rect 4847 42072 4859 42075
rect 8128 42072 8156 42112
rect 4847 42044 8156 42072
rect 4847 42041 4859 42044
rect 4801 42035 4859 42041
rect 8202 42032 8208 42084
rect 8260 42072 8266 42084
rect 10137 42075 10195 42081
rect 10137 42072 10149 42075
rect 8260 42044 10149 42072
rect 8260 42032 8266 42044
rect 10137 42041 10149 42044
rect 10183 42041 10195 42075
rect 10137 42035 10195 42041
rect 6362 41964 6368 42016
rect 6420 42004 6426 42016
rect 9309 42007 9367 42013
rect 9309 42004 9321 42007
rect 6420 41976 9321 42004
rect 6420 41964 6426 41976
rect 9309 41973 9321 41976
rect 9355 41973 9367 42007
rect 11241 42007 11299 42013
rect 11241 42004 11253 42007
rect 9309 41967 9367 41973
rect 10888 41976 11253 42004
rect 1104 41914 10856 41936
rect 1104 41862 2582 41914
rect 2634 41862 2646 41914
rect 2698 41862 2710 41914
rect 2762 41862 2774 41914
rect 2826 41862 2838 41914
rect 2890 41862 5845 41914
rect 5897 41862 5909 41914
rect 5961 41862 5973 41914
rect 6025 41862 6037 41914
rect 6089 41862 6101 41914
rect 6153 41862 9109 41914
rect 9161 41862 9173 41914
rect 9225 41862 9237 41914
rect 9289 41862 9301 41914
rect 9353 41862 9365 41914
rect 9417 41862 10856 41914
rect 1104 41840 10856 41862
rect 1581 41803 1639 41809
rect 1581 41769 1593 41803
rect 1627 41800 1639 41803
rect 2406 41800 2412 41812
rect 1627 41772 2412 41800
rect 1627 41769 1639 41772
rect 1581 41763 1639 41769
rect 2406 41760 2412 41772
rect 2464 41760 2470 41812
rect 934 41692 940 41744
rect 992 41732 998 41744
rect 6362 41732 6368 41744
rect 992 41704 6368 41732
rect 992 41692 998 41704
rect 6362 41692 6368 41704
rect 6420 41692 6426 41744
rect 8938 41692 8944 41744
rect 8996 41732 9002 41744
rect 9398 41732 9404 41744
rect 8996 41704 9404 41732
rect 8996 41692 9002 41704
rect 9398 41692 9404 41704
rect 9456 41692 9462 41744
rect 3510 41624 3516 41676
rect 3568 41664 3574 41676
rect 10134 41664 10140 41676
rect 3568 41636 10140 41664
rect 3568 41624 3574 41636
rect 10134 41624 10140 41636
rect 10192 41624 10198 41676
rect 1394 41596 1400 41608
rect 1355 41568 1400 41596
rect 1394 41556 1400 41568
rect 1452 41556 1458 41608
rect 3786 41556 3792 41608
rect 3844 41596 3850 41608
rect 9858 41596 9864 41608
rect 3844 41568 9864 41596
rect 3844 41556 3850 41568
rect 9858 41556 9864 41568
rect 9916 41556 9922 41608
rect 10686 41556 10692 41608
rect 10744 41596 10750 41608
rect 10888 41596 10916 41976
rect 11241 41973 11253 41976
rect 11287 41973 11299 42007
rect 11882 42004 11888 42016
rect 11241 41967 11299 41973
rect 11716 41976 11888 42004
rect 10965 41939 11023 41945
rect 10965 41905 10977 41939
rect 11011 41936 11023 41939
rect 11011 41908 11468 41936
rect 11011 41905 11023 41908
rect 10965 41899 11023 41905
rect 11330 41868 11336 41880
rect 10980 41840 11336 41868
rect 10980 41605 11008 41840
rect 11330 41828 11336 41840
rect 11388 41828 11394 41880
rect 11330 41692 11336 41744
rect 11388 41732 11394 41744
rect 11440 41732 11468 41908
rect 11517 41871 11575 41877
rect 11517 41837 11529 41871
rect 11563 41868 11575 41871
rect 11606 41868 11612 41880
rect 11563 41840 11612 41868
rect 11563 41837 11575 41840
rect 11517 41831 11575 41837
rect 11606 41828 11612 41840
rect 11664 41828 11670 41880
rect 11388 41704 11468 41732
rect 11517 41735 11575 41741
rect 11388 41692 11394 41704
rect 11517 41701 11529 41735
rect 11563 41732 11575 41735
rect 11716 41732 11744 41976
rect 11882 41964 11888 41976
rect 11940 41964 11946 42016
rect 11793 41939 11851 41945
rect 11793 41905 11805 41939
rect 11839 41905 11851 41939
rect 11793 41899 11851 41905
rect 11563 41704 11744 41732
rect 11563 41701 11575 41704
rect 11517 41695 11575 41701
rect 11808 41673 11836 41899
rect 11885 41803 11943 41809
rect 11885 41769 11897 41803
rect 11931 41769 11943 41803
rect 11885 41763 11943 41769
rect 11793 41667 11851 41673
rect 11793 41633 11805 41667
rect 11839 41633 11851 41667
rect 11793 41627 11851 41633
rect 10744 41568 10916 41596
rect 10965 41599 11023 41605
rect 10744 41556 10750 41568
rect 10965 41565 10977 41599
rect 11011 41565 11023 41599
rect 10965 41559 11023 41565
rect 11146 41556 11152 41608
rect 11204 41556 11210 41608
rect 3326 41488 3332 41540
rect 3384 41528 3390 41540
rect 5442 41528 5448 41540
rect 3384 41500 5448 41528
rect 3384 41488 3390 41500
rect 5442 41488 5448 41500
rect 5500 41488 5506 41540
rect 8570 41488 8576 41540
rect 8628 41528 8634 41540
rect 9950 41528 9956 41540
rect 8628 41500 8800 41528
rect 9911 41500 9956 41528
rect 8628 41488 8634 41500
rect 8772 41472 8800 41500
rect 9950 41488 9956 41500
rect 10008 41488 10014 41540
rect 10134 41488 10140 41540
rect 10192 41528 10198 41540
rect 10778 41528 10784 41540
rect 10192 41500 10784 41528
rect 10192 41488 10198 41500
rect 10778 41488 10784 41500
rect 10836 41488 10842 41540
rect 3786 41420 3792 41472
rect 3844 41460 3850 41472
rect 6914 41460 6920 41472
rect 3844 41432 6920 41460
rect 3844 41420 3850 41432
rect 6914 41420 6920 41432
rect 6972 41420 6978 41472
rect 8754 41420 8760 41472
rect 8812 41420 8818 41472
rect 10045 41463 10103 41469
rect 10045 41429 10057 41463
rect 10091 41460 10103 41463
rect 11164 41460 11192 41556
rect 11900 41540 11928 41763
rect 11882 41488 11888 41540
rect 11940 41488 11946 41540
rect 11238 41460 11244 41472
rect 10091 41432 11100 41460
rect 11164 41432 11244 41460
rect 10091 41429 10103 41432
rect 10045 41423 10103 41429
rect 11072 41392 11100 41432
rect 11238 41420 11244 41432
rect 11296 41420 11302 41472
rect 1104 41370 10856 41392
rect 1104 41318 4213 41370
rect 4265 41318 4277 41370
rect 4329 41318 4341 41370
rect 4393 41318 4405 41370
rect 4457 41318 4469 41370
rect 4521 41318 7477 41370
rect 7529 41318 7541 41370
rect 7593 41318 7605 41370
rect 7657 41318 7669 41370
rect 7721 41318 7733 41370
rect 7785 41318 10856 41370
rect 11072 41364 11744 41392
rect 1104 41296 10856 41318
rect 11054 41284 11060 41336
rect 11112 41324 11118 41336
rect 11146 41324 11152 41336
rect 11112 41296 11152 41324
rect 11112 41284 11118 41296
rect 11146 41284 11152 41296
rect 11204 41284 11210 41336
rect 2498 41216 2504 41268
rect 2556 41256 2562 41268
rect 5534 41256 5540 41268
rect 2556 41228 5540 41256
rect 2556 41216 2562 41228
rect 5534 41216 5540 41228
rect 5592 41216 5598 41268
rect 10873 41259 10931 41265
rect 10873 41256 10885 41259
rect 7484 41228 10885 41256
rect 7484 41200 7512 41228
rect 10873 41225 10885 41228
rect 10919 41225 10931 41259
rect 11425 41259 11483 41265
rect 11425 41256 11437 41259
rect 10873 41219 10931 41225
rect 11348 41228 11437 41256
rect 2041 41191 2099 41197
rect 2041 41157 2053 41191
rect 2087 41188 2099 41191
rect 2130 41188 2136 41200
rect 2087 41160 2136 41188
rect 2087 41157 2099 41160
rect 2041 41151 2099 41157
rect 2130 41148 2136 41160
rect 2188 41148 2194 41200
rect 7466 41148 7472 41200
rect 7524 41148 7530 41200
rect 11054 41148 11060 41200
rect 11112 41188 11118 41200
rect 11348 41188 11376 41228
rect 11425 41225 11437 41228
rect 11471 41225 11483 41259
rect 11425 41219 11483 41225
rect 11112 41160 11376 41188
rect 11112 41148 11118 41160
rect 1854 41120 1860 41132
rect 1815 41092 1860 41120
rect 1854 41080 1860 41092
rect 1912 41080 1918 41132
rect 6454 41080 6460 41132
rect 6512 41120 6518 41132
rect 6822 41120 6828 41132
rect 6512 41092 6828 41120
rect 6512 41080 6518 41092
rect 6822 41080 6828 41092
rect 6880 41080 6886 41132
rect 9950 41120 9956 41132
rect 9911 41092 9956 41120
rect 9950 41080 9956 41092
rect 10008 41080 10014 41132
rect 10962 41120 10968 41132
rect 10923 41092 10968 41120
rect 10962 41080 10968 41092
rect 11020 41080 11026 41132
rect 11716 41129 11744 41364
rect 11701 41123 11759 41129
rect 11701 41089 11713 41123
rect 11747 41089 11759 41123
rect 11701 41083 11759 41089
rect 1302 41012 1308 41064
rect 1360 41052 1366 41064
rect 9490 41052 9496 41064
rect 1360 41024 9496 41052
rect 1360 41012 1366 41024
rect 9490 41012 9496 41024
rect 9548 41012 9554 41064
rect 11057 41055 11115 41061
rect 11057 41021 11069 41055
rect 11103 41052 11115 41055
rect 11333 41055 11391 41061
rect 11333 41052 11345 41055
rect 11103 41024 11345 41052
rect 11103 41021 11115 41024
rect 11057 41015 11115 41021
rect 11333 41021 11345 41024
rect 11379 41021 11391 41055
rect 11333 41015 11391 41021
rect 11514 41012 11520 41064
rect 11572 41052 11578 41064
rect 11790 41052 11796 41064
rect 11572 41024 11796 41052
rect 11572 41012 11578 41024
rect 11790 41012 11796 41024
rect 11848 41012 11854 41064
rect 6822 40944 6828 40996
rect 6880 40984 6886 40996
rect 7190 40984 7196 40996
rect 6880 40956 7196 40984
rect 6880 40944 6886 40956
rect 7190 40944 7196 40956
rect 7248 40944 7254 40996
rect 8846 40944 8852 40996
rect 8904 40984 8910 40996
rect 9398 40984 9404 40996
rect 8904 40956 9404 40984
rect 8904 40944 8910 40956
rect 9398 40944 9404 40956
rect 9456 40944 9462 40996
rect 10137 40987 10195 40993
rect 10137 40953 10149 40987
rect 10183 40984 10195 40987
rect 10962 40984 10968 40996
rect 10183 40956 10968 40984
rect 10183 40953 10195 40956
rect 10137 40947 10195 40953
rect 10962 40944 10968 40956
rect 11020 40944 11026 40996
rect 6914 40876 6920 40928
rect 6972 40916 6978 40928
rect 7834 40916 7840 40928
rect 6972 40888 7840 40916
rect 6972 40876 6978 40888
rect 7834 40876 7840 40888
rect 7892 40876 7898 40928
rect 8570 40876 8576 40928
rect 8628 40916 8634 40928
rect 9490 40916 9496 40928
rect 8628 40888 9496 40916
rect 8628 40876 8634 40888
rect 9490 40876 9496 40888
rect 9548 40876 9554 40928
rect 10870 40876 10876 40928
rect 10928 40916 10934 40928
rect 11057 40919 11115 40925
rect 11057 40916 11069 40919
rect 10928 40888 11069 40916
rect 10928 40876 10934 40888
rect 11057 40885 11069 40888
rect 11103 40885 11115 40919
rect 11057 40879 11115 40885
rect 1104 40826 10856 40848
rect 1104 40774 2582 40826
rect 2634 40774 2646 40826
rect 2698 40774 2710 40826
rect 2762 40774 2774 40826
rect 2826 40774 2838 40826
rect 2890 40774 5845 40826
rect 5897 40774 5909 40826
rect 5961 40774 5973 40826
rect 6025 40774 6037 40826
rect 6089 40774 6101 40826
rect 6153 40774 9109 40826
rect 9161 40774 9173 40826
rect 9225 40774 9237 40826
rect 9289 40774 9301 40826
rect 9353 40774 9365 40826
rect 9417 40774 10856 40826
rect 1104 40752 10856 40774
rect 4982 40672 4988 40724
rect 5040 40712 5046 40724
rect 5442 40712 5448 40724
rect 5040 40684 5448 40712
rect 5040 40672 5046 40684
rect 5442 40672 5448 40684
rect 5500 40672 5506 40724
rect 7190 40672 7196 40724
rect 7248 40712 7254 40724
rect 7926 40712 7932 40724
rect 7248 40684 7932 40712
rect 7248 40672 7254 40684
rect 7926 40672 7932 40684
rect 7984 40672 7990 40724
rect 10870 40672 10876 40724
rect 10928 40712 10934 40724
rect 11149 40715 11207 40721
rect 11149 40712 11161 40715
rect 10928 40684 11161 40712
rect 10928 40672 10934 40684
rect 11149 40681 11161 40684
rect 11195 40681 11207 40715
rect 11149 40675 11207 40681
rect 2038 40644 2044 40656
rect 1999 40616 2044 40644
rect 2038 40604 2044 40616
rect 2096 40604 2102 40656
rect 9122 40604 9128 40656
rect 9180 40644 9186 40656
rect 11606 40644 11612 40656
rect 9180 40616 11612 40644
rect 9180 40604 9186 40616
rect 11606 40604 11612 40616
rect 11664 40604 11670 40656
rect 11885 40647 11943 40653
rect 11885 40613 11897 40647
rect 11931 40613 11943 40647
rect 11885 40607 11943 40613
rect 10134 40536 10140 40588
rect 10192 40536 10198 40588
rect 11057 40579 11115 40585
rect 11057 40545 11069 40579
rect 11103 40576 11115 40579
rect 11900 40576 11928 40607
rect 11103 40548 11928 40576
rect 11103 40545 11115 40548
rect 11057 40539 11115 40545
rect 5626 40468 5632 40520
rect 5684 40508 5690 40520
rect 9125 40511 9183 40517
rect 9125 40508 9137 40511
rect 5684 40480 9137 40508
rect 5684 40468 5690 40480
rect 9125 40477 9137 40480
rect 9171 40477 9183 40511
rect 9858 40508 9864 40520
rect 9819 40480 9864 40508
rect 9125 40471 9183 40477
rect 9858 40468 9864 40480
rect 9916 40468 9922 40520
rect 10152 40508 10180 40536
rect 11885 40511 11943 40517
rect 11885 40508 11897 40511
rect 10152 40480 11897 40508
rect 11885 40477 11897 40480
rect 11931 40477 11943 40511
rect 11885 40471 11943 40477
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 7466 40400 7472 40452
rect 7524 40400 7530 40452
rect 7926 40400 7932 40452
rect 7984 40440 7990 40452
rect 8202 40440 8208 40452
rect 7984 40412 8208 40440
rect 7984 40400 7990 40412
rect 8202 40400 8208 40412
rect 8260 40400 8266 40452
rect 10778 40440 10784 40452
rect 8496 40412 10784 40440
rect 5626 40332 5632 40384
rect 5684 40372 5690 40384
rect 7484 40372 7512 40400
rect 5684 40344 7512 40372
rect 5684 40332 5690 40344
rect 8018 40332 8024 40384
rect 8076 40372 8082 40384
rect 8496 40372 8524 40412
rect 10778 40400 10784 40412
rect 10836 40400 10842 40452
rect 9306 40372 9312 40384
rect 8076 40344 8524 40372
rect 9267 40344 9312 40372
rect 8076 40332 8082 40344
rect 9306 40332 9312 40344
rect 9364 40332 9370 40384
rect 10042 40372 10048 40384
rect 10003 40344 10048 40372
rect 10042 40332 10048 40344
rect 10100 40332 10106 40384
rect 10410 40332 10416 40384
rect 10468 40372 10474 40384
rect 11790 40372 11796 40384
rect 10468 40344 11796 40372
rect 10468 40332 10474 40344
rect 11790 40332 11796 40344
rect 11848 40332 11854 40384
rect 1104 40282 10856 40304
rect 1104 40230 4213 40282
rect 4265 40230 4277 40282
rect 4329 40230 4341 40282
rect 4393 40230 4405 40282
rect 4457 40230 4469 40282
rect 4521 40230 7477 40282
rect 7529 40230 7541 40282
rect 7593 40230 7605 40282
rect 7657 40230 7669 40282
rect 7721 40230 7733 40282
rect 7785 40230 10856 40282
rect 1104 40208 10856 40230
rect 9483 40171 9541 40177
rect 6380 40140 9444 40168
rect 1578 40060 1584 40112
rect 1636 40100 1642 40112
rect 3878 40100 3884 40112
rect 1636 40072 3884 40100
rect 1636 40060 1642 40072
rect 3878 40060 3884 40072
rect 3936 40060 3942 40112
rect 1670 40032 1676 40044
rect 1631 40004 1676 40032
rect 1670 39992 1676 40004
rect 1728 39992 1734 40044
rect 2038 39992 2044 40044
rect 2096 40032 2102 40044
rect 3326 40032 3332 40044
rect 2096 40004 3332 40032
rect 2096 39992 2102 40004
rect 3326 39992 3332 40004
rect 3384 39992 3390 40044
rect 1394 39964 1400 39976
rect 1355 39936 1400 39964
rect 1394 39924 1400 39936
rect 1452 39924 1458 39976
rect 6380 39964 6408 40140
rect 6454 40060 6460 40112
rect 6512 40100 6518 40112
rect 6825 40103 6883 40109
rect 6825 40100 6837 40103
rect 6512 40072 6837 40100
rect 6512 40060 6518 40072
rect 6825 40069 6837 40072
rect 6871 40069 6883 40103
rect 8570 40100 8576 40112
rect 6825 40063 6883 40069
rect 8496 40072 8576 40100
rect 8496 40041 8524 40072
rect 8570 40060 8576 40072
rect 8628 40060 8634 40112
rect 9416 40100 9444 40140
rect 9483 40137 9495 40171
rect 9529 40168 9541 40171
rect 9529 40140 11928 40168
rect 9529 40137 9541 40140
rect 9483 40131 9541 40137
rect 9858 40100 9864 40112
rect 9416 40072 9864 40100
rect 9858 40060 9864 40072
rect 9916 40060 9922 40112
rect 9953 40103 10011 40109
rect 9953 40069 9965 40103
rect 9999 40069 10011 40103
rect 9953 40063 10011 40069
rect 8481 40035 8539 40041
rect 8481 40001 8493 40035
rect 8527 40001 8539 40035
rect 8481 39995 8539 40001
rect 9125 40035 9183 40041
rect 9125 40001 9137 40035
rect 9171 40032 9183 40035
rect 9309 40035 9367 40041
rect 9309 40032 9321 40035
rect 9171 40004 9321 40032
rect 9171 40001 9183 40004
rect 9125 39995 9183 40001
rect 9309 40001 9321 40004
rect 9355 40032 9367 40035
rect 9968 40032 9996 40063
rect 10778 40060 10784 40112
rect 10836 40100 10842 40112
rect 11425 40103 11483 40109
rect 11425 40100 11437 40103
rect 10836 40072 11437 40100
rect 10836 40060 10842 40072
rect 11425 40069 11437 40072
rect 11471 40069 11483 40103
rect 11425 40063 11483 40069
rect 10134 40032 10140 40044
rect 9355 40004 10140 40032
rect 9355 40001 9367 40004
rect 9309 39995 9367 40001
rect 10134 39992 10140 40004
rect 10192 39992 10198 40044
rect 6380 39936 6500 39964
rect 6472 39905 6500 39936
rect 6546 39924 6552 39976
rect 6604 39964 6610 39976
rect 6917 39967 6975 39973
rect 6917 39964 6929 39967
rect 6604 39936 6929 39964
rect 6604 39924 6610 39936
rect 6917 39933 6929 39936
rect 6963 39933 6975 39967
rect 6917 39927 6975 39933
rect 7009 39967 7067 39973
rect 7009 39933 7021 39967
rect 7055 39933 7067 39967
rect 7009 39927 7067 39933
rect 9953 39967 10011 39973
rect 9953 39933 9965 39967
rect 9999 39933 10011 39967
rect 9953 39927 10011 39933
rect 10045 39967 10103 39973
rect 10045 39933 10057 39967
rect 10091 39964 10103 39967
rect 10410 39964 10416 39976
rect 10091 39936 10416 39964
rect 10091 39933 10103 39936
rect 10045 39927 10103 39933
rect 6457 39899 6515 39905
rect 6457 39865 6469 39899
rect 6503 39865 6515 39899
rect 7024 39896 7052 39927
rect 6457 39859 6515 39865
rect 6564 39868 7052 39896
rect 6564 39840 6592 39868
rect 7466 39856 7472 39908
rect 7524 39896 7530 39908
rect 9122 39896 9128 39908
rect 7524 39868 9128 39896
rect 7524 39856 7530 39868
rect 9122 39856 9128 39868
rect 9180 39856 9186 39908
rect 9968 39896 9996 39927
rect 10410 39924 10416 39936
rect 10468 39924 10474 39976
rect 9968 39868 10364 39896
rect 6546 39788 6552 39840
rect 6604 39788 6610 39840
rect 8662 39828 8668 39840
rect 8623 39800 8668 39828
rect 8662 39788 8668 39800
rect 8720 39788 8726 39840
rect 10336 39837 10364 39868
rect 10321 39831 10379 39837
rect 10321 39797 10333 39831
rect 10367 39828 10379 39831
rect 10686 39828 10692 39840
rect 10367 39800 10692 39828
rect 10367 39797 10379 39800
rect 10321 39791 10379 39797
rect 10686 39788 10692 39800
rect 10744 39788 10750 39840
rect 1104 39738 10856 39760
rect 1104 39686 2582 39738
rect 2634 39686 2646 39738
rect 2698 39686 2710 39738
rect 2762 39686 2774 39738
rect 2826 39686 2838 39738
rect 2890 39686 5845 39738
rect 5897 39686 5909 39738
rect 5961 39686 5973 39738
rect 6025 39686 6037 39738
rect 6089 39686 6101 39738
rect 6153 39686 9109 39738
rect 9161 39686 9173 39738
rect 9225 39686 9237 39738
rect 9289 39686 9301 39738
rect 9353 39686 9365 39738
rect 9417 39686 10856 39738
rect 1104 39664 10856 39686
rect 1857 39627 1915 39633
rect 1857 39593 1869 39627
rect 1903 39624 1915 39627
rect 2498 39624 2504 39636
rect 1903 39596 2504 39624
rect 1903 39593 1915 39596
rect 1857 39587 1915 39593
rect 2498 39584 2504 39596
rect 2556 39584 2562 39636
rect 2746 39596 5304 39624
rect 1670 39516 1676 39568
rect 1728 39556 1734 39568
rect 2746 39556 2774 39596
rect 1728 39528 2774 39556
rect 5276 39556 5304 39596
rect 7006 39584 7012 39636
rect 7064 39624 7070 39636
rect 9217 39627 9275 39633
rect 9217 39624 9229 39627
rect 7064 39596 9229 39624
rect 7064 39584 7070 39596
rect 9217 39593 9229 39596
rect 9263 39593 9275 39627
rect 9217 39587 9275 39593
rect 9950 39584 9956 39636
rect 10008 39584 10014 39636
rect 9968 39556 9996 39584
rect 11900 39568 11928 40140
rect 5276 39528 9996 39556
rect 1728 39516 1734 39528
rect 11882 39516 11888 39568
rect 11940 39516 11946 39568
rect 2314 39488 2320 39500
rect 2275 39460 2320 39488
rect 2314 39448 2320 39460
rect 2372 39448 2378 39500
rect 3234 39488 3240 39500
rect 2516 39460 3240 39488
rect 2516 39364 2544 39460
rect 3234 39448 3240 39460
rect 3292 39488 3298 39500
rect 5261 39491 5319 39497
rect 5261 39488 5273 39491
rect 3292 39460 5273 39488
rect 3292 39448 3298 39460
rect 5261 39457 5273 39460
rect 5307 39488 5319 39491
rect 6546 39488 6552 39500
rect 5307 39460 6552 39488
rect 5307 39457 5319 39460
rect 5261 39451 5319 39457
rect 6546 39448 6552 39460
rect 6604 39448 6610 39500
rect 9490 39448 9496 39500
rect 9548 39488 9554 39500
rect 9950 39488 9956 39500
rect 9548 39460 9956 39488
rect 9548 39448 9554 39460
rect 9950 39448 9956 39460
rect 10008 39448 10014 39500
rect 5166 39420 5172 39432
rect 5127 39392 5172 39420
rect 5166 39380 5172 39392
rect 5224 39380 5230 39432
rect 10134 39420 10140 39432
rect 9324 39392 10140 39420
rect 2409 39355 2467 39361
rect 2409 39321 2421 39355
rect 2455 39352 2467 39355
rect 2498 39352 2504 39364
rect 2455 39324 2504 39352
rect 2455 39321 2467 39324
rect 2409 39315 2467 39321
rect 2498 39312 2504 39324
rect 2556 39312 2562 39364
rect 9324 39352 9352 39392
rect 10134 39380 10140 39392
rect 10192 39380 10198 39432
rect 4724 39324 9352 39352
rect 2222 39244 2228 39296
rect 2280 39284 2286 39296
rect 4724 39293 4752 39324
rect 9398 39312 9404 39364
rect 9456 39352 9462 39364
rect 9493 39355 9551 39361
rect 9493 39352 9505 39355
rect 9456 39324 9505 39352
rect 9456 39312 9462 39324
rect 9493 39321 9505 39324
rect 9539 39321 9551 39355
rect 9769 39355 9827 39361
rect 9769 39352 9781 39355
rect 9493 39315 9551 39321
rect 9600 39324 9781 39352
rect 2317 39287 2375 39293
rect 2317 39284 2329 39287
rect 2280 39256 2329 39284
rect 2280 39244 2286 39256
rect 2317 39253 2329 39256
rect 2363 39253 2375 39287
rect 2317 39247 2375 39253
rect 4709 39287 4767 39293
rect 4709 39253 4721 39287
rect 4755 39253 4767 39287
rect 4709 39247 4767 39253
rect 4982 39244 4988 39296
rect 5040 39284 5046 39296
rect 5077 39287 5135 39293
rect 5077 39284 5089 39287
rect 5040 39256 5089 39284
rect 5040 39244 5046 39256
rect 5077 39253 5089 39256
rect 5123 39253 5135 39287
rect 5077 39247 5135 39253
rect 5166 39244 5172 39296
rect 5224 39284 5230 39296
rect 5626 39284 5632 39296
rect 5224 39256 5632 39284
rect 5224 39244 5230 39256
rect 5626 39244 5632 39256
rect 5684 39244 5690 39296
rect 6546 39244 6552 39296
rect 6604 39284 6610 39296
rect 9600 39284 9628 39324
rect 9769 39321 9781 39324
rect 9815 39352 9827 39355
rect 10410 39352 10416 39364
rect 9815 39324 10416 39352
rect 9815 39321 9827 39324
rect 9769 39315 9827 39321
rect 10410 39312 10416 39324
rect 10468 39312 10474 39364
rect 6604 39256 9628 39284
rect 9677 39287 9735 39293
rect 6604 39244 6610 39256
rect 9677 39253 9689 39287
rect 9723 39284 9735 39287
rect 9858 39284 9864 39296
rect 9723 39256 9864 39284
rect 9723 39253 9735 39256
rect 9677 39247 9735 39253
rect 9858 39244 9864 39256
rect 9916 39244 9922 39296
rect 1104 39194 10856 39216
rect 1104 39142 4213 39194
rect 4265 39142 4277 39194
rect 4329 39142 4341 39194
rect 4393 39142 4405 39194
rect 4457 39142 4469 39194
rect 4521 39142 7477 39194
rect 7529 39142 7541 39194
rect 7593 39142 7605 39194
rect 7657 39142 7669 39194
rect 7721 39142 7733 39194
rect 7785 39142 10856 39194
rect 1104 39120 10856 39142
rect 1578 39080 1584 39092
rect 1539 39052 1584 39080
rect 1578 39040 1584 39052
rect 1636 39040 1642 39092
rect 6822 38972 6828 39024
rect 6880 39012 6886 39024
rect 8018 39012 8024 39024
rect 6880 38984 8024 39012
rect 6880 38972 6886 38984
rect 8018 38972 8024 38984
rect 8076 38972 8082 39024
rect 8662 38972 8668 39024
rect 8720 39012 8726 39024
rect 9585 39015 9643 39021
rect 9585 39012 9597 39015
rect 8720 38984 9597 39012
rect 8720 38972 8726 38984
rect 9585 38981 9597 38984
rect 9631 38981 9643 39015
rect 9585 38975 9643 38981
rect 9677 39015 9735 39021
rect 9677 38981 9689 39015
rect 9723 39012 9735 39015
rect 10410 39012 10416 39024
rect 9723 38984 10416 39012
rect 9723 38981 9735 38984
rect 9677 38975 9735 38981
rect 1394 38944 1400 38956
rect 1355 38916 1400 38944
rect 1394 38904 1400 38916
rect 1452 38904 1458 38956
rect 3694 38904 3700 38956
rect 3752 38944 3758 38956
rect 8297 38947 8355 38953
rect 8297 38944 8309 38947
rect 3752 38916 8309 38944
rect 3752 38904 3758 38916
rect 8297 38913 8309 38916
rect 8343 38913 8355 38947
rect 8297 38907 8355 38913
rect 10060 38888 10088 38984
rect 10410 38972 10416 38984
rect 10468 38972 10474 39024
rect 9490 38876 9496 38888
rect 2746 38848 9496 38876
rect 1946 38768 1952 38820
rect 2004 38808 2010 38820
rect 2746 38808 2774 38848
rect 9490 38836 9496 38848
rect 9548 38836 9554 38888
rect 10042 38836 10048 38888
rect 10100 38836 10106 38888
rect 9122 38808 9128 38820
rect 2004 38780 2774 38808
rect 9083 38780 9128 38808
rect 2004 38768 2010 38780
rect 9122 38768 9128 38780
rect 9180 38768 9186 38820
rect 8110 38700 8116 38752
rect 8168 38740 8174 38752
rect 8481 38743 8539 38749
rect 8481 38740 8493 38743
rect 8168 38712 8493 38740
rect 8168 38700 8174 38712
rect 8481 38709 8493 38712
rect 8527 38709 8539 38743
rect 8481 38703 8539 38709
rect 1104 38650 10856 38672
rect 1104 38598 2582 38650
rect 2634 38598 2646 38650
rect 2698 38598 2710 38650
rect 2762 38598 2774 38650
rect 2826 38598 2838 38650
rect 2890 38598 5845 38650
rect 5897 38598 5909 38650
rect 5961 38598 5973 38650
rect 6025 38598 6037 38650
rect 6089 38598 6101 38650
rect 6153 38598 9109 38650
rect 9161 38598 9173 38650
rect 9225 38598 9237 38650
rect 9289 38598 9301 38650
rect 9353 38598 9365 38650
rect 9417 38598 10856 38650
rect 1104 38576 10856 38598
rect 566 38496 572 38548
rect 624 38536 630 38548
rect 1581 38539 1639 38545
rect 1581 38536 1593 38539
rect 624 38508 1593 38536
rect 624 38496 630 38508
rect 1581 38505 1593 38508
rect 1627 38505 1639 38539
rect 1581 38499 1639 38505
rect 7098 38496 7104 38548
rect 7156 38536 7162 38548
rect 9033 38539 9091 38545
rect 9033 38536 9045 38539
rect 7156 38508 9045 38536
rect 7156 38496 7162 38508
rect 9033 38505 9045 38508
rect 9079 38505 9091 38539
rect 9582 38536 9588 38548
rect 9033 38499 9091 38505
rect 9324 38508 9588 38536
rect 9324 38480 9352 38508
rect 9582 38496 9588 38508
rect 9640 38496 9646 38548
rect 9306 38428 9312 38480
rect 9364 38428 9370 38480
rect 6362 38360 6368 38412
rect 6420 38400 6426 38412
rect 7742 38400 7748 38412
rect 6420 38372 7748 38400
rect 6420 38360 6426 38372
rect 7742 38360 7748 38372
rect 7800 38400 7806 38412
rect 9401 38403 9459 38409
rect 9401 38400 9413 38403
rect 7800 38372 9413 38400
rect 7800 38360 7806 38372
rect 9401 38369 9413 38372
rect 9447 38369 9459 38403
rect 9401 38363 9459 38369
rect 9582 38360 9588 38412
rect 9640 38400 9646 38412
rect 10042 38400 10048 38412
rect 9640 38372 10048 38400
rect 9640 38360 9646 38372
rect 10042 38360 10048 38372
rect 10100 38360 10106 38412
rect 1394 38332 1400 38344
rect 1355 38304 1400 38332
rect 1394 38292 1400 38304
rect 1452 38292 1458 38344
rect 4798 38292 4804 38344
rect 4856 38332 4862 38344
rect 8113 38335 8171 38341
rect 8113 38332 8125 38335
rect 4856 38304 8125 38332
rect 4856 38292 4862 38304
rect 8113 38301 8125 38304
rect 8159 38301 8171 38335
rect 8113 38295 8171 38301
rect 8110 38156 8116 38208
rect 8168 38196 8174 38208
rect 8297 38199 8355 38205
rect 8297 38196 8309 38199
rect 8168 38168 8309 38196
rect 8168 38156 8174 38168
rect 8297 38165 8309 38168
rect 8343 38165 8355 38199
rect 8297 38159 8355 38165
rect 9214 38156 9220 38208
rect 9272 38196 9278 38208
rect 9493 38199 9551 38205
rect 9493 38196 9505 38199
rect 9272 38168 9505 38196
rect 9272 38156 9278 38168
rect 9493 38165 9505 38168
rect 9539 38165 9551 38199
rect 9493 38159 9551 38165
rect 1104 38106 10856 38128
rect 1104 38054 4213 38106
rect 4265 38054 4277 38106
rect 4329 38054 4341 38106
rect 4393 38054 4405 38106
rect 4457 38054 4469 38106
rect 4521 38054 7477 38106
rect 7529 38054 7541 38106
rect 7593 38054 7605 38106
rect 7657 38054 7669 38106
rect 7721 38054 7733 38106
rect 7785 38054 10856 38106
rect 1104 38032 10856 38054
rect 9033 37995 9091 38001
rect 9033 37961 9045 37995
rect 9079 37961 9091 37995
rect 9490 37992 9496 38004
rect 9451 37964 9496 37992
rect 9033 37955 9091 37961
rect 9048 37924 9076 37955
rect 9490 37952 9496 37964
rect 9548 37952 9554 38004
rect 9950 37924 9956 37936
rect 9048 37896 9956 37924
rect 9950 37884 9956 37896
rect 10008 37884 10014 37936
rect 1302 37816 1308 37868
rect 1360 37856 1366 37868
rect 1397 37859 1455 37865
rect 1397 37856 1409 37859
rect 1360 37828 1409 37856
rect 1360 37816 1366 37828
rect 1397 37825 1409 37828
rect 1443 37825 1455 37859
rect 1397 37819 1455 37825
rect 4890 37816 4896 37868
rect 4948 37856 4954 37868
rect 8297 37859 8355 37865
rect 8297 37856 8309 37859
rect 4948 37828 8309 37856
rect 4948 37816 4954 37828
rect 8297 37825 8309 37828
rect 8343 37825 8355 37859
rect 8297 37819 8355 37825
rect 8662 37816 8668 37868
rect 8720 37816 8726 37868
rect 9401 37859 9459 37865
rect 9401 37825 9413 37859
rect 9447 37825 9459 37859
rect 9401 37819 9459 37825
rect 8018 37748 8024 37800
rect 8076 37788 8082 37800
rect 8680 37788 8708 37816
rect 9416 37788 9444 37819
rect 9582 37788 9588 37800
rect 8076 37760 9444 37788
rect 9543 37760 9588 37788
rect 8076 37748 8082 37760
rect 9582 37748 9588 37760
rect 9640 37748 9646 37800
rect 1581 37723 1639 37729
rect 1581 37689 1593 37723
rect 1627 37720 1639 37723
rect 2682 37720 2688 37732
rect 1627 37692 2688 37720
rect 1627 37689 1639 37692
rect 1581 37683 1639 37689
rect 2682 37680 2688 37692
rect 2740 37680 2746 37732
rect 7742 37680 7748 37732
rect 7800 37720 7806 37732
rect 9122 37720 9128 37732
rect 7800 37692 9128 37720
rect 7800 37680 7806 37692
rect 9122 37680 9128 37692
rect 9180 37680 9186 37732
rect 8481 37655 8539 37661
rect 8481 37621 8493 37655
rect 8527 37652 8539 37655
rect 9582 37652 9588 37664
rect 8527 37624 9588 37652
rect 8527 37621 8539 37624
rect 8481 37615 8539 37621
rect 9582 37612 9588 37624
rect 9640 37612 9646 37664
rect 1104 37562 10856 37584
rect 1104 37510 2582 37562
rect 2634 37510 2646 37562
rect 2698 37510 2710 37562
rect 2762 37510 2774 37562
rect 2826 37510 2838 37562
rect 2890 37510 5845 37562
rect 5897 37510 5909 37562
rect 5961 37510 5973 37562
rect 6025 37510 6037 37562
rect 6089 37510 6101 37562
rect 6153 37510 9109 37562
rect 9161 37510 9173 37562
rect 9225 37510 9237 37562
rect 9289 37510 9301 37562
rect 9353 37510 9365 37562
rect 9417 37510 10856 37562
rect 1104 37488 10856 37510
rect 7742 37408 7748 37460
rect 7800 37448 7806 37460
rect 7800 37420 8294 37448
rect 7800 37408 7806 37420
rect 8110 37340 8116 37392
rect 8168 37340 8174 37392
rect 2409 37315 2467 37321
rect 2409 37281 2421 37315
rect 2455 37312 2467 37315
rect 2498 37312 2504 37324
rect 2455 37284 2504 37312
rect 2455 37281 2467 37284
rect 2409 37275 2467 37281
rect 2498 37272 2504 37284
rect 2556 37272 2562 37324
rect 8128 37312 8156 37340
rect 7944 37284 8156 37312
rect 8266 37312 8294 37420
rect 8386 37408 8392 37460
rect 8444 37448 8450 37460
rect 8570 37448 8576 37460
rect 8444 37420 8576 37448
rect 8444 37408 8450 37420
rect 8570 37408 8576 37420
rect 8628 37408 8634 37460
rect 8266 37284 9628 37312
rect 2133 37247 2191 37253
rect 2133 37213 2145 37247
rect 2179 37244 2191 37247
rect 2222 37244 2228 37256
rect 2179 37216 2228 37244
rect 2179 37213 2191 37216
rect 2133 37207 2191 37213
rect 2222 37204 2228 37216
rect 2280 37204 2286 37256
rect 6914 37204 6920 37256
rect 6972 37244 6978 37256
rect 7944 37244 7972 37284
rect 8110 37244 8116 37256
rect 6972 37216 7972 37244
rect 8071 37216 8116 37244
rect 6972 37204 6978 37216
rect 8110 37204 8116 37216
rect 8168 37204 8174 37256
rect 8294 37204 8300 37256
rect 8352 37244 8358 37256
rect 8478 37244 8484 37256
rect 8352 37216 8484 37244
rect 8352 37204 8358 37216
rect 8478 37204 8484 37216
rect 8536 37204 8542 37256
rect 9600 37253 9628 37284
rect 9674 37272 9680 37324
rect 9732 37312 9738 37324
rect 9732 37284 9777 37312
rect 9732 37272 9738 37284
rect 9585 37247 9643 37253
rect 9585 37213 9597 37247
rect 9631 37213 9643 37247
rect 9585 37207 9643 37213
rect 5626 37136 5632 37188
rect 5684 37176 5690 37188
rect 9493 37179 9551 37185
rect 9493 37176 9505 37179
rect 5684 37148 9505 37176
rect 5684 37136 5690 37148
rect 9493 37145 9505 37148
rect 9539 37176 9551 37179
rect 9539 37148 9674 37176
rect 9539 37145 9551 37148
rect 9493 37139 9551 37145
rect 1762 37108 1768 37120
rect 1723 37080 1768 37108
rect 1762 37068 1768 37080
rect 1820 37068 1826 37120
rect 2225 37111 2283 37117
rect 2225 37077 2237 37111
rect 2271 37108 2283 37111
rect 2314 37108 2320 37120
rect 2271 37080 2320 37108
rect 2271 37077 2283 37080
rect 2225 37071 2283 37077
rect 2314 37068 2320 37080
rect 2372 37068 2378 37120
rect 8110 37068 8116 37120
rect 8168 37108 8174 37120
rect 8297 37111 8355 37117
rect 8297 37108 8309 37111
rect 8168 37080 8309 37108
rect 8168 37068 8174 37080
rect 8297 37077 8309 37080
rect 8343 37077 8355 37111
rect 8297 37071 8355 37077
rect 8478 37068 8484 37120
rect 8536 37108 8542 37120
rect 9125 37111 9183 37117
rect 9125 37108 9137 37111
rect 8536 37080 9137 37108
rect 8536 37068 8542 37080
rect 9125 37077 9137 37080
rect 9171 37077 9183 37111
rect 9646 37108 9674 37148
rect 9858 37108 9864 37120
rect 9646 37080 9864 37108
rect 9125 37071 9183 37077
rect 9858 37068 9864 37080
rect 9916 37068 9922 37120
rect 11330 37068 11336 37120
rect 11388 37068 11394 37120
rect 11348 37040 11376 37068
rect 1104 37018 10856 37040
rect 1104 36966 4213 37018
rect 4265 36966 4277 37018
rect 4329 36966 4341 37018
rect 4393 36966 4405 37018
rect 4457 36966 4469 37018
rect 4521 36966 7477 37018
rect 7529 36966 7541 37018
rect 7593 36966 7605 37018
rect 7657 36966 7669 37018
rect 7721 36966 7733 37018
rect 7785 36966 10856 37018
rect 1104 36944 10856 36966
rect 11072 37012 11376 37040
rect 1762 36864 1768 36916
rect 1820 36904 1826 36916
rect 6270 36904 6276 36916
rect 1820 36876 6276 36904
rect 1820 36864 1826 36876
rect 6270 36864 6276 36876
rect 6328 36864 6334 36916
rect 8846 36864 8852 36916
rect 8904 36904 8910 36916
rect 9953 36907 10011 36913
rect 9953 36904 9965 36907
rect 8904 36876 9965 36904
rect 8904 36864 8910 36876
rect 9953 36873 9965 36876
rect 9999 36873 10011 36907
rect 9953 36867 10011 36873
rect 3418 36796 3424 36848
rect 3476 36836 3482 36848
rect 3476 36808 8708 36836
rect 3476 36796 3482 36808
rect 1578 36728 1584 36780
rect 1636 36768 1642 36780
rect 8680 36777 8708 36808
rect 9582 36796 9588 36848
rect 9640 36836 9646 36848
rect 9674 36836 9680 36848
rect 9640 36808 9680 36836
rect 9640 36796 9646 36808
rect 9674 36796 9680 36808
rect 9732 36836 9738 36848
rect 10045 36839 10103 36845
rect 10045 36836 10057 36839
rect 9732 36808 10057 36836
rect 9732 36796 9738 36808
rect 10045 36805 10057 36808
rect 10091 36805 10103 36839
rect 10045 36799 10103 36805
rect 7929 36771 7987 36777
rect 7929 36768 7941 36771
rect 1636 36740 7941 36768
rect 1636 36728 1642 36740
rect 7929 36737 7941 36740
rect 7975 36737 7987 36771
rect 7929 36731 7987 36737
rect 8665 36771 8723 36777
rect 8665 36737 8677 36771
rect 8711 36737 8723 36771
rect 8665 36731 8723 36737
rect 1394 36700 1400 36712
rect 1355 36672 1400 36700
rect 1394 36660 1400 36672
rect 1452 36660 1458 36712
rect 1673 36703 1731 36709
rect 1673 36669 1685 36703
rect 1719 36700 1731 36703
rect 6914 36700 6920 36712
rect 1719 36672 6920 36700
rect 1719 36669 1731 36672
rect 1673 36663 1731 36669
rect 6914 36660 6920 36672
rect 6972 36660 6978 36712
rect 9309 36703 9367 36709
rect 9309 36669 9321 36703
rect 9355 36700 9367 36703
rect 9953 36703 10011 36709
rect 9953 36700 9965 36703
rect 9355 36672 9965 36700
rect 9355 36669 9367 36672
rect 9309 36663 9367 36669
rect 9953 36669 9965 36672
rect 9999 36700 10011 36703
rect 11072 36700 11100 37012
rect 11330 36932 11336 36984
rect 11388 36972 11394 36984
rect 11606 36972 11612 36984
rect 11388 36944 11612 36972
rect 11388 36932 11394 36944
rect 11606 36932 11612 36944
rect 11664 36932 11670 36984
rect 11149 36839 11207 36845
rect 11149 36805 11161 36839
rect 11195 36836 11207 36839
rect 11606 36836 11612 36848
rect 11195 36808 11612 36836
rect 11195 36805 11207 36808
rect 11149 36799 11207 36805
rect 11606 36796 11612 36808
rect 11664 36796 11670 36848
rect 11149 36703 11207 36709
rect 11149 36700 11161 36703
rect 9999 36672 10364 36700
rect 11072 36672 11161 36700
rect 9999 36669 10011 36672
rect 9953 36663 10011 36669
rect 8110 36632 8116 36644
rect 8071 36604 8116 36632
rect 8110 36592 8116 36604
rect 8168 36592 8174 36644
rect 8846 36564 8852 36576
rect 8807 36536 8852 36564
rect 8846 36524 8852 36536
rect 8904 36524 8910 36576
rect 9490 36564 9496 36576
rect 9451 36536 9496 36564
rect 9490 36524 9496 36536
rect 9548 36524 9554 36576
rect 10336 36573 10364 36672
rect 11149 36669 11161 36672
rect 11195 36669 11207 36703
rect 11149 36663 11207 36669
rect 10321 36567 10379 36573
rect 10321 36533 10333 36567
rect 10367 36564 10379 36567
rect 11606 36564 11612 36576
rect 10367 36536 11612 36564
rect 10367 36533 10379 36536
rect 10321 36527 10379 36533
rect 11606 36524 11612 36536
rect 11664 36524 11670 36576
rect 1104 36474 10856 36496
rect 1104 36422 2582 36474
rect 2634 36422 2646 36474
rect 2698 36422 2710 36474
rect 2762 36422 2774 36474
rect 2826 36422 2838 36474
rect 2890 36422 5845 36474
rect 5897 36422 5909 36474
rect 5961 36422 5973 36474
rect 6025 36422 6037 36474
rect 6089 36422 6101 36474
rect 6153 36422 9109 36474
rect 9161 36422 9173 36474
rect 9225 36422 9237 36474
rect 9289 36422 9301 36474
rect 9353 36422 9365 36474
rect 9417 36422 10856 36474
rect 1104 36400 10856 36422
rect 1397 36363 1455 36369
rect 1397 36329 1409 36363
rect 1443 36360 1455 36363
rect 8018 36360 8024 36372
rect 1443 36332 8024 36360
rect 1443 36329 1455 36332
rect 1397 36323 1455 36329
rect 8018 36320 8024 36332
rect 8076 36320 8082 36372
rect 5534 36252 5540 36304
rect 5592 36292 5598 36304
rect 7834 36292 7840 36304
rect 5592 36264 7840 36292
rect 5592 36252 5598 36264
rect 7834 36252 7840 36264
rect 7892 36252 7898 36304
rect 8941 36295 8999 36301
rect 8941 36261 8953 36295
rect 8987 36292 8999 36295
rect 10226 36292 10232 36304
rect 8987 36264 10232 36292
rect 8987 36261 8999 36264
rect 8941 36255 8999 36261
rect 10226 36252 10232 36264
rect 10284 36252 10290 36304
rect 2314 36224 2320 36236
rect 2275 36196 2320 36224
rect 2314 36184 2320 36196
rect 2372 36184 2378 36236
rect 2498 36184 2504 36236
rect 2556 36224 2562 36236
rect 3050 36224 3056 36236
rect 2556 36196 2636 36224
rect 3011 36196 3056 36224
rect 2556 36184 2562 36196
rect 1578 36156 1584 36168
rect 1539 36128 1584 36156
rect 1578 36116 1584 36128
rect 1636 36116 1642 36168
rect 2406 36116 2412 36168
rect 2464 36156 2470 36168
rect 2608 36165 2636 36196
rect 3050 36184 3056 36196
rect 3108 36184 3114 36236
rect 6270 36184 6276 36236
rect 6328 36224 6334 36236
rect 8018 36224 8024 36236
rect 6328 36196 8024 36224
rect 6328 36184 6334 36196
rect 8018 36184 8024 36196
rect 8076 36184 8082 36236
rect 9398 36224 9404 36236
rect 9359 36196 9404 36224
rect 9398 36184 9404 36196
rect 9456 36184 9462 36236
rect 9582 36224 9588 36236
rect 9495 36196 9588 36224
rect 9582 36184 9588 36196
rect 9640 36224 9646 36236
rect 9674 36224 9680 36236
rect 9640 36196 9680 36224
rect 9640 36184 9646 36196
rect 9674 36184 9680 36196
rect 9732 36184 9738 36236
rect 2593 36159 2651 36165
rect 2464 36128 2509 36156
rect 2464 36116 2470 36128
rect 2593 36125 2605 36159
rect 2639 36125 2651 36159
rect 2593 36119 2651 36125
rect 1394 35980 1400 36032
rect 1452 36020 1458 36032
rect 8846 36020 8852 36032
rect 1452 35992 8852 36020
rect 1452 35980 1458 35992
rect 8846 35980 8852 35992
rect 8904 36020 8910 36032
rect 9309 36023 9367 36029
rect 9309 36020 9321 36023
rect 8904 35992 9321 36020
rect 8904 35980 8910 35992
rect 9309 35989 9321 35992
rect 9355 35989 9367 36023
rect 9309 35983 9367 35989
rect 1104 35930 10856 35952
rect 1104 35878 4213 35930
rect 4265 35878 4277 35930
rect 4329 35878 4341 35930
rect 4393 35878 4405 35930
rect 4457 35878 4469 35930
rect 4521 35878 7477 35930
rect 7529 35878 7541 35930
rect 7593 35878 7605 35930
rect 7657 35878 7669 35930
rect 7721 35878 7733 35930
rect 7785 35878 10856 35930
rect 1104 35856 10856 35878
rect 1397 35819 1455 35825
rect 1397 35785 1409 35819
rect 1443 35816 1455 35819
rect 5626 35816 5632 35828
rect 1443 35788 5632 35816
rect 1443 35785 1455 35788
rect 1397 35779 1455 35785
rect 5626 35776 5632 35788
rect 5684 35776 5690 35828
rect 9858 35776 9864 35828
rect 9916 35816 9922 35828
rect 10134 35816 10140 35828
rect 9916 35788 10140 35816
rect 9916 35776 9922 35788
rect 10134 35776 10140 35788
rect 10192 35776 10198 35828
rect 6362 35708 6368 35760
rect 6420 35748 6426 35760
rect 6420 35720 9904 35748
rect 6420 35708 6426 35720
rect 1578 35680 1584 35692
rect 1539 35652 1584 35680
rect 1578 35640 1584 35652
rect 1636 35640 1642 35692
rect 7190 35640 7196 35692
rect 7248 35680 7254 35692
rect 9876 35689 9904 35720
rect 9125 35683 9183 35689
rect 9125 35680 9137 35683
rect 7248 35652 9137 35680
rect 7248 35640 7254 35652
rect 9125 35649 9137 35652
rect 9171 35649 9183 35683
rect 9125 35643 9183 35649
rect 9861 35683 9919 35689
rect 9861 35649 9873 35683
rect 9907 35649 9919 35683
rect 9861 35643 9919 35649
rect 7190 35504 7196 35556
rect 7248 35544 7254 35556
rect 11149 35547 11207 35553
rect 11149 35544 11161 35547
rect 7248 35516 11161 35544
rect 7248 35504 7254 35516
rect 11149 35513 11161 35516
rect 11195 35513 11207 35547
rect 11149 35507 11207 35513
rect 8110 35436 8116 35488
rect 8168 35476 8174 35488
rect 9309 35479 9367 35485
rect 9309 35476 9321 35479
rect 8168 35448 9321 35476
rect 8168 35436 8174 35448
rect 9309 35445 9321 35448
rect 9355 35445 9367 35479
rect 9309 35439 9367 35445
rect 10045 35479 10103 35485
rect 10045 35445 10057 35479
rect 10091 35476 10103 35479
rect 10134 35476 10140 35488
rect 10091 35448 10140 35476
rect 10091 35445 10103 35448
rect 10045 35439 10103 35445
rect 10134 35436 10140 35448
rect 10192 35436 10198 35488
rect 1104 35386 10856 35408
rect 1104 35334 2582 35386
rect 2634 35334 2646 35386
rect 2698 35334 2710 35386
rect 2762 35334 2774 35386
rect 2826 35334 2838 35386
rect 2890 35334 5845 35386
rect 5897 35334 5909 35386
rect 5961 35334 5973 35386
rect 6025 35334 6037 35386
rect 6089 35334 6101 35386
rect 6153 35334 9109 35386
rect 9161 35334 9173 35386
rect 9225 35334 9237 35386
rect 9289 35334 9301 35386
rect 9353 35334 9365 35386
rect 9417 35334 10856 35386
rect 1104 35312 10856 35334
rect 1394 35272 1400 35284
rect 1355 35244 1400 35272
rect 1394 35232 1400 35244
rect 1452 35232 1458 35284
rect 8846 35232 8852 35284
rect 8904 35272 8910 35284
rect 9309 35275 9367 35281
rect 9309 35272 9321 35275
rect 8904 35244 9321 35272
rect 8904 35232 8910 35244
rect 9309 35241 9321 35244
rect 9355 35241 9367 35275
rect 9309 35235 9367 35241
rect 2314 35096 2320 35148
rect 2372 35136 2378 35148
rect 2501 35139 2559 35145
rect 2501 35136 2513 35139
rect 2372 35108 2513 35136
rect 2372 35096 2378 35108
rect 2501 35105 2513 35108
rect 2547 35105 2559 35139
rect 2501 35099 2559 35105
rect 2590 35096 2596 35148
rect 2648 35136 2654 35148
rect 2648 35108 2693 35136
rect 2648 35096 2654 35108
rect 9306 35096 9312 35148
rect 9364 35136 9370 35148
rect 10042 35136 10048 35148
rect 9364 35108 10048 35136
rect 9364 35096 9370 35108
rect 10042 35096 10048 35108
rect 10100 35096 10106 35148
rect 1578 35068 1584 35080
rect 1539 35040 1584 35068
rect 1578 35028 1584 35040
rect 1636 35028 1642 35080
rect 2038 35028 2044 35080
rect 2096 35068 2102 35080
rect 2406 35068 2412 35080
rect 2096 35040 2412 35068
rect 2096 35028 2102 35040
rect 2406 35028 2412 35040
rect 2464 35028 2470 35080
rect 4614 35028 4620 35080
rect 4672 35068 4678 35080
rect 9125 35071 9183 35077
rect 9125 35068 9137 35071
rect 4672 35040 9137 35068
rect 4672 35028 4678 35040
rect 9125 35037 9137 35040
rect 9171 35037 9183 35071
rect 9125 35031 9183 35037
rect 9766 35028 9772 35080
rect 9824 35068 9830 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9824 35040 9873 35068
rect 9824 35028 9830 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 8110 35000 8116 35012
rect 2056 34972 8116 35000
rect 2056 34941 2084 34972
rect 8110 34960 8116 34972
rect 8168 34960 8174 35012
rect 2041 34935 2099 34941
rect 2041 34901 2053 34935
rect 2087 34901 2099 34935
rect 10042 34932 10048 34944
rect 10003 34904 10048 34932
rect 2041 34895 2099 34901
rect 10042 34892 10048 34904
rect 10100 34892 10106 34944
rect 1104 34842 10856 34864
rect 1104 34790 4213 34842
rect 4265 34790 4277 34842
rect 4329 34790 4341 34842
rect 4393 34790 4405 34842
rect 4457 34790 4469 34842
rect 4521 34790 7477 34842
rect 7529 34790 7541 34842
rect 7593 34790 7605 34842
rect 7657 34790 7669 34842
rect 7721 34790 7733 34842
rect 7785 34790 10856 34842
rect 1104 34768 10856 34790
rect 4798 34688 4804 34740
rect 4856 34728 4862 34740
rect 9401 34731 9459 34737
rect 9401 34728 9413 34731
rect 4856 34700 9413 34728
rect 4856 34688 4862 34700
rect 9401 34697 9413 34700
rect 9447 34697 9459 34731
rect 9401 34691 9459 34697
rect 3142 34660 3148 34672
rect 3103 34632 3148 34660
rect 3142 34620 3148 34632
rect 3200 34620 3206 34672
rect 9306 34620 9312 34672
rect 9364 34660 9370 34672
rect 9861 34663 9919 34669
rect 9861 34660 9873 34663
rect 9364 34632 9873 34660
rect 9364 34620 9370 34632
rect 9861 34629 9873 34632
rect 9907 34629 9919 34663
rect 9861 34623 9919 34629
rect 2498 34592 2504 34604
rect 2459 34564 2504 34592
rect 2498 34552 2504 34564
rect 2556 34552 2562 34604
rect 2590 34552 2596 34604
rect 2648 34592 2654 34604
rect 2685 34595 2743 34601
rect 2685 34592 2697 34595
rect 2648 34564 2697 34592
rect 2648 34552 2654 34564
rect 2685 34561 2697 34564
rect 2731 34561 2743 34595
rect 2685 34555 2743 34561
rect 8662 34552 8668 34604
rect 8720 34592 8726 34604
rect 8846 34592 8852 34604
rect 8720 34564 8852 34592
rect 8720 34552 8726 34564
rect 8846 34552 8852 34564
rect 8904 34552 8910 34604
rect 9769 34595 9827 34601
rect 9769 34561 9781 34595
rect 9815 34561 9827 34595
rect 9769 34555 9827 34561
rect 658 34484 664 34536
rect 716 34524 722 34536
rect 2314 34524 2320 34536
rect 716 34496 2320 34524
rect 716 34484 722 34496
rect 2314 34484 2320 34496
rect 2372 34524 2378 34536
rect 2409 34527 2467 34533
rect 2409 34524 2421 34527
rect 2372 34496 2421 34524
rect 2372 34484 2378 34496
rect 2409 34493 2421 34496
rect 2455 34493 2467 34527
rect 2409 34487 2467 34493
rect 7834 34484 7840 34536
rect 7892 34524 7898 34536
rect 9217 34527 9275 34533
rect 9217 34524 9229 34527
rect 7892 34496 9229 34524
rect 7892 34484 7898 34496
rect 9217 34493 9229 34496
rect 9263 34524 9275 34527
rect 9784 34524 9812 34555
rect 9263 34496 9812 34524
rect 10045 34527 10103 34533
rect 9263 34493 9275 34496
rect 9217 34487 9275 34493
rect 10045 34493 10057 34527
rect 10091 34524 10103 34527
rect 10134 34524 10140 34536
rect 10091 34496 10140 34524
rect 10091 34493 10103 34496
rect 10045 34487 10103 34493
rect 9582 34416 9588 34468
rect 9640 34456 9646 34468
rect 10060 34456 10088 34487
rect 10134 34484 10140 34496
rect 10192 34484 10198 34536
rect 9640 34428 10088 34456
rect 9640 34416 9646 34428
rect 1104 34298 10856 34320
rect 1104 34246 2582 34298
rect 2634 34246 2646 34298
rect 2698 34246 2710 34298
rect 2762 34246 2774 34298
rect 2826 34246 2838 34298
rect 2890 34246 5845 34298
rect 5897 34246 5909 34298
rect 5961 34246 5973 34298
rect 6025 34246 6037 34298
rect 6089 34246 6101 34298
rect 6153 34246 9109 34298
rect 9161 34246 9173 34298
rect 9225 34246 9237 34298
rect 9289 34246 9301 34298
rect 9353 34246 9365 34298
rect 9417 34246 10856 34298
rect 1104 34224 10856 34246
rect 8018 34144 8024 34196
rect 8076 34184 8082 34196
rect 9766 34184 9772 34196
rect 8076 34156 9772 34184
rect 8076 34144 8082 34156
rect 9766 34144 9772 34156
rect 9824 34144 9830 34196
rect 1673 34051 1731 34057
rect 1673 34017 1685 34051
rect 1719 34048 1731 34051
rect 6454 34048 6460 34060
rect 1719 34020 6460 34048
rect 1719 34017 1731 34020
rect 1673 34011 1731 34017
rect 6454 34008 6460 34020
rect 6512 34008 6518 34060
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 7098 33940 7104 33992
rect 7156 33980 7162 33992
rect 9125 33983 9183 33989
rect 9125 33980 9137 33983
rect 7156 33952 9137 33980
rect 7156 33940 7162 33952
rect 9125 33949 9137 33952
rect 9171 33949 9183 33983
rect 9125 33943 9183 33949
rect 9861 33983 9919 33989
rect 9861 33949 9873 33983
rect 9907 33980 9919 33983
rect 10870 33980 10876 33992
rect 9907 33952 10876 33980
rect 9907 33949 9919 33952
rect 9861 33943 9919 33949
rect 10870 33940 10876 33952
rect 10928 33940 10934 33992
rect 9306 33844 9312 33856
rect 9267 33816 9312 33844
rect 9306 33804 9312 33816
rect 9364 33804 9370 33856
rect 10042 33844 10048 33856
rect 10003 33816 10048 33844
rect 10042 33804 10048 33816
rect 10100 33804 10106 33856
rect 1104 33754 10856 33776
rect 1104 33702 4213 33754
rect 4265 33702 4277 33754
rect 4329 33702 4341 33754
rect 4393 33702 4405 33754
rect 4457 33702 4469 33754
rect 4521 33702 7477 33754
rect 7529 33702 7541 33754
rect 7593 33702 7605 33754
rect 7657 33702 7669 33754
rect 7721 33702 7733 33754
rect 7785 33702 10856 33754
rect 1104 33680 10856 33702
rect 3418 33600 3424 33652
rect 3476 33640 3482 33652
rect 9401 33643 9459 33649
rect 9401 33640 9413 33643
rect 3476 33612 9413 33640
rect 3476 33600 3482 33612
rect 9401 33609 9413 33612
rect 9447 33609 9459 33643
rect 9401 33603 9459 33609
rect 9861 33643 9919 33649
rect 9861 33609 9873 33643
rect 9907 33640 9919 33643
rect 10778 33640 10784 33652
rect 9907 33612 10784 33640
rect 9907 33609 9919 33612
rect 9861 33603 9919 33609
rect 10778 33600 10784 33612
rect 10836 33600 10842 33652
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33504 1731 33507
rect 4982 33504 4988 33516
rect 1719 33476 4988 33504
rect 1719 33473 1731 33476
rect 1673 33467 1731 33473
rect 4982 33464 4988 33476
rect 5040 33464 5046 33516
rect 8662 33504 8668 33516
rect 8623 33476 8668 33504
rect 8662 33464 8668 33476
rect 8720 33464 8726 33516
rect 9125 33507 9183 33513
rect 9125 33473 9137 33507
rect 9171 33504 9183 33507
rect 9769 33507 9827 33513
rect 9769 33504 9781 33507
rect 9171 33476 9781 33504
rect 9171 33473 9183 33476
rect 9125 33467 9183 33473
rect 9769 33473 9781 33476
rect 9815 33473 9827 33507
rect 9769 33467 9827 33473
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 10045 33439 10103 33445
rect 10045 33405 10057 33439
rect 10091 33436 10103 33439
rect 10134 33436 10140 33448
rect 10091 33408 10140 33436
rect 10091 33405 10103 33408
rect 10045 33399 10103 33405
rect 10134 33396 10140 33408
rect 10192 33396 10198 33448
rect 8849 33371 8907 33377
rect 8849 33337 8861 33371
rect 8895 33368 8907 33371
rect 9582 33368 9588 33380
rect 8895 33340 9588 33368
rect 8895 33337 8907 33340
rect 8849 33331 8907 33337
rect 9582 33328 9588 33340
rect 9640 33328 9646 33380
rect 11149 33371 11207 33377
rect 11149 33337 11161 33371
rect 11195 33368 11207 33371
rect 11885 33371 11943 33377
rect 11885 33368 11897 33371
rect 11195 33340 11897 33368
rect 11195 33337 11207 33340
rect 11149 33331 11207 33337
rect 11885 33337 11897 33340
rect 11931 33337 11943 33371
rect 11885 33331 11943 33337
rect 8018 33260 8024 33312
rect 8076 33300 8082 33312
rect 9125 33303 9183 33309
rect 9125 33300 9137 33303
rect 8076 33272 9137 33300
rect 8076 33260 8082 33272
rect 9125 33269 9137 33272
rect 9171 33300 9183 33303
rect 9217 33303 9275 33309
rect 9217 33300 9229 33303
rect 9171 33272 9229 33300
rect 9171 33269 9183 33272
rect 9125 33263 9183 33269
rect 9217 33269 9229 33272
rect 9263 33269 9275 33303
rect 9217 33263 9275 33269
rect 10686 33260 10692 33312
rect 10744 33300 10750 33312
rect 11333 33303 11391 33309
rect 11333 33300 11345 33303
rect 10744 33272 11345 33300
rect 10744 33260 10750 33272
rect 11333 33269 11345 33272
rect 11379 33269 11391 33303
rect 11333 33263 11391 33269
rect 1104 33210 10856 33232
rect 1104 33158 2582 33210
rect 2634 33158 2646 33210
rect 2698 33158 2710 33210
rect 2762 33158 2774 33210
rect 2826 33158 2838 33210
rect 2890 33158 5845 33210
rect 5897 33158 5909 33210
rect 5961 33158 5973 33210
rect 6025 33158 6037 33210
rect 6089 33158 6101 33210
rect 6153 33158 9109 33210
rect 9161 33158 9173 33210
rect 9225 33158 9237 33210
rect 9289 33158 9301 33210
rect 9353 33158 9365 33210
rect 9417 33158 10856 33210
rect 1104 33136 10856 33158
rect 1397 33099 1455 33105
rect 1397 33065 1409 33099
rect 1443 33096 1455 33099
rect 2222 33096 2228 33108
rect 1443 33068 2228 33096
rect 1443 33065 1455 33068
rect 1397 33059 1455 33065
rect 2222 33056 2228 33068
rect 2280 33056 2286 33108
rect 8110 33056 8116 33108
rect 8168 33096 8174 33108
rect 8478 33096 8484 33108
rect 8168 33068 8484 33096
rect 8168 33056 8174 33068
rect 8478 33056 8484 33068
rect 8536 33056 8542 33108
rect 10413 33099 10471 33105
rect 10413 33065 10425 33099
rect 10459 33096 10471 33099
rect 10594 33096 10600 33108
rect 10459 33068 10600 33096
rect 10459 33065 10471 33068
rect 10413 33059 10471 33065
rect 10594 33056 10600 33068
rect 10652 33056 10658 33108
rect 4890 32988 4896 33040
rect 4948 33028 4954 33040
rect 9401 33031 9459 33037
rect 9401 33028 9413 33031
rect 4948 33000 9413 33028
rect 4948 32988 4954 33000
rect 9401 32997 9413 33000
rect 9447 32997 9459 33031
rect 9401 32991 9459 32997
rect 9674 32988 9680 33040
rect 9732 33028 9738 33040
rect 9858 33028 9864 33040
rect 9732 33000 9864 33028
rect 9732 32988 9738 33000
rect 9858 32988 9864 33000
rect 9916 32988 9922 33040
rect 11330 33028 11336 33040
rect 9968 33000 11336 33028
rect 2498 32920 2504 32972
rect 2556 32960 2562 32972
rect 2685 32963 2743 32969
rect 2685 32960 2697 32963
rect 2556 32932 2697 32960
rect 2556 32920 2562 32932
rect 2685 32929 2697 32932
rect 2731 32929 2743 32963
rect 2685 32923 2743 32929
rect 8110 32920 8116 32972
rect 8168 32960 8174 32972
rect 8846 32960 8852 32972
rect 8168 32932 8852 32960
rect 8168 32920 8174 32932
rect 8846 32920 8852 32932
rect 8904 32920 8910 32972
rect 1578 32892 1584 32904
rect 1539 32864 1584 32892
rect 1578 32852 1584 32864
rect 1636 32852 1642 32904
rect 2314 32852 2320 32904
rect 2372 32892 2378 32904
rect 2593 32895 2651 32901
rect 2593 32892 2605 32895
rect 2372 32864 2605 32892
rect 2372 32852 2378 32864
rect 2593 32861 2605 32864
rect 2639 32861 2651 32895
rect 2593 32855 2651 32861
rect 7006 32852 7012 32904
rect 7064 32892 7070 32904
rect 9033 32895 9091 32901
rect 9033 32892 9045 32895
rect 7064 32864 9045 32892
rect 7064 32852 7070 32864
rect 9033 32861 9045 32864
rect 9079 32861 9091 32895
rect 9033 32855 9091 32861
rect 9861 32895 9919 32901
rect 9861 32861 9873 32895
rect 9907 32892 9919 32895
rect 9968 32892 9996 33000
rect 11330 32988 11336 33000
rect 11388 32988 11394 33040
rect 10045 32963 10103 32969
rect 10045 32929 10057 32963
rect 10091 32960 10103 32963
rect 10134 32960 10140 32972
rect 10091 32932 10140 32960
rect 10091 32929 10103 32932
rect 10045 32923 10103 32929
rect 9907 32864 9996 32892
rect 9907 32861 9919 32864
rect 9861 32855 9919 32861
rect 7098 32784 7104 32836
rect 7156 32824 7162 32836
rect 9490 32824 9496 32836
rect 7156 32796 9496 32824
rect 7156 32784 7162 32796
rect 9490 32784 9496 32796
rect 9548 32784 9554 32836
rect 10060 32824 10088 32923
rect 10134 32920 10140 32932
rect 10192 32920 10198 32972
rect 10594 32920 10600 32972
rect 10652 32960 10658 32972
rect 11514 32960 11520 32972
rect 10652 32932 11520 32960
rect 10652 32920 10658 32932
rect 11514 32920 11520 32932
rect 11572 32920 11578 32972
rect 10229 32895 10287 32901
rect 10229 32861 10241 32895
rect 10275 32892 10287 32895
rect 11425 32895 11483 32901
rect 11425 32892 11437 32895
rect 10275 32864 11437 32892
rect 10275 32861 10287 32864
rect 10229 32855 10287 32861
rect 11425 32861 11437 32864
rect 11471 32861 11483 32895
rect 11425 32855 11483 32861
rect 11333 32827 11391 32833
rect 11333 32824 11345 32827
rect 10060 32796 11345 32824
rect 11333 32793 11345 32796
rect 11379 32793 11391 32827
rect 11333 32787 11391 32793
rect 2130 32756 2136 32768
rect 2091 32728 2136 32756
rect 2130 32716 2136 32728
rect 2188 32716 2194 32768
rect 2498 32756 2504 32768
rect 2459 32728 2504 32756
rect 2498 32716 2504 32728
rect 2556 32716 2562 32768
rect 9214 32756 9220 32768
rect 9175 32728 9220 32756
rect 9214 32716 9220 32728
rect 9272 32716 9278 32768
rect 9398 32716 9404 32768
rect 9456 32756 9462 32768
rect 9769 32759 9827 32765
rect 9769 32756 9781 32759
rect 9456 32728 9781 32756
rect 9456 32716 9462 32728
rect 9769 32725 9781 32728
rect 9815 32725 9827 32759
rect 9769 32719 9827 32725
rect 11425 32759 11483 32765
rect 11425 32725 11437 32759
rect 11471 32756 11483 32759
rect 11698 32756 11704 32768
rect 11471 32728 11704 32756
rect 11471 32725 11483 32728
rect 11425 32719 11483 32725
rect 11698 32716 11704 32728
rect 11756 32716 11762 32768
rect 11057 32691 11115 32697
rect 1104 32666 10856 32688
rect 1104 32614 4213 32666
rect 4265 32614 4277 32666
rect 4329 32614 4341 32666
rect 4393 32614 4405 32666
rect 4457 32614 4469 32666
rect 4521 32614 7477 32666
rect 7529 32614 7541 32666
rect 7593 32614 7605 32666
rect 7657 32614 7669 32666
rect 7721 32614 7733 32666
rect 7785 32614 10856 32666
rect 11057 32657 11069 32691
rect 11103 32688 11115 32691
rect 11330 32688 11336 32700
rect 11103 32660 11336 32688
rect 11103 32657 11115 32660
rect 11057 32651 11115 32657
rect 11330 32648 11336 32660
rect 11388 32648 11394 32700
rect 11882 32648 11888 32700
rect 11940 32688 11946 32700
rect 11940 32660 11985 32688
rect 11940 32648 11946 32660
rect 1104 32592 10856 32614
rect 1397 32555 1455 32561
rect 1397 32521 1409 32555
rect 1443 32552 1455 32555
rect 2038 32552 2044 32564
rect 1443 32524 2044 32552
rect 1443 32521 1455 32524
rect 1397 32515 1455 32521
rect 2038 32512 2044 32524
rect 2096 32512 2102 32564
rect 2130 32512 2136 32564
rect 2188 32552 2194 32564
rect 10042 32552 10048 32564
rect 2188 32524 10048 32552
rect 2188 32512 2194 32524
rect 10042 32512 10048 32524
rect 10100 32512 10106 32564
rect 10134 32444 10140 32496
rect 10192 32484 10198 32496
rect 11054 32484 11060 32496
rect 10192 32456 11060 32484
rect 10192 32444 10198 32456
rect 11054 32444 11060 32456
rect 11112 32444 11118 32496
rect 1578 32416 1584 32428
rect 1539 32388 1584 32416
rect 1578 32376 1584 32388
rect 1636 32376 1642 32428
rect 5442 32376 5448 32428
rect 5500 32416 5506 32428
rect 8665 32419 8723 32425
rect 8665 32416 8677 32419
rect 5500 32388 8677 32416
rect 5500 32376 5506 32388
rect 8665 32385 8677 32388
rect 8711 32385 8723 32419
rect 8665 32379 8723 32385
rect 11422 32376 11428 32428
rect 11480 32416 11486 32428
rect 11480 32388 11836 32416
rect 11480 32376 11486 32388
rect 9309 32351 9367 32357
rect 9309 32317 9321 32351
rect 9355 32348 9367 32351
rect 9398 32348 9404 32360
rect 9355 32320 9404 32348
rect 9355 32317 9367 32320
rect 9309 32311 9367 32317
rect 9398 32308 9404 32320
rect 9456 32348 9462 32360
rect 9456 32320 9674 32348
rect 9456 32308 9462 32320
rect 5166 32240 5172 32292
rect 5224 32280 5230 32292
rect 5442 32280 5448 32292
rect 5224 32252 5448 32280
rect 5224 32240 5230 32252
rect 5442 32240 5448 32252
rect 5500 32240 5506 32292
rect 9646 32280 9674 32320
rect 10229 32283 10287 32289
rect 10229 32280 10241 32283
rect 9646 32252 10241 32280
rect 10229 32249 10241 32252
rect 10275 32249 10287 32283
rect 10229 32243 10287 32249
rect 11146 32240 11152 32292
rect 11204 32240 11210 32292
rect 8846 32212 8852 32224
rect 8807 32184 8852 32212
rect 8846 32172 8852 32184
rect 8904 32172 8910 32224
rect 11057 32147 11115 32153
rect 1104 32122 10856 32144
rect 1104 32070 2582 32122
rect 2634 32070 2646 32122
rect 2698 32070 2710 32122
rect 2762 32070 2774 32122
rect 2826 32070 2838 32122
rect 2890 32070 5845 32122
rect 5897 32070 5909 32122
rect 5961 32070 5973 32122
rect 6025 32070 6037 32122
rect 6089 32070 6101 32122
rect 6153 32070 9109 32122
rect 9161 32070 9173 32122
rect 9225 32070 9237 32122
rect 9289 32070 9301 32122
rect 9353 32070 9365 32122
rect 9417 32070 10856 32122
rect 11057 32113 11069 32147
rect 11103 32113 11115 32147
rect 11057 32107 11115 32113
rect 1104 32048 10856 32070
rect 1397 32011 1455 32017
rect 1397 31977 1409 32011
rect 1443 32008 1455 32011
rect 2498 32008 2504 32020
rect 1443 31980 2504 32008
rect 1443 31977 1455 31980
rect 1397 31971 1455 31977
rect 2498 31968 2504 31980
rect 2556 31968 2562 32020
rect 10778 31968 10784 32020
rect 10836 32008 10842 32020
rect 11072 32017 11100 32107
rect 10873 32011 10931 32017
rect 10873 32008 10885 32011
rect 10836 31980 10885 32008
rect 10836 31968 10842 31980
rect 10873 31977 10885 31980
rect 10919 31977 10931 32011
rect 10873 31971 10931 31977
rect 11057 32011 11115 32017
rect 11057 31977 11069 32011
rect 11103 31977 11115 32011
rect 11057 31971 11115 31977
rect 11164 31949 11192 32240
rect 11808 32088 11836 32388
rect 11790 32036 11796 32088
rect 11848 32036 11854 32088
rect 11238 31968 11244 32020
rect 11296 31968 11302 32020
rect 11330 31968 11336 32020
rect 11388 31968 11394 32020
rect 11149 31943 11207 31949
rect 11149 31909 11161 31943
rect 11195 31909 11207 31943
rect 11149 31903 11207 31909
rect 6178 31832 6184 31884
rect 6236 31872 6242 31884
rect 6236 31844 10916 31872
rect 6236 31832 6242 31844
rect 10888 31816 10916 31844
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 9309 31807 9367 31813
rect 9309 31773 9321 31807
rect 9355 31804 9367 31807
rect 10229 31807 10287 31813
rect 10229 31804 10241 31807
rect 9355 31776 10241 31804
rect 9355 31773 9367 31776
rect 9309 31767 9367 31773
rect 10229 31773 10241 31776
rect 10275 31804 10287 31807
rect 10594 31804 10600 31816
rect 10275 31776 10600 31804
rect 10275 31773 10287 31776
rect 10229 31767 10287 31773
rect 10594 31764 10600 31776
rect 10652 31764 10658 31816
rect 10870 31764 10876 31816
rect 10928 31764 10934 31816
rect 9950 31696 9956 31748
rect 10008 31736 10014 31748
rect 10134 31736 10140 31748
rect 10008 31708 10140 31736
rect 10008 31696 10014 31708
rect 10134 31696 10140 31708
rect 10192 31696 10198 31748
rect 11256 31736 11284 31968
rect 11348 31816 11376 31968
rect 11606 31900 11612 31952
rect 11664 31940 11670 31952
rect 11701 31943 11759 31949
rect 11701 31940 11713 31943
rect 11664 31912 11713 31940
rect 11664 31900 11670 31912
rect 11701 31909 11713 31912
rect 11747 31909 11759 31943
rect 11701 31903 11759 31909
rect 11330 31764 11336 31816
rect 11388 31764 11394 31816
rect 11701 31807 11759 31813
rect 11701 31773 11713 31807
rect 11747 31804 11759 31807
rect 11882 31804 11888 31816
rect 11747 31776 11888 31804
rect 11747 31773 11759 31776
rect 11701 31767 11759 31773
rect 11882 31764 11888 31776
rect 11940 31764 11946 31816
rect 11072 31708 11284 31736
rect 1104 31578 10856 31600
rect 1104 31526 4213 31578
rect 4265 31526 4277 31578
rect 4329 31526 4341 31578
rect 4393 31526 4405 31578
rect 4457 31526 4469 31578
rect 4521 31526 7477 31578
rect 7529 31526 7541 31578
rect 7593 31526 7605 31578
rect 7657 31526 7669 31578
rect 7721 31526 7733 31578
rect 7785 31526 10856 31578
rect 1104 31504 10856 31526
rect 9861 31467 9919 31473
rect 9861 31433 9873 31467
rect 9907 31464 9919 31467
rect 9950 31464 9956 31476
rect 9907 31436 9956 31464
rect 9907 31433 9919 31436
rect 9861 31427 9919 31433
rect 9950 31424 9956 31436
rect 10008 31424 10014 31476
rect 10686 31464 10692 31476
rect 10269 31436 10692 31464
rect 10269 31337 10297 31436
rect 10686 31424 10692 31436
rect 10744 31424 10750 31476
rect 9769 31331 9827 31337
rect 9769 31297 9781 31331
rect 9815 31297 9827 31331
rect 9769 31291 9827 31297
rect 10254 31331 10312 31337
rect 10254 31297 10266 31331
rect 10300 31297 10312 31331
rect 10254 31291 10312 31297
rect 9784 31192 9812 31291
rect 10042 31260 10048 31272
rect 10003 31232 10048 31260
rect 10042 31220 10048 31232
rect 10100 31220 10106 31272
rect 10134 31220 10140 31272
rect 10192 31260 10198 31272
rect 10410 31260 10416 31272
rect 10192 31232 10416 31260
rect 10192 31220 10198 31232
rect 10410 31220 10416 31232
rect 10468 31220 10474 31272
rect 10962 31220 10968 31272
rect 11020 31260 11026 31272
rect 11072 31260 11100 31708
rect 11793 31671 11851 31677
rect 11793 31668 11805 31671
rect 11624 31640 11805 31668
rect 11149 31603 11207 31609
rect 11149 31569 11161 31603
rect 11195 31600 11207 31603
rect 11422 31600 11428 31612
rect 11195 31572 11428 31600
rect 11195 31569 11207 31572
rect 11149 31563 11207 31569
rect 11422 31560 11428 31572
rect 11480 31560 11486 31612
rect 11514 31492 11520 31544
rect 11572 31532 11578 31544
rect 11624 31532 11652 31640
rect 11793 31637 11805 31640
rect 11839 31637 11851 31671
rect 11793 31631 11851 31637
rect 11698 31560 11704 31612
rect 11756 31600 11762 31612
rect 11756 31572 11836 31600
rect 11756 31560 11762 31572
rect 11572 31504 11652 31532
rect 11572 31492 11578 31504
rect 11808 31337 11836 31572
rect 11793 31331 11851 31337
rect 11793 31297 11805 31331
rect 11839 31297 11851 31331
rect 11793 31291 11851 31297
rect 11885 31331 11943 31337
rect 11885 31297 11897 31331
rect 11931 31297 11943 31331
rect 11885 31291 11943 31297
rect 11020 31232 11100 31260
rect 11020 31220 11026 31232
rect 11606 31220 11612 31272
rect 11664 31260 11670 31272
rect 11900 31260 11928 31291
rect 11664 31232 11928 31260
rect 11664 31220 11670 31232
rect 10686 31192 10692 31204
rect 9784 31164 10692 31192
rect 10686 31152 10692 31164
rect 10744 31152 10750 31204
rect 8846 31084 8852 31136
rect 8904 31124 8910 31136
rect 9401 31127 9459 31133
rect 9401 31124 9413 31127
rect 8904 31096 9413 31124
rect 8904 31084 8910 31096
rect 9401 31093 9413 31096
rect 9447 31093 9459 31127
rect 10410 31124 10416 31136
rect 10371 31096 10416 31124
rect 9401 31087 9459 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 1104 31034 10856 31056
rect 1104 30982 2582 31034
rect 2634 30982 2646 31034
rect 2698 30982 2710 31034
rect 2762 30982 2774 31034
rect 2826 30982 2838 31034
rect 2890 30982 5845 31034
rect 5897 30982 5909 31034
rect 5961 30982 5973 31034
rect 6025 30982 6037 31034
rect 6089 30982 6101 31034
rect 6153 30982 9109 31034
rect 9161 30982 9173 31034
rect 9225 30982 9237 31034
rect 9289 30982 9301 31034
rect 9353 30982 9365 31034
rect 9417 30982 10856 31034
rect 1104 30960 10856 30982
rect 11333 30923 11391 30929
rect 11333 30889 11345 30923
rect 11379 30889 11391 30923
rect 11333 30883 11391 30889
rect 11348 30852 11376 30883
rect 10336 30824 11376 30852
rect 10134 30784 10140 30796
rect 1412 30756 10140 30784
rect 1412 30725 1440 30756
rect 10134 30744 10140 30756
rect 10192 30744 10198 30796
rect 1397 30719 1455 30725
rect 1397 30685 1409 30719
rect 1443 30685 1455 30719
rect 1397 30679 1455 30685
rect 7374 30676 7380 30728
rect 7432 30716 7438 30728
rect 9861 30719 9919 30725
rect 9861 30716 9873 30719
rect 7432 30688 9873 30716
rect 7432 30676 7438 30688
rect 9861 30685 9873 30688
rect 9907 30685 9919 30719
rect 9861 30679 9919 30685
rect 10042 30676 10048 30728
rect 10100 30716 10106 30728
rect 10336 30716 10364 30824
rect 10410 30744 10416 30796
rect 10468 30784 10474 30796
rect 11333 30787 11391 30793
rect 11333 30784 11345 30787
rect 10468 30756 11345 30784
rect 10468 30744 10474 30756
rect 11333 30753 11345 30756
rect 11379 30753 11391 30787
rect 11333 30747 11391 30753
rect 10100 30688 10456 30716
rect 10100 30676 10106 30688
rect 10428 30660 10456 30688
rect 10410 30608 10416 30660
rect 10468 30608 10474 30660
rect 1578 30580 1584 30592
rect 1539 30552 1584 30580
rect 1578 30540 1584 30552
rect 1636 30540 1642 30592
rect 10042 30580 10048 30592
rect 10003 30552 10048 30580
rect 10042 30540 10048 30552
rect 10100 30540 10106 30592
rect 1104 30490 10856 30512
rect 1104 30438 4213 30490
rect 4265 30438 4277 30490
rect 4329 30438 4341 30490
rect 4393 30438 4405 30490
rect 4457 30438 4469 30490
rect 4521 30438 7477 30490
rect 7529 30438 7541 30490
rect 7593 30438 7605 30490
rect 7657 30438 7669 30490
rect 7721 30438 7733 30490
rect 7785 30438 10856 30490
rect 1104 30416 10856 30438
rect 10134 30308 10140 30320
rect 2746 30280 10140 30308
rect 1397 30243 1455 30249
rect 1397 30209 1409 30243
rect 1443 30240 1455 30243
rect 2746 30240 2774 30280
rect 10134 30268 10140 30280
rect 10192 30268 10198 30320
rect 1443 30212 2774 30240
rect 9861 30243 9919 30249
rect 1443 30209 1455 30212
rect 1397 30203 1455 30209
rect 9861 30209 9873 30243
rect 9907 30240 9919 30243
rect 10594 30240 10600 30252
rect 9907 30212 10600 30240
rect 9907 30209 9919 30212
rect 9861 30203 9919 30209
rect 10594 30200 10600 30212
rect 10652 30200 10658 30252
rect 1578 30036 1584 30048
rect 1539 30008 1584 30036
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 10042 30036 10048 30048
rect 10003 30008 10048 30036
rect 10042 29996 10048 30008
rect 10100 29996 10106 30048
rect 1104 29946 10856 29968
rect 1104 29894 2582 29946
rect 2634 29894 2646 29946
rect 2698 29894 2710 29946
rect 2762 29894 2774 29946
rect 2826 29894 2838 29946
rect 2890 29894 5845 29946
rect 5897 29894 5909 29946
rect 5961 29894 5973 29946
rect 6025 29894 6037 29946
rect 6089 29894 6101 29946
rect 6153 29894 9109 29946
rect 9161 29894 9173 29946
rect 9225 29894 9237 29946
rect 9289 29894 9301 29946
rect 9353 29894 9365 29946
rect 9417 29894 10856 29946
rect 1104 29872 10856 29894
rect 10042 29696 10048 29708
rect 9140 29668 10048 29696
rect 9140 29637 9168 29668
rect 10042 29656 10048 29668
rect 10100 29656 10106 29708
rect 11882 29696 11888 29708
rect 11843 29668 11888 29696
rect 11882 29656 11888 29668
rect 11940 29656 11946 29708
rect 1397 29631 1455 29637
rect 1397 29597 1409 29631
rect 1443 29628 1455 29631
rect 9125 29631 9183 29637
rect 1443 29600 2774 29628
rect 1443 29597 1455 29600
rect 1397 29591 1455 29597
rect 2746 29560 2774 29600
rect 9125 29597 9137 29631
rect 9171 29597 9183 29631
rect 9858 29628 9864 29640
rect 9819 29600 9864 29628
rect 9125 29591 9183 29597
rect 9858 29588 9864 29600
rect 9916 29588 9922 29640
rect 10134 29560 10140 29572
rect 2746 29532 10140 29560
rect 10134 29520 10140 29532
rect 10192 29520 10198 29572
rect 1578 29492 1584 29504
rect 1539 29464 1584 29492
rect 1578 29452 1584 29464
rect 1636 29452 1642 29504
rect 9306 29492 9312 29504
rect 9267 29464 9312 29492
rect 9306 29452 9312 29464
rect 9364 29452 9370 29504
rect 10042 29492 10048 29504
rect 10003 29464 10048 29492
rect 10042 29452 10048 29464
rect 10100 29452 10106 29504
rect 1104 29402 10856 29424
rect 1104 29350 4213 29402
rect 4265 29350 4277 29402
rect 4329 29350 4341 29402
rect 4393 29350 4405 29402
rect 4457 29350 4469 29402
rect 4521 29350 7477 29402
rect 7529 29350 7541 29402
rect 7593 29350 7605 29402
rect 7657 29350 7669 29402
rect 7721 29350 7733 29402
rect 7785 29350 10856 29402
rect 1104 29328 10856 29350
rect 7374 29248 7380 29300
rect 7432 29288 7438 29300
rect 9401 29291 9459 29297
rect 9401 29288 9413 29291
rect 7432 29260 9413 29288
rect 7432 29248 7438 29260
rect 9401 29257 9413 29260
rect 9447 29257 9459 29291
rect 9858 29288 9864 29300
rect 9819 29260 9864 29288
rect 9401 29251 9459 29257
rect 9858 29248 9864 29260
rect 9916 29248 9922 29300
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29152 1455 29155
rect 1946 29152 1952 29164
rect 1443 29124 1952 29152
rect 1443 29121 1455 29124
rect 1397 29115 1455 29121
rect 1946 29112 1952 29124
rect 2004 29112 2010 29164
rect 7282 29112 7288 29164
rect 7340 29152 7346 29164
rect 8665 29155 8723 29161
rect 8665 29152 8677 29155
rect 7340 29124 8677 29152
rect 7340 29112 7346 29124
rect 8665 29121 8677 29124
rect 8711 29121 8723 29155
rect 8665 29115 8723 29121
rect 9769 29155 9827 29161
rect 9769 29121 9781 29155
rect 9815 29121 9827 29155
rect 9769 29115 9827 29121
rect 9217 29087 9275 29093
rect 9217 29084 9229 29087
rect 7300 29056 9229 29084
rect 7300 29028 7328 29056
rect 9217 29053 9229 29056
rect 9263 29084 9275 29087
rect 9784 29084 9812 29115
rect 9263 29056 9812 29084
rect 9263 29053 9275 29056
rect 9217 29047 9275 29053
rect 9858 29044 9864 29096
rect 9916 29084 9922 29096
rect 9953 29087 10011 29093
rect 9953 29084 9965 29087
rect 9916 29056 9965 29084
rect 9916 29044 9922 29056
rect 9953 29053 9965 29056
rect 9999 29084 10011 29087
rect 10410 29084 10416 29096
rect 9999 29056 10416 29084
rect 9999 29053 10011 29056
rect 9953 29047 10011 29053
rect 10410 29044 10416 29056
rect 10468 29044 10474 29096
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 7282 28976 7288 29028
rect 7340 28976 7346 29028
rect 8849 29019 8907 29025
rect 8849 28985 8861 29019
rect 8895 29016 8907 29019
rect 9122 29016 9128 29028
rect 8895 28988 9128 29016
rect 8895 28985 8907 28988
rect 8849 28979 8907 28985
rect 9122 28976 9128 28988
rect 9180 28976 9186 29028
rect 1104 28858 10856 28880
rect 1104 28806 2582 28858
rect 2634 28806 2646 28858
rect 2698 28806 2710 28858
rect 2762 28806 2774 28858
rect 2826 28806 2838 28858
rect 2890 28806 5845 28858
rect 5897 28806 5909 28858
rect 5961 28806 5973 28858
rect 6025 28806 6037 28858
rect 6089 28806 6101 28858
rect 6153 28806 9109 28858
rect 9161 28806 9173 28858
rect 9225 28806 9237 28858
rect 9289 28806 9301 28858
rect 9353 28806 9365 28858
rect 9417 28806 10856 28858
rect 1104 28784 10856 28806
rect 1397 28543 1455 28549
rect 1397 28509 1409 28543
rect 1443 28540 1455 28543
rect 7190 28540 7196 28552
rect 1443 28512 7196 28540
rect 1443 28509 1455 28512
rect 1397 28503 1455 28509
rect 7190 28500 7196 28512
rect 7248 28500 7254 28552
rect 8662 28500 8668 28552
rect 8720 28540 8726 28552
rect 9125 28543 9183 28549
rect 9125 28540 9137 28543
rect 8720 28512 9137 28540
rect 8720 28500 8726 28512
rect 9125 28509 9137 28512
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 9861 28543 9919 28549
rect 9861 28509 9873 28543
rect 9907 28540 9919 28543
rect 10226 28540 10232 28552
rect 9907 28512 10232 28540
rect 9907 28509 9919 28512
rect 9861 28503 9919 28509
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 1578 28404 1584 28416
rect 1539 28376 1584 28404
rect 1578 28364 1584 28376
rect 1636 28364 1642 28416
rect 9306 28404 9312 28416
rect 9267 28376 9312 28404
rect 9306 28364 9312 28376
rect 9364 28364 9370 28416
rect 10045 28407 10103 28413
rect 10045 28373 10057 28407
rect 10091 28404 10103 28407
rect 10134 28404 10140 28416
rect 10091 28376 10140 28404
rect 10091 28373 10103 28376
rect 10045 28367 10103 28373
rect 10134 28364 10140 28376
rect 10192 28364 10198 28416
rect 1104 28314 10856 28336
rect 1104 28262 4213 28314
rect 4265 28262 4277 28314
rect 4329 28262 4341 28314
rect 4393 28262 4405 28314
rect 4457 28262 4469 28314
rect 4521 28262 7477 28314
rect 7529 28262 7541 28314
rect 7593 28262 7605 28314
rect 7657 28262 7669 28314
rect 7721 28262 7733 28314
rect 7785 28262 10856 28314
rect 1104 28240 10856 28262
rect 9769 28203 9827 28209
rect 9769 28169 9781 28203
rect 9815 28200 9827 28203
rect 10226 28200 10232 28212
rect 9815 28172 10232 28200
rect 9815 28169 9827 28172
rect 9769 28163 9827 28169
rect 9876 28073 9904 28172
rect 10226 28160 10232 28172
rect 10284 28160 10290 28212
rect 11238 28160 11244 28212
rect 11296 28200 11302 28212
rect 11882 28200 11888 28212
rect 11296 28172 11888 28200
rect 11296 28160 11302 28172
rect 11882 28160 11888 28172
rect 11940 28160 11946 28212
rect 9861 28067 9919 28073
rect 9861 28033 9873 28067
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 10042 27860 10048 27872
rect 10003 27832 10048 27860
rect 10042 27820 10048 27832
rect 10100 27820 10106 27872
rect 1104 27770 10856 27792
rect 1104 27718 2582 27770
rect 2634 27718 2646 27770
rect 2698 27718 2710 27770
rect 2762 27718 2774 27770
rect 2826 27718 2838 27770
rect 2890 27718 5845 27770
rect 5897 27718 5909 27770
rect 5961 27718 5973 27770
rect 6025 27718 6037 27770
rect 6089 27718 6101 27770
rect 6153 27718 9109 27770
rect 9161 27718 9173 27770
rect 9225 27718 9237 27770
rect 9289 27718 9301 27770
rect 9353 27718 9365 27770
rect 9417 27718 10856 27770
rect 1104 27696 10856 27718
rect 1397 27455 1455 27461
rect 1397 27421 1409 27455
rect 1443 27452 1455 27455
rect 7006 27452 7012 27464
rect 1443 27424 7012 27452
rect 1443 27421 1455 27424
rect 1397 27415 1455 27421
rect 7006 27412 7012 27424
rect 7064 27412 7070 27464
rect 9674 27412 9680 27464
rect 9732 27452 9738 27464
rect 9861 27455 9919 27461
rect 9861 27452 9873 27455
rect 9732 27424 9873 27452
rect 9732 27412 9738 27424
rect 9861 27421 9873 27424
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 10045 27319 10103 27325
rect 10045 27285 10057 27319
rect 10091 27316 10103 27319
rect 10134 27316 10140 27328
rect 10091 27288 10140 27316
rect 10091 27285 10103 27288
rect 10045 27279 10103 27285
rect 10134 27276 10140 27288
rect 10192 27276 10198 27328
rect 1104 27226 10856 27248
rect 1104 27174 4213 27226
rect 4265 27174 4277 27226
rect 4329 27174 4341 27226
rect 4393 27174 4405 27226
rect 4457 27174 4469 27226
rect 4521 27174 7477 27226
rect 7529 27174 7541 27226
rect 7593 27174 7605 27226
rect 7657 27174 7669 27226
rect 7721 27174 7733 27226
rect 7785 27174 10856 27226
rect 1104 27152 10856 27174
rect 8110 27044 8116 27056
rect 2746 27016 8116 27044
rect 1397 26979 1455 26985
rect 1397 26945 1409 26979
rect 1443 26976 1455 26979
rect 2746 26976 2774 27016
rect 8110 27004 8116 27016
rect 8168 27004 8174 27056
rect 8846 27004 8852 27056
rect 8904 27044 8910 27056
rect 8904 27016 9076 27044
rect 8904 27004 8910 27016
rect 1443 26948 2774 26976
rect 1443 26945 1455 26948
rect 1397 26939 1455 26945
rect 7190 26936 7196 26988
rect 7248 26976 7254 26988
rect 7926 26976 7932 26988
rect 7248 26948 7932 26976
rect 7248 26936 7254 26948
rect 7926 26936 7932 26948
rect 7984 26936 7990 26988
rect 8662 26936 8668 26988
rect 8720 26976 8726 26988
rect 8938 26976 8944 26988
rect 8720 26948 8944 26976
rect 8720 26936 8726 26948
rect 8938 26936 8944 26948
rect 8996 26936 9002 26988
rect 9048 26784 9076 27016
rect 9766 26936 9772 26988
rect 9824 26976 9830 26988
rect 9861 26979 9919 26985
rect 9861 26976 9873 26979
rect 9824 26948 9873 26976
rect 9824 26936 9830 26948
rect 9861 26945 9873 26948
rect 9907 26945 9919 26979
rect 9861 26939 9919 26945
rect 1578 26772 1584 26784
rect 1539 26744 1584 26772
rect 1578 26732 1584 26744
rect 1636 26732 1642 26784
rect 9030 26732 9036 26784
rect 9088 26732 9094 26784
rect 10042 26772 10048 26784
rect 10003 26744 10048 26772
rect 10042 26732 10048 26744
rect 10100 26732 10106 26784
rect 1104 26682 10856 26704
rect 1104 26630 2582 26682
rect 2634 26630 2646 26682
rect 2698 26630 2710 26682
rect 2762 26630 2774 26682
rect 2826 26630 2838 26682
rect 2890 26630 5845 26682
rect 5897 26630 5909 26682
rect 5961 26630 5973 26682
rect 6025 26630 6037 26682
rect 6089 26630 6101 26682
rect 6153 26630 9109 26682
rect 9161 26630 9173 26682
rect 9225 26630 9237 26682
rect 9289 26630 9301 26682
rect 9353 26630 9365 26682
rect 9417 26630 10856 26682
rect 1104 26608 10856 26630
rect 8938 26528 8944 26580
rect 8996 26568 9002 26580
rect 9490 26568 9496 26580
rect 8996 26540 9496 26568
rect 8996 26528 9002 26540
rect 9490 26528 9496 26540
rect 9548 26528 9554 26580
rect 7926 26460 7932 26512
rect 7984 26500 7990 26512
rect 8110 26500 8116 26512
rect 7984 26472 8116 26500
rect 7984 26460 7990 26472
rect 8110 26460 8116 26472
rect 8168 26460 8174 26512
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26364 1455 26367
rect 3602 26364 3608 26376
rect 1443 26336 3608 26364
rect 1443 26333 1455 26336
rect 1397 26327 1455 26333
rect 3602 26324 3608 26336
rect 3660 26324 3666 26376
rect 9861 26367 9919 26373
rect 9861 26333 9873 26367
rect 9907 26364 9919 26367
rect 9950 26364 9956 26376
rect 9907 26336 9956 26364
rect 9907 26333 9919 26336
rect 9861 26327 9919 26333
rect 9950 26324 9956 26336
rect 10008 26324 10014 26376
rect 10594 26324 10600 26376
rect 10652 26364 10658 26376
rect 10965 26367 11023 26373
rect 10965 26364 10977 26367
rect 10652 26336 10977 26364
rect 10652 26324 10658 26336
rect 10965 26333 10977 26336
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 1578 26228 1584 26240
rect 1539 26200 1584 26228
rect 1578 26188 1584 26200
rect 1636 26188 1642 26240
rect 10045 26231 10103 26237
rect 10045 26197 10057 26231
rect 10091 26228 10103 26231
rect 10965 26231 11023 26237
rect 10965 26228 10977 26231
rect 10091 26200 10977 26228
rect 10091 26197 10103 26200
rect 10045 26191 10103 26197
rect 10965 26197 10977 26200
rect 11011 26197 11023 26231
rect 10965 26191 11023 26197
rect 1104 26138 10856 26160
rect 1104 26086 4213 26138
rect 4265 26086 4277 26138
rect 4329 26086 4341 26138
rect 4393 26086 4405 26138
rect 4457 26086 4469 26138
rect 4521 26086 7477 26138
rect 7529 26086 7541 26138
rect 7593 26086 7605 26138
rect 7657 26086 7669 26138
rect 7721 26086 7733 26138
rect 7785 26086 10856 26138
rect 1104 26064 10856 26086
rect 6730 25984 6736 26036
rect 6788 26024 6794 26036
rect 10045 26027 10103 26033
rect 10045 26024 10057 26027
rect 6788 25996 10057 26024
rect 6788 25984 6794 25996
rect 10045 25993 10057 25996
rect 10091 25993 10103 26027
rect 10045 25987 10103 25993
rect 11606 25956 11612 25968
rect 2746 25928 11612 25956
rect 1397 25891 1455 25897
rect 1397 25857 1409 25891
rect 1443 25888 1455 25891
rect 2746 25888 2774 25928
rect 11606 25916 11612 25928
rect 11664 25916 11670 25968
rect 1443 25860 2774 25888
rect 1443 25857 1455 25860
rect 1397 25851 1455 25857
rect 8478 25848 8484 25900
rect 8536 25888 8542 25900
rect 9125 25891 9183 25897
rect 9125 25888 9137 25891
rect 8536 25860 9137 25888
rect 8536 25848 8542 25860
rect 9125 25857 9137 25860
rect 9171 25857 9183 25891
rect 9858 25888 9864 25900
rect 9819 25860 9864 25888
rect 9125 25851 9183 25857
rect 9858 25848 9864 25860
rect 9916 25848 9922 25900
rect 1578 25684 1584 25696
rect 1539 25656 1584 25684
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 9309 25687 9367 25693
rect 9309 25653 9321 25687
rect 9355 25684 9367 25687
rect 9490 25684 9496 25696
rect 9355 25656 9496 25684
rect 9355 25653 9367 25656
rect 9309 25647 9367 25653
rect 9490 25644 9496 25656
rect 9548 25644 9554 25696
rect 1104 25594 10856 25616
rect 1104 25542 2582 25594
rect 2634 25542 2646 25594
rect 2698 25542 2710 25594
rect 2762 25542 2774 25594
rect 2826 25542 2838 25594
rect 2890 25542 5845 25594
rect 5897 25542 5909 25594
rect 5961 25542 5973 25594
rect 6025 25542 6037 25594
rect 6089 25542 6101 25594
rect 6153 25542 9109 25594
rect 9161 25542 9173 25594
rect 9225 25542 9237 25594
rect 9289 25542 9301 25594
rect 9353 25542 9365 25594
rect 9417 25542 10856 25594
rect 1104 25520 10856 25542
rect 10410 25372 10416 25424
rect 10468 25412 10474 25424
rect 10962 25412 10968 25424
rect 10468 25384 10968 25412
rect 10468 25372 10474 25384
rect 10962 25372 10968 25384
rect 11020 25372 11026 25424
rect 9950 25344 9956 25356
rect 9911 25316 9956 25344
rect 9950 25304 9956 25316
rect 10008 25304 10014 25356
rect 10962 25276 10968 25288
rect 10923 25248 10968 25276
rect 10962 25236 10968 25248
rect 11020 25236 11026 25288
rect 1026 25168 1032 25220
rect 1084 25208 1090 25220
rect 9861 25211 9919 25217
rect 9861 25208 9873 25211
rect 1084 25180 9873 25208
rect 1084 25168 1090 25180
rect 9861 25177 9873 25180
rect 9907 25177 9919 25211
rect 9861 25171 9919 25177
rect 8478 25100 8484 25152
rect 8536 25140 8542 25152
rect 9401 25143 9459 25149
rect 9401 25140 9413 25143
rect 8536 25112 9413 25140
rect 8536 25100 8542 25112
rect 9401 25109 9413 25112
rect 9447 25109 9459 25143
rect 9766 25140 9772 25152
rect 9727 25112 9772 25140
rect 9401 25103 9459 25109
rect 9766 25100 9772 25112
rect 9824 25100 9830 25152
rect 1104 25050 10856 25072
rect 1104 24998 4213 25050
rect 4265 24998 4277 25050
rect 4329 24998 4341 25050
rect 4393 24998 4405 25050
rect 4457 24998 4469 25050
rect 4521 24998 7477 25050
rect 7529 24998 7541 25050
rect 7593 24998 7605 25050
rect 7657 24998 7669 25050
rect 7721 24998 7733 25050
rect 7785 24998 10856 25050
rect 1104 24976 10856 24998
rect 1397 24803 1455 24809
rect 1397 24769 1409 24803
rect 1443 24800 1455 24803
rect 7098 24800 7104 24812
rect 1443 24772 7104 24800
rect 1443 24769 1455 24772
rect 1397 24763 1455 24769
rect 7098 24760 7104 24772
rect 7156 24760 7162 24812
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24800 9183 24803
rect 9490 24800 9496 24812
rect 9171 24772 9496 24800
rect 9171 24769 9183 24772
rect 9125 24763 9183 24769
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 9950 24800 9956 24812
rect 9911 24772 9956 24800
rect 9950 24760 9956 24772
rect 10008 24760 10014 24812
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24800 10195 24803
rect 10318 24800 10324 24812
rect 10183 24772 10324 24800
rect 10183 24769 10195 24772
rect 10137 24763 10195 24769
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 1578 24664 1584 24676
rect 1539 24636 1584 24664
rect 1578 24624 1584 24636
rect 1636 24624 1642 24676
rect 9309 24667 9367 24673
rect 9309 24633 9321 24667
rect 9355 24664 9367 24667
rect 11790 24664 11796 24676
rect 9355 24636 11796 24664
rect 9355 24633 9367 24636
rect 9309 24627 9367 24633
rect 11790 24624 11796 24636
rect 11848 24624 11854 24676
rect 1104 24506 10856 24528
rect 1104 24454 2582 24506
rect 2634 24454 2646 24506
rect 2698 24454 2710 24506
rect 2762 24454 2774 24506
rect 2826 24454 2838 24506
rect 2890 24454 5845 24506
rect 5897 24454 5909 24506
rect 5961 24454 5973 24506
rect 6025 24454 6037 24506
rect 6089 24454 6101 24506
rect 6153 24454 9109 24506
rect 9161 24454 9173 24506
rect 9225 24454 9237 24506
rect 9289 24454 9301 24506
rect 9353 24454 9365 24506
rect 9417 24454 10856 24506
rect 1104 24432 10856 24454
rect 4062 24352 4068 24404
rect 4120 24392 4126 24404
rect 9309 24395 9367 24401
rect 9309 24392 9321 24395
rect 4120 24364 9321 24392
rect 4120 24352 4126 24364
rect 9309 24361 9321 24364
rect 9355 24361 9367 24395
rect 9309 24355 9367 24361
rect 10137 24327 10195 24333
rect 10137 24293 10149 24327
rect 10183 24324 10195 24327
rect 10502 24324 10508 24336
rect 10183 24296 10508 24324
rect 10183 24293 10195 24296
rect 10137 24287 10195 24293
rect 10502 24284 10508 24296
rect 10560 24284 10566 24336
rect 1397 24191 1455 24197
rect 1397 24157 1409 24191
rect 1443 24188 1455 24191
rect 4798 24188 4804 24200
rect 1443 24160 4804 24188
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 9122 24188 9128 24200
rect 9083 24160 9128 24188
rect 9122 24148 9128 24160
rect 9180 24148 9186 24200
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10042 24188 10048 24200
rect 9999 24160 10048 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 10042 24148 10048 24160
rect 10100 24148 10106 24200
rect 11241 24191 11299 24197
rect 11241 24157 11253 24191
rect 11287 24188 11299 24191
rect 11790 24188 11796 24200
rect 11287 24160 11796 24188
rect 11287 24157 11299 24160
rect 11241 24151 11299 24157
rect 11790 24148 11796 24160
rect 11848 24148 11854 24200
rect 9490 24080 9496 24132
rect 9548 24120 9554 24132
rect 11698 24120 11704 24132
rect 9548 24092 11704 24120
rect 9548 24080 9554 24092
rect 11698 24080 11704 24092
rect 11756 24080 11762 24132
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 1104 23962 10856 23984
rect 1104 23910 4213 23962
rect 4265 23910 4277 23962
rect 4329 23910 4341 23962
rect 4393 23910 4405 23962
rect 4457 23910 4469 23962
rect 4521 23910 7477 23962
rect 7529 23910 7541 23962
rect 7593 23910 7605 23962
rect 7657 23910 7669 23962
rect 7721 23910 7733 23962
rect 7785 23910 10856 23962
rect 1104 23888 10856 23910
rect 8754 23808 8760 23860
rect 8812 23848 8818 23860
rect 8849 23851 8907 23857
rect 8849 23848 8861 23851
rect 8812 23820 8861 23848
rect 8812 23808 8818 23820
rect 8849 23817 8861 23820
rect 8895 23817 8907 23851
rect 8849 23811 8907 23817
rect 9309 23851 9367 23857
rect 9309 23817 9321 23851
rect 9355 23848 9367 23851
rect 9861 23851 9919 23857
rect 9861 23848 9873 23851
rect 9355 23820 9873 23848
rect 9355 23817 9367 23820
rect 9309 23811 9367 23817
rect 9861 23817 9873 23820
rect 9907 23848 9919 23851
rect 11514 23848 11520 23860
rect 9907 23820 11520 23848
rect 9907 23817 9919 23820
rect 9861 23811 9919 23817
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23712 1455 23715
rect 3418 23712 3424 23724
rect 1443 23684 3424 23712
rect 1443 23681 1455 23684
rect 1397 23675 1455 23681
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 8754 23712 8760 23724
rect 8715 23684 8760 23712
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 9674 23672 9680 23724
rect 9732 23712 9738 23724
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 9732 23684 9781 23712
rect 9732 23672 9738 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 10045 23647 10103 23653
rect 10045 23613 10057 23647
rect 10091 23644 10103 23647
rect 10134 23644 10140 23656
rect 10091 23616 10140 23644
rect 10091 23613 10103 23616
rect 10045 23607 10103 23613
rect 10134 23604 10140 23616
rect 10192 23604 10198 23656
rect 6730 23536 6736 23588
rect 6788 23576 6794 23588
rect 9401 23579 9459 23585
rect 9401 23576 9413 23579
rect 6788 23548 9413 23576
rect 6788 23536 6794 23548
rect 9401 23545 9413 23548
rect 9447 23545 9459 23579
rect 9401 23539 9459 23545
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 1104 23418 10856 23440
rect 1104 23366 2582 23418
rect 2634 23366 2646 23418
rect 2698 23366 2710 23418
rect 2762 23366 2774 23418
rect 2826 23366 2838 23418
rect 2890 23366 5845 23418
rect 5897 23366 5909 23418
rect 5961 23366 5973 23418
rect 6025 23366 6037 23418
rect 6089 23366 6101 23418
rect 6153 23366 9109 23418
rect 9161 23366 9173 23418
rect 9225 23366 9237 23418
rect 9289 23366 9301 23418
rect 9353 23366 9365 23418
rect 9417 23366 10856 23418
rect 1104 23344 10856 23366
rect 5442 23128 5448 23180
rect 5500 23168 5506 23180
rect 9861 23171 9919 23177
rect 9861 23168 9873 23171
rect 5500 23140 9873 23168
rect 5500 23128 5506 23140
rect 9861 23137 9873 23140
rect 9907 23137 9919 23171
rect 9861 23131 9919 23137
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23168 10103 23171
rect 10134 23168 10140 23180
rect 10091 23140 10140 23168
rect 10091 23137 10103 23140
rect 10045 23131 10103 23137
rect 10134 23128 10140 23140
rect 10192 23128 10198 23180
rect 1397 23103 1455 23109
rect 1397 23069 1409 23103
rect 1443 23100 1455 23103
rect 9030 23100 9036 23112
rect 1443 23072 9036 23100
rect 1443 23069 1455 23072
rect 1397 23063 1455 23069
rect 9030 23060 9036 23072
rect 9088 23060 9094 23112
rect 9769 23035 9827 23041
rect 9769 23001 9781 23035
rect 9815 23032 9827 23035
rect 10134 23032 10140 23044
rect 9815 23004 10140 23032
rect 9815 23001 9827 23004
rect 9769 22995 9827 23001
rect 10134 22992 10140 23004
rect 10192 22992 10198 23044
rect 1578 22964 1584 22976
rect 1539 22936 1584 22964
rect 1578 22924 1584 22936
rect 1636 22924 1642 22976
rect 5626 22924 5632 22976
rect 5684 22964 5690 22976
rect 9401 22967 9459 22973
rect 9401 22964 9413 22967
rect 5684 22936 9413 22964
rect 5684 22924 5690 22936
rect 9401 22933 9413 22936
rect 9447 22933 9459 22967
rect 9401 22927 9459 22933
rect 1104 22874 10856 22896
rect 1104 22822 4213 22874
rect 4265 22822 4277 22874
rect 4329 22822 4341 22874
rect 4393 22822 4405 22874
rect 4457 22822 4469 22874
rect 4521 22822 7477 22874
rect 7529 22822 7541 22874
rect 7593 22822 7605 22874
rect 7657 22822 7669 22874
rect 7721 22822 7733 22874
rect 7785 22822 10856 22874
rect 1104 22800 10856 22822
rect 3786 22720 3792 22772
rect 3844 22760 3850 22772
rect 8665 22763 8723 22769
rect 8665 22760 8677 22763
rect 3844 22732 8677 22760
rect 3844 22720 3850 22732
rect 8665 22729 8677 22732
rect 8711 22729 8723 22763
rect 8665 22723 8723 22729
rect 11146 22720 11152 22772
rect 11204 22760 11210 22772
rect 11885 22763 11943 22769
rect 11885 22760 11897 22763
rect 11204 22732 11897 22760
rect 11204 22720 11210 22732
rect 11885 22729 11897 22732
rect 11931 22729 11943 22763
rect 11885 22723 11943 22729
rect 6546 22652 6552 22704
rect 6604 22692 6610 22704
rect 9861 22695 9919 22701
rect 9861 22692 9873 22695
rect 6604 22664 9873 22692
rect 6604 22652 6610 22664
rect 9861 22661 9873 22664
rect 9907 22661 9919 22695
rect 9861 22655 9919 22661
rect 10318 22652 10324 22704
rect 10376 22692 10382 22704
rect 11425 22695 11483 22701
rect 11425 22692 11437 22695
rect 10376 22664 11437 22692
rect 10376 22652 10382 22664
rect 11425 22661 11437 22664
rect 11471 22661 11483 22695
rect 11425 22655 11483 22661
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22624 1455 22627
rect 4890 22624 4896 22636
rect 1443 22596 4896 22624
rect 1443 22593 1455 22596
rect 1397 22587 1455 22593
rect 4890 22584 4896 22596
rect 4948 22584 4954 22636
rect 7098 22584 7104 22636
rect 7156 22624 7162 22636
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 7156 22596 8585 22624
rect 7156 22584 7162 22596
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 9766 22624 9772 22636
rect 9727 22596 9772 22624
rect 8573 22587 8631 22593
rect 9766 22584 9772 22596
rect 9824 22584 9830 22636
rect 11149 22627 11207 22633
rect 11149 22593 11161 22627
rect 11195 22593 11207 22627
rect 11149 22587 11207 22593
rect 8754 22516 8760 22568
rect 8812 22556 8818 22568
rect 8849 22559 8907 22565
rect 8849 22556 8861 22559
rect 8812 22528 8861 22556
rect 8812 22516 8818 22528
rect 8849 22525 8861 22528
rect 8895 22556 8907 22559
rect 10045 22559 10103 22565
rect 10045 22556 10057 22559
rect 8895 22528 10057 22556
rect 8895 22525 8907 22528
rect 8849 22519 8907 22525
rect 10045 22525 10057 22528
rect 10091 22556 10103 22559
rect 10226 22556 10232 22568
rect 10091 22528 10232 22556
rect 10091 22525 10103 22528
rect 10045 22519 10103 22525
rect 10226 22516 10232 22528
rect 10284 22516 10290 22568
rect 6178 22448 6184 22500
rect 6236 22488 6242 22500
rect 9401 22491 9459 22497
rect 9401 22488 9413 22491
rect 6236 22460 9413 22488
rect 6236 22448 6242 22460
rect 9401 22457 9413 22460
rect 9447 22457 9459 22491
rect 9401 22451 9459 22457
rect 10778 22448 10784 22500
rect 10836 22488 10842 22500
rect 10836 22460 11100 22488
rect 10836 22448 10842 22460
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 7834 22380 7840 22432
rect 7892 22420 7898 22432
rect 8205 22423 8263 22429
rect 8205 22420 8217 22423
rect 7892 22392 8217 22420
rect 7892 22380 7898 22392
rect 8205 22389 8217 22392
rect 8251 22389 8263 22423
rect 8205 22383 8263 22389
rect 1104 22330 10856 22352
rect 1104 22278 2582 22330
rect 2634 22278 2646 22330
rect 2698 22278 2710 22330
rect 2762 22278 2774 22330
rect 2826 22278 2838 22330
rect 2890 22278 5845 22330
rect 5897 22278 5909 22330
rect 5961 22278 5973 22330
rect 6025 22278 6037 22330
rect 6089 22278 6101 22330
rect 6153 22278 9109 22330
rect 9161 22278 9173 22330
rect 9225 22278 9237 22330
rect 9289 22278 9301 22330
rect 9353 22278 9365 22330
rect 9417 22278 10856 22330
rect 11072 22296 11100 22460
rect 11164 22420 11192 22587
rect 11238 22420 11244 22432
rect 11164 22392 11244 22420
rect 11238 22380 11244 22392
rect 11296 22380 11302 22432
rect 1104 22256 10856 22278
rect 11054 22244 11060 22296
rect 11112 22244 11118 22296
rect 11330 22244 11336 22296
rect 11388 22244 11394 22296
rect 11609 22287 11667 22293
rect 11609 22253 11621 22287
rect 11655 22284 11667 22287
rect 11698 22284 11704 22296
rect 11655 22256 11704 22284
rect 11655 22253 11667 22256
rect 11609 22247 11667 22253
rect 11698 22244 11704 22256
rect 11756 22244 11762 22296
rect 11348 22216 11376 22244
rect 11348 22188 11652 22216
rect 10962 22108 10968 22160
rect 11020 22148 11026 22160
rect 11624 22157 11652 22188
rect 11333 22151 11391 22157
rect 11333 22148 11345 22151
rect 11020 22120 11345 22148
rect 11020 22108 11026 22120
rect 11333 22117 11345 22120
rect 11379 22117 11391 22151
rect 11333 22111 11391 22117
rect 11609 22151 11667 22157
rect 11609 22117 11621 22151
rect 11655 22117 11667 22151
rect 11609 22111 11667 22117
rect 8294 22040 8300 22092
rect 8352 22080 8358 22092
rect 8389 22083 8447 22089
rect 8389 22080 8401 22083
rect 8352 22052 8401 22080
rect 8352 22040 8358 22052
rect 8389 22049 8401 22052
rect 8435 22049 8447 22083
rect 8389 22043 8447 22049
rect 9585 22083 9643 22089
rect 9585 22049 9597 22083
rect 9631 22080 9643 22083
rect 10318 22080 10324 22092
rect 9631 22052 10324 22080
rect 9631 22049 9643 22052
rect 9585 22043 9643 22049
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 11514 22040 11520 22092
rect 11572 22080 11578 22092
rect 11572 22052 11617 22080
rect 11572 22040 11578 22052
rect 9306 22012 9312 22024
rect 9267 21984 9312 22012
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 10410 21972 10416 22024
rect 10468 22012 10474 22024
rect 10965 22015 11023 22021
rect 10965 22012 10977 22015
rect 10468 21984 10977 22012
rect 10468 21972 10474 21984
rect 10965 21981 10977 21984
rect 11011 21981 11023 22015
rect 10965 21975 11023 21981
rect 8110 21904 8116 21956
rect 8168 21944 8174 21956
rect 8205 21947 8263 21953
rect 8205 21944 8217 21947
rect 8168 21916 8217 21944
rect 8168 21904 8174 21916
rect 8205 21913 8217 21916
rect 8251 21913 8263 21947
rect 8205 21907 8263 21913
rect 11149 21947 11207 21953
rect 11149 21913 11161 21947
rect 11195 21944 11207 21947
rect 11238 21944 11244 21956
rect 11195 21916 11244 21944
rect 11195 21913 11207 21916
rect 11149 21907 11207 21913
rect 11238 21904 11244 21916
rect 11296 21904 11302 21956
rect 11333 21947 11391 21953
rect 11333 21913 11345 21947
rect 11379 21913 11391 21947
rect 11333 21907 11391 21913
rect 11425 21947 11483 21953
rect 11425 21913 11437 21947
rect 11471 21913 11483 21947
rect 11425 21907 11483 21913
rect 5258 21836 5264 21888
rect 5316 21876 5322 21888
rect 9766 21876 9772 21888
rect 5316 21848 9772 21876
rect 5316 21836 5322 21848
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 11348 21817 11376 21907
rect 11440 21817 11468 21907
rect 11790 21904 11796 21956
rect 11848 21944 11854 21956
rect 11885 21947 11943 21953
rect 11885 21944 11897 21947
rect 11848 21916 11897 21944
rect 11848 21904 11854 21916
rect 11885 21913 11897 21916
rect 11931 21913 11943 21947
rect 11885 21907 11943 21913
rect 11517 21879 11575 21885
rect 11517 21845 11529 21879
rect 11563 21876 11575 21879
rect 11606 21876 11612 21888
rect 11563 21848 11612 21876
rect 11563 21845 11575 21848
rect 11517 21839 11575 21845
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 11333 21811 11391 21817
rect 1104 21786 10856 21808
rect 1104 21734 4213 21786
rect 4265 21734 4277 21786
rect 4329 21734 4341 21786
rect 4393 21734 4405 21786
rect 4457 21734 4469 21786
rect 4521 21734 7477 21786
rect 7529 21734 7541 21786
rect 7593 21734 7605 21786
rect 7657 21734 7669 21786
rect 7721 21734 7733 21786
rect 7785 21734 10856 21786
rect 11333 21777 11345 21811
rect 11379 21777 11391 21811
rect 11333 21771 11391 21777
rect 11425 21811 11483 21817
rect 11425 21777 11437 21811
rect 11471 21777 11483 21811
rect 11425 21771 11483 21777
rect 1104 21712 10856 21734
rect 11054 21700 11060 21752
rect 11112 21740 11118 21752
rect 11517 21743 11575 21749
rect 11517 21740 11529 21743
rect 11112 21712 11529 21740
rect 11112 21700 11118 21712
rect 11517 21709 11529 21712
rect 11563 21709 11575 21743
rect 11517 21703 11575 21709
rect 11609 21743 11667 21749
rect 11609 21709 11621 21743
rect 11655 21740 11667 21743
rect 11698 21740 11704 21752
rect 11655 21712 11704 21740
rect 11655 21709 11667 21712
rect 11609 21703 11667 21709
rect 11698 21700 11704 21712
rect 11756 21700 11762 21752
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 8573 21675 8631 21681
rect 8573 21672 8585 21675
rect 3568 21644 8585 21672
rect 3568 21632 3574 21644
rect 8573 21641 8585 21644
rect 8619 21641 8631 21675
rect 8573 21635 8631 21641
rect 8481 21607 8539 21613
rect 8481 21573 8493 21607
rect 8527 21604 8539 21607
rect 10226 21604 10232 21616
rect 8527 21576 10232 21604
rect 8527 21573 8539 21576
rect 8481 21567 8539 21573
rect 10226 21564 10232 21576
rect 10284 21564 10290 21616
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21536 1455 21539
rect 7374 21536 7380 21548
rect 1443 21508 7380 21536
rect 1443 21505 1455 21508
rect 1397 21499 1455 21505
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 10778 21536 10784 21548
rect 9631 21508 10784 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 10778 21496 10784 21508
rect 10836 21496 10842 21548
rect 8754 21468 8760 21480
rect 8715 21440 8760 21468
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 9309 21471 9367 21477
rect 9309 21437 9321 21471
rect 9355 21468 9367 21471
rect 9490 21468 9496 21480
rect 9355 21440 9496 21468
rect 9355 21437 9367 21440
rect 9309 21431 9367 21437
rect 9490 21428 9496 21440
rect 9548 21428 9554 21480
rect 1578 21400 1584 21412
rect 1539 21372 1584 21400
rect 1578 21360 1584 21372
rect 1636 21360 1642 21412
rect 8772 21400 8800 21428
rect 9950 21400 9956 21412
rect 8772 21372 9956 21400
rect 9950 21360 9956 21372
rect 10008 21360 10014 21412
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 1762 21332 1768 21344
rect 1452 21304 1768 21332
rect 1452 21292 1458 21304
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 8113 21335 8171 21341
rect 8113 21332 8125 21335
rect 6972 21304 8125 21332
rect 6972 21292 6978 21304
rect 8113 21301 8125 21304
rect 8159 21301 8171 21335
rect 8113 21295 8171 21301
rect 8754 21292 8760 21344
rect 8812 21332 8818 21344
rect 9582 21332 9588 21344
rect 8812 21304 9588 21332
rect 8812 21292 8818 21304
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 1104 21242 10856 21264
rect 1104 21190 2582 21242
rect 2634 21190 2646 21242
rect 2698 21190 2710 21242
rect 2762 21190 2774 21242
rect 2826 21190 2838 21242
rect 2890 21190 5845 21242
rect 5897 21190 5909 21242
rect 5961 21190 5973 21242
rect 6025 21190 6037 21242
rect 6089 21190 6101 21242
rect 6153 21190 9109 21242
rect 9161 21190 9173 21242
rect 9225 21190 9237 21242
rect 9289 21190 9301 21242
rect 9353 21190 9365 21242
rect 9417 21190 10856 21242
rect 1104 21168 10856 21190
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20992 9643 20995
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 9631 20964 11161 20992
rect 9631 20961 9643 20964
rect 9585 20955 9643 20961
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 1397 20927 1455 20933
rect 1397 20893 1409 20927
rect 1443 20924 1455 20927
rect 8478 20924 8484 20936
rect 1443 20896 8484 20924
rect 1443 20893 1455 20896
rect 1397 20887 1455 20893
rect 8478 20884 8484 20896
rect 8536 20884 8542 20936
rect 9306 20924 9312 20936
rect 9267 20896 9312 20924
rect 9306 20884 9312 20896
rect 9364 20884 9370 20936
rect 11146 20856 11152 20868
rect 11107 20828 11152 20856
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 1578 20788 1584 20800
rect 1539 20760 1584 20788
rect 1578 20748 1584 20760
rect 1636 20748 1642 20800
rect 1104 20698 10856 20720
rect 1104 20646 4213 20698
rect 4265 20646 4277 20698
rect 4329 20646 4341 20698
rect 4393 20646 4405 20698
rect 4457 20646 4469 20698
rect 4521 20646 7477 20698
rect 7529 20646 7541 20698
rect 7593 20646 7605 20698
rect 7657 20646 7669 20698
rect 7721 20646 7733 20698
rect 7785 20646 10856 20698
rect 1104 20624 10856 20646
rect 8018 20544 8024 20596
rect 8076 20584 8082 20596
rect 8113 20587 8171 20593
rect 8113 20584 8125 20587
rect 8076 20556 8125 20584
rect 8076 20544 8082 20556
rect 8113 20553 8125 20556
rect 8159 20553 8171 20587
rect 8113 20547 8171 20553
rect 8757 20587 8815 20593
rect 8757 20553 8769 20587
rect 8803 20584 8815 20587
rect 10594 20584 10600 20596
rect 8803 20556 10600 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 10594 20544 10600 20556
rect 10652 20544 10658 20596
rect 8662 20476 8668 20528
rect 8720 20516 8726 20528
rect 9217 20519 9275 20525
rect 9217 20516 9229 20519
rect 8720 20488 9229 20516
rect 8720 20476 8726 20488
rect 9217 20485 9229 20488
rect 9263 20516 9275 20519
rect 9582 20516 9588 20528
rect 9263 20488 9588 20516
rect 9263 20485 9275 20488
rect 9217 20479 9275 20485
rect 9582 20476 9588 20488
rect 9640 20516 9646 20528
rect 10229 20519 10287 20525
rect 10229 20516 10241 20519
rect 9640 20488 10241 20516
rect 9640 20476 9646 20488
rect 10229 20485 10241 20488
rect 10275 20485 10287 20519
rect 10229 20479 10287 20485
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20448 1455 20451
rect 6730 20448 6736 20460
rect 1443 20420 6736 20448
rect 1443 20417 1455 20420
rect 1397 20411 1455 20417
rect 6730 20408 6736 20420
rect 6788 20408 6794 20460
rect 8110 20408 8116 20460
rect 8168 20448 8174 20460
rect 8297 20451 8355 20457
rect 8297 20448 8309 20451
rect 8168 20420 8309 20448
rect 8168 20408 8174 20420
rect 8297 20417 8309 20420
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20448 8999 20451
rect 9490 20448 9496 20460
rect 8987 20420 9496 20448
rect 8987 20417 8999 20420
rect 8941 20411 8999 20417
rect 9490 20408 9496 20420
rect 9548 20408 9554 20460
rect 8294 20272 8300 20324
rect 8352 20312 8358 20324
rect 8938 20312 8944 20324
rect 8352 20284 8944 20312
rect 8352 20272 8358 20284
rect 8938 20272 8944 20284
rect 8996 20272 9002 20324
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1104 20154 10856 20176
rect 1104 20102 2582 20154
rect 2634 20102 2646 20154
rect 2698 20102 2710 20154
rect 2762 20102 2774 20154
rect 2826 20102 2838 20154
rect 2890 20102 5845 20154
rect 5897 20102 5909 20154
rect 5961 20102 5973 20154
rect 6025 20102 6037 20154
rect 6089 20102 6101 20154
rect 6153 20102 9109 20154
rect 9161 20102 9173 20154
rect 9225 20102 9237 20154
rect 9289 20102 9301 20154
rect 9353 20102 9365 20154
rect 9417 20102 10856 20154
rect 1104 20080 10856 20102
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 8205 20043 8263 20049
rect 8205 20040 8217 20043
rect 7984 20012 8217 20040
rect 7984 20000 7990 20012
rect 8205 20009 8217 20012
rect 8251 20009 8263 20043
rect 8205 20003 8263 20009
rect 8754 19932 8760 19984
rect 8812 19972 8818 19984
rect 9306 19972 9312 19984
rect 8812 19944 9312 19972
rect 8812 19932 8818 19944
rect 9306 19932 9312 19944
rect 9364 19932 9370 19984
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 9640 19876 9873 19904
rect 9640 19864 9646 19876
rect 9861 19873 9873 19876
rect 9907 19873 9919 19907
rect 9861 19867 9919 19873
rect 9950 19864 9956 19916
rect 10008 19904 10014 19916
rect 10318 19904 10324 19916
rect 10008 19876 10324 19904
rect 10008 19864 10014 19876
rect 10318 19864 10324 19876
rect 10376 19864 10382 19916
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19836 1455 19839
rect 7834 19836 7840 19848
rect 1443 19808 7840 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 8168 19808 8401 19836
rect 8168 19796 8174 19808
rect 8389 19805 8401 19808
rect 8435 19805 8447 19839
rect 8389 19799 8447 19805
rect 1578 19700 1584 19712
rect 1539 19672 1584 19700
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 9401 19703 9459 19709
rect 9401 19700 9413 19703
rect 7064 19672 9413 19700
rect 7064 19660 7070 19672
rect 9401 19669 9413 19672
rect 9447 19669 9459 19703
rect 9401 19663 9459 19669
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 10042 19700 10048 19712
rect 9815 19672 10048 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 1104 19610 10856 19632
rect 1104 19558 4213 19610
rect 4265 19558 4277 19610
rect 4329 19558 4341 19610
rect 4393 19558 4405 19610
rect 4457 19558 4469 19610
rect 4521 19558 7477 19610
rect 7529 19558 7541 19610
rect 7593 19558 7605 19610
rect 7657 19558 7669 19610
rect 7721 19558 7733 19610
rect 7785 19558 10856 19610
rect 1104 19536 10856 19558
rect 8113 19499 8171 19505
rect 8113 19465 8125 19499
rect 8159 19496 8171 19499
rect 8294 19496 8300 19508
rect 8159 19468 8300 19496
rect 8159 19465 8171 19468
rect 8113 19459 8171 19465
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 8757 19499 8815 19505
rect 8757 19465 8769 19499
rect 8803 19465 8815 19499
rect 8757 19459 8815 19465
rect 9125 19499 9183 19505
rect 9125 19465 9137 19499
rect 9171 19496 9183 19499
rect 9171 19468 9812 19496
rect 9171 19465 9183 19468
rect 9125 19459 9183 19465
rect 7926 19388 7932 19440
rect 7984 19428 7990 19440
rect 8772 19428 8800 19459
rect 9674 19428 9680 19440
rect 7984 19400 8708 19428
rect 8772 19400 9680 19428
rect 7984 19388 7990 19400
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19360 1455 19363
rect 6914 19360 6920 19372
rect 1443 19332 6920 19360
rect 1443 19329 1455 19332
rect 1397 19323 1455 19329
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 8294 19360 8300 19372
rect 8255 19332 8300 19360
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 8680 19360 8708 19400
rect 9674 19388 9680 19400
rect 9732 19388 9738 19440
rect 8941 19363 8999 19369
rect 8941 19360 8953 19363
rect 8680 19332 8953 19360
rect 8941 19329 8953 19332
rect 8987 19329 8999 19363
rect 8941 19323 8999 19329
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9784 19369 9812 19468
rect 9950 19428 9956 19440
rect 9911 19400 9956 19428
rect 9950 19388 9956 19400
rect 10008 19388 10014 19440
rect 10045 19431 10103 19437
rect 10045 19397 10057 19431
rect 10091 19428 10103 19431
rect 10318 19428 10324 19440
rect 10091 19400 10324 19428
rect 10091 19397 10103 19400
rect 10045 19391 10103 19397
rect 10318 19388 10324 19400
rect 10376 19388 10382 19440
rect 9309 19363 9367 19369
rect 9309 19360 9321 19363
rect 9088 19332 9321 19360
rect 9088 19320 9094 19332
rect 9309 19329 9321 19332
rect 9355 19329 9367 19363
rect 9309 19323 9367 19329
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 9858 19360 9864 19372
rect 9815 19332 9864 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 10502 19360 10508 19372
rect 9968 19332 10508 19360
rect 9968 19292 9996 19332
rect 10502 19320 10508 19332
rect 10560 19320 10566 19372
rect 9508 19264 9996 19292
rect 9508 19233 9536 19264
rect 9493 19227 9551 19233
rect 9493 19193 9505 19227
rect 9539 19193 9551 19227
rect 9493 19187 9551 19193
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 1104 19066 10856 19088
rect 1104 19014 2582 19066
rect 2634 19014 2646 19066
rect 2698 19014 2710 19066
rect 2762 19014 2774 19066
rect 2826 19014 2838 19066
rect 2890 19014 5845 19066
rect 5897 19014 5909 19066
rect 5961 19014 5973 19066
rect 6025 19014 6037 19066
rect 6089 19014 6101 19066
rect 6153 19014 9109 19066
rect 9161 19014 9173 19066
rect 9225 19014 9237 19066
rect 9289 19014 9301 19066
rect 9353 19014 9365 19066
rect 9417 19014 10856 19066
rect 1104 18992 10856 19014
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 7561 18955 7619 18961
rect 7561 18952 7573 18955
rect 7340 18924 7573 18952
rect 7340 18912 7346 18924
rect 7561 18921 7573 18924
rect 7607 18921 7619 18955
rect 7561 18915 7619 18921
rect 8205 18955 8263 18961
rect 8205 18921 8217 18955
rect 8251 18952 8263 18955
rect 9766 18952 9772 18964
rect 8251 18924 9772 18952
rect 8251 18921 8263 18924
rect 8205 18915 8263 18921
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 10226 18952 10232 18964
rect 10187 18924 10232 18952
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10318 18816 10324 18828
rect 10091 18788 10324 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18748 7803 18751
rect 7834 18748 7840 18760
rect 7791 18720 7840 18748
rect 7791 18717 7803 18720
rect 7745 18711 7803 18717
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 8662 18748 8668 18760
rect 8435 18720 8668 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18748 9367 18751
rect 10413 18751 10471 18757
rect 9355 18720 9904 18748
rect 9355 18717 9367 18720
rect 9309 18711 9367 18717
rect 9876 18689 9904 18720
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 10459 18720 11161 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 9861 18683 9919 18689
rect 2746 18652 9444 18680
rect 1394 18572 1400 18624
rect 1452 18612 1458 18624
rect 2746 18612 2774 18652
rect 9416 18621 9444 18652
rect 9861 18649 9873 18683
rect 9907 18680 9919 18683
rect 11609 18683 11667 18689
rect 11609 18680 11621 18683
rect 9907 18652 11621 18680
rect 9907 18649 9919 18652
rect 9861 18643 9919 18649
rect 11609 18649 11621 18652
rect 11655 18649 11667 18683
rect 11609 18643 11667 18649
rect 1452 18584 2774 18612
rect 9401 18615 9459 18621
rect 1452 18572 1458 18584
rect 9401 18581 9413 18615
rect 9447 18581 9459 18615
rect 9401 18575 9459 18581
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 9769 18615 9827 18621
rect 9769 18612 9781 18615
rect 9732 18584 9781 18612
rect 9732 18572 9738 18584
rect 9769 18581 9781 18584
rect 9815 18581 9827 18615
rect 9769 18575 9827 18581
rect 1104 18522 10856 18544
rect 1104 18470 4213 18522
rect 4265 18470 4277 18522
rect 4329 18470 4341 18522
rect 4393 18470 4405 18522
rect 4457 18470 4469 18522
rect 4521 18470 7477 18522
rect 7529 18470 7541 18522
rect 7593 18470 7605 18522
rect 7657 18470 7669 18522
rect 7721 18470 7733 18522
rect 7785 18470 10856 18522
rect 1104 18448 10856 18470
rect 7098 18408 7104 18420
rect 7059 18380 7104 18408
rect 7098 18368 7104 18380
rect 7156 18368 7162 18420
rect 8846 18368 8852 18420
rect 8904 18408 8910 18420
rect 9217 18411 9275 18417
rect 9217 18408 9229 18411
rect 8904 18380 9229 18408
rect 8904 18368 8910 18380
rect 9217 18377 9229 18380
rect 9263 18408 9275 18411
rect 9582 18408 9588 18420
rect 9263 18380 9588 18408
rect 9263 18377 9275 18380
rect 9217 18371 9275 18377
rect 9582 18368 9588 18380
rect 9640 18408 9646 18420
rect 10229 18411 10287 18417
rect 10229 18408 10241 18411
rect 9640 18380 10241 18408
rect 9640 18368 9646 18380
rect 10229 18377 10241 18380
rect 10275 18377 10287 18411
rect 10229 18371 10287 18377
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 7282 18272 7288 18284
rect 7243 18244 7288 18272
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 8386 18272 8392 18284
rect 8347 18244 8392 18272
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 1578 18136 1584 18148
rect 1539 18108 1584 18136
rect 1578 18096 1584 18108
rect 1636 18096 1642 18148
rect 7834 18028 7840 18080
rect 7892 18068 7898 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 7892 18040 8217 18068
rect 7892 18028 7898 18040
rect 8205 18037 8217 18040
rect 8251 18037 8263 18071
rect 8205 18031 8263 18037
rect 1104 17978 10856 18000
rect 1104 17926 2582 17978
rect 2634 17926 2646 17978
rect 2698 17926 2710 17978
rect 2762 17926 2774 17978
rect 2826 17926 2838 17978
rect 2890 17926 5845 17978
rect 5897 17926 5909 17978
rect 5961 17926 5973 17978
rect 6025 17926 6037 17978
rect 6089 17926 6101 17978
rect 6153 17926 9109 17978
rect 9161 17926 9173 17978
rect 9225 17926 9237 17978
rect 9289 17926 9301 17978
rect 9353 17926 9365 17978
rect 9417 17926 10856 17978
rect 1104 17904 10856 17926
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 9030 17864 9036 17876
rect 8435 17836 9036 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 5350 17756 5356 17808
rect 5408 17796 5414 17808
rect 5408 17768 9720 17796
rect 5408 17756 5414 17768
rect 5626 17728 5632 17740
rect 1412 17700 5632 17728
rect 1412 17669 1440 17700
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 2958 17620 2964 17672
rect 3016 17660 3022 17672
rect 6549 17663 6607 17669
rect 6549 17660 6561 17663
rect 3016 17632 6561 17660
rect 3016 17620 3022 17632
rect 6549 17629 6561 17632
rect 6595 17660 6607 17663
rect 7006 17660 7012 17672
rect 6595 17632 7012 17660
rect 6595 17629 6607 17632
rect 6549 17623 6607 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 7745 17663 7803 17669
rect 7745 17660 7757 17663
rect 7432 17632 7757 17660
rect 7432 17620 7438 17632
rect 7745 17629 7757 17632
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 8230 17595 8288 17601
rect 8230 17561 8242 17595
rect 8276 17592 8288 17595
rect 9122 17592 9128 17604
rect 8276 17564 9128 17592
rect 8276 17561 8288 17564
rect 8230 17555 8288 17561
rect 9122 17552 9128 17564
rect 9180 17552 9186 17604
rect 9692 17592 9720 17768
rect 9858 17728 9864 17740
rect 9819 17700 9864 17728
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10318 17728 10324 17740
rect 10091 17700 10324 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 9692 17564 9904 17592
rect 9876 17536 9904 17564
rect 1578 17524 1584 17536
rect 1539 17496 1584 17524
rect 1578 17484 1584 17496
rect 1636 17484 1642 17536
rect 6454 17484 6460 17536
rect 6512 17524 6518 17536
rect 6641 17527 6699 17533
rect 6641 17524 6653 17527
rect 6512 17496 6653 17524
rect 6512 17484 6518 17496
rect 6641 17493 6653 17496
rect 6687 17493 6699 17527
rect 8018 17524 8024 17536
rect 7979 17496 8024 17524
rect 6641 17487 6699 17493
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8168 17496 8213 17524
rect 8168 17484 8174 17496
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 9401 17527 9459 17533
rect 9401 17524 9413 17527
rect 8812 17496 9413 17524
rect 8812 17484 8818 17496
rect 9401 17493 9413 17496
rect 9447 17493 9459 17527
rect 9766 17524 9772 17536
rect 9727 17496 9772 17524
rect 9401 17487 9459 17493
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 9858 17484 9864 17536
rect 9916 17484 9922 17536
rect 1104 17434 10856 17456
rect 1104 17382 4213 17434
rect 4265 17382 4277 17434
rect 4329 17382 4341 17434
rect 4393 17382 4405 17434
rect 4457 17382 4469 17434
rect 4521 17382 7477 17434
rect 7529 17382 7541 17434
rect 7593 17382 7605 17434
rect 7657 17382 7669 17434
rect 7721 17382 7733 17434
rect 7785 17382 10856 17434
rect 1104 17360 10856 17382
rect 11333 17391 11391 17397
rect 11333 17357 11345 17391
rect 11379 17388 11391 17391
rect 11609 17391 11667 17397
rect 11609 17388 11621 17391
rect 11379 17360 11621 17388
rect 11379 17357 11391 17360
rect 11333 17351 11391 17357
rect 11609 17357 11621 17360
rect 11655 17357 11667 17391
rect 11609 17351 11667 17357
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9401 17323 9459 17329
rect 9401 17320 9413 17323
rect 9263 17292 9413 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 9401 17289 9413 17292
rect 9447 17289 9459 17323
rect 9401 17283 9459 17289
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 9861 17323 9919 17329
rect 9861 17320 9873 17323
rect 9640 17292 9873 17320
rect 9640 17280 9646 17292
rect 9861 17289 9873 17292
rect 9907 17289 9919 17323
rect 9861 17283 9919 17289
rect 3970 17212 3976 17264
rect 4028 17252 4034 17264
rect 7650 17252 7656 17264
rect 4028 17224 7656 17252
rect 4028 17212 4034 17224
rect 7650 17212 7656 17224
rect 7708 17212 7714 17264
rect 7742 17212 7748 17264
rect 7800 17252 7806 17264
rect 10321 17255 10379 17261
rect 10321 17252 10333 17255
rect 7800 17224 10333 17252
rect 7800 17212 7806 17224
rect 10321 17221 10333 17224
rect 10367 17221 10379 17255
rect 10321 17215 10379 17221
rect 11333 17255 11391 17261
rect 11333 17221 11345 17255
rect 11379 17252 11391 17255
rect 11701 17255 11759 17261
rect 11701 17252 11713 17255
rect 11379 17224 11713 17252
rect 11379 17221 11391 17224
rect 11333 17215 11391 17221
rect 11701 17221 11713 17224
rect 11747 17221 11759 17255
rect 11701 17215 11759 17221
rect 1397 17187 1455 17193
rect 1397 17153 1409 17187
rect 1443 17184 1455 17187
rect 6178 17184 6184 17196
rect 1443 17156 6184 17184
rect 1443 17153 1455 17156
rect 1397 17147 1455 17153
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 6454 17184 6460 17196
rect 6415 17156 6460 17184
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6656 17156 7113 17184
rect 6656 17057 6684 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 8001 17187 8059 17193
rect 8001 17184 8013 17187
rect 7248 17156 8013 17184
rect 7248 17144 7254 17156
rect 8001 17153 8013 17156
rect 8047 17153 8059 17187
rect 8001 17147 8059 17153
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8352 17156 9229 17184
rect 8352 17144 8358 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 9769 17187 9827 17193
rect 9769 17153 9781 17187
rect 9815 17153 9827 17187
rect 10226 17184 10232 17196
rect 10187 17156 10232 17184
rect 9769 17147 9827 17153
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7300 17088 7757 17116
rect 7300 17057 7328 17088
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17017 6699 17051
rect 6641 17011 6699 17017
rect 7285 17051 7343 17057
rect 7285 17017 7297 17051
rect 7331 17017 7343 17051
rect 9784 17048 9812 17147
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 10318 17116 10324 17128
rect 10091 17088 10324 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 11287 17088 11621 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 11609 17085 11621 17088
rect 11655 17085 11667 17119
rect 11609 17079 11667 17085
rect 7285 17011 7343 17017
rect 8680 17020 9812 17048
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 6270 16940 6276 16992
rect 6328 16980 6334 16992
rect 8680 16980 8708 17020
rect 6328 16952 8708 16980
rect 6328 16940 6334 16952
rect 1104 16890 10856 16912
rect 1104 16838 2582 16890
rect 2634 16838 2646 16890
rect 2698 16838 2710 16890
rect 2762 16838 2774 16890
rect 2826 16838 2838 16890
rect 2890 16838 5845 16890
rect 5897 16838 5909 16890
rect 5961 16838 5973 16890
rect 6025 16838 6037 16890
rect 6089 16838 6101 16890
rect 6153 16838 9109 16890
rect 9161 16838 9173 16890
rect 9225 16838 9237 16890
rect 9289 16838 9301 16890
rect 9353 16838 9365 16890
rect 9417 16838 10856 16890
rect 1104 16816 10856 16838
rect 6457 16779 6515 16785
rect 6457 16745 6469 16779
rect 6503 16776 6515 16779
rect 7190 16776 7196 16788
rect 6503 16748 7196 16776
rect 6503 16745 6515 16748
rect 6457 16739 6515 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 9950 16776 9956 16788
rect 7708 16748 9956 16776
rect 7708 16736 7714 16748
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 6656 16680 7420 16708
rect 6656 16581 6684 16680
rect 7392 16652 7420 16680
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 7064 16612 7144 16640
rect 7064 16600 7070 16612
rect 7116 16581 7144 16612
rect 7374 16600 7380 16652
rect 7432 16640 7438 16652
rect 7745 16643 7803 16649
rect 7745 16640 7757 16643
rect 7432 16612 7757 16640
rect 7432 16600 7438 16612
rect 7745 16609 7757 16612
rect 7791 16640 7803 16643
rect 7926 16640 7932 16652
rect 7791 16612 7932 16640
rect 7791 16609 7803 16612
rect 7745 16603 7803 16609
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 9585 16643 9643 16649
rect 9585 16640 9597 16643
rect 8536 16612 9597 16640
rect 8536 16600 8542 16612
rect 9585 16609 9597 16612
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 10318 16640 10324 16652
rect 9815 16612 10324 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16541 6515 16575
rect 6457 16535 6515 16541
rect 6641 16575 6699 16581
rect 6641 16541 6653 16575
rect 6687 16541 6699 16575
rect 6641 16535 6699 16541
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 8128 16572 8156 16600
rect 8128 16544 9168 16572
rect 7101 16535 7159 16541
rect 1412 16504 1440 16535
rect 6472 16504 6500 16535
rect 7742 16504 7748 16516
rect 1412 16476 2774 16504
rect 6472 16476 7748 16504
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 2746 16436 2774 16476
rect 7742 16464 7748 16476
rect 7800 16504 7806 16516
rect 8110 16504 8116 16516
rect 7800 16476 8116 16504
rect 7800 16464 7806 16476
rect 8110 16464 8116 16476
rect 8168 16504 8174 16516
rect 8230 16507 8288 16513
rect 8230 16504 8242 16507
rect 8168 16476 8242 16504
rect 8168 16464 8174 16476
rect 8230 16473 8242 16476
rect 8276 16473 8288 16507
rect 8230 16467 8288 16473
rect 6914 16436 6920 16448
rect 2746 16408 6920 16436
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7190 16436 7196 16448
rect 7151 16408 7196 16436
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 8386 16436 8392 16448
rect 8347 16408 8392 16436
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 9140 16445 9168 16544
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 9493 16575 9551 16581
rect 9493 16572 9505 16575
rect 9272 16544 9505 16572
rect 9272 16532 9278 16544
rect 9493 16541 9505 16544
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 11241 16575 11299 16581
rect 11241 16541 11253 16575
rect 11287 16572 11299 16575
rect 11606 16572 11612 16584
rect 11287 16544 11612 16572
rect 11287 16541 11299 16544
rect 11241 16535 11299 16541
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16405 9183 16439
rect 9125 16399 9183 16405
rect 1104 16346 10856 16368
rect 1104 16294 4213 16346
rect 4265 16294 4277 16346
rect 4329 16294 4341 16346
rect 4393 16294 4405 16346
rect 4457 16294 4469 16346
rect 4521 16294 7477 16346
rect 7529 16294 7541 16346
rect 7593 16294 7605 16346
rect 7657 16294 7669 16346
rect 7721 16294 7733 16346
rect 7785 16294 10856 16346
rect 1104 16272 10856 16294
rect 11054 16260 11060 16312
rect 11112 16300 11118 16312
rect 11149 16303 11207 16309
rect 11149 16300 11161 16303
rect 11112 16272 11161 16300
rect 11112 16260 11118 16272
rect 11149 16269 11161 16272
rect 11195 16269 11207 16303
rect 11149 16263 11207 16269
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 8941 16235 8999 16241
rect 5675 16204 7972 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 7834 16173 7840 16176
rect 7828 16164 7840 16173
rect 7795 16136 7840 16164
rect 7828 16127 7840 16136
rect 7834 16124 7840 16127
rect 7892 16124 7898 16176
rect 7944 16164 7972 16204
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 10226 16232 10232 16244
rect 8987 16204 10232 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 9674 16164 9680 16176
rect 7944 16136 9680 16164
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 9769 16167 9827 16173
rect 9769 16133 9781 16167
rect 9815 16164 9827 16167
rect 11149 16167 11207 16173
rect 11149 16164 11161 16167
rect 9815 16136 11161 16164
rect 9815 16133 9827 16136
rect 9769 16127 9827 16133
rect 11149 16133 11161 16136
rect 11195 16164 11207 16167
rect 11882 16164 11888 16176
rect 11195 16136 11888 16164
rect 11195 16133 11207 16136
rect 11149 16127 11207 16133
rect 11882 16124 11888 16136
rect 11940 16124 11946 16176
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6914 16096 6920 16108
rect 5859 16068 6920 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7098 16096 7104 16108
rect 7059 16068 7104 16096
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7561 16099 7619 16105
rect 7561 16096 7573 16099
rect 7248 16068 7573 16096
rect 7248 16056 7254 16068
rect 7561 16065 7573 16068
rect 7607 16065 7619 16099
rect 7561 16059 7619 16065
rect 7668 16068 8616 16096
rect 6730 15988 6736 16040
rect 6788 16028 6794 16040
rect 7668 16028 7696 16068
rect 6788 16000 7696 16028
rect 6788 15988 6794 16000
rect 8588 15960 8616 16068
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 9861 16031 9919 16037
rect 9861 16028 9873 16031
rect 9640 16000 9873 16028
rect 9640 15988 9646 16000
rect 9861 15997 9873 16000
rect 9907 15997 9919 16031
rect 9861 15991 9919 15997
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 16028 10011 16031
rect 10318 16028 10324 16040
rect 9999 16000 10324 16028
rect 9999 15997 10011 16000
rect 9953 15991 10011 15997
rect 10318 15988 10324 16000
rect 10376 15988 10382 16040
rect 10042 15960 10048 15972
rect 8588 15932 10048 15960
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 474 15852 480 15904
rect 532 15892 538 15904
rect 5350 15892 5356 15904
rect 532 15864 5356 15892
rect 532 15852 538 15864
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 6917 15895 6975 15901
rect 6917 15861 6929 15895
rect 6963 15892 6975 15895
rect 7282 15892 7288 15904
rect 6963 15864 7288 15892
rect 6963 15861 6975 15864
rect 6917 15855 6975 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 7984 15864 9413 15892
rect 7984 15852 7990 15864
rect 9401 15861 9413 15864
rect 9447 15861 9459 15895
rect 9401 15855 9459 15861
rect 1104 15802 10856 15824
rect 1104 15750 2582 15802
rect 2634 15750 2646 15802
rect 2698 15750 2710 15802
rect 2762 15750 2774 15802
rect 2826 15750 2838 15802
rect 2890 15750 5845 15802
rect 5897 15750 5909 15802
rect 5961 15750 5973 15802
rect 6025 15750 6037 15802
rect 6089 15750 6101 15802
rect 6153 15750 9109 15802
rect 9161 15750 9173 15802
rect 9225 15750 9237 15802
rect 9289 15750 9301 15802
rect 9353 15750 9365 15802
rect 9417 15750 10856 15802
rect 1104 15728 10856 15750
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 8113 15691 8171 15697
rect 8113 15688 8125 15691
rect 5408 15660 8125 15688
rect 5408 15648 5414 15660
rect 8113 15657 8125 15660
rect 8159 15657 8171 15691
rect 8113 15651 8171 15657
rect 8294 15620 8300 15632
rect 2746 15592 8300 15620
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15453 1455 15487
rect 1397 15447 1455 15453
rect 1412 15416 1440 15447
rect 2746 15416 2774 15592
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 10134 15620 10140 15632
rect 8772 15592 10140 15620
rect 7190 15552 7196 15564
rect 6748 15524 7196 15552
rect 6748 15493 6776 15524
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 8772 15552 8800 15592
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 7340 15524 8800 15552
rect 9309 15555 9367 15561
rect 7340 15512 7346 15524
rect 9309 15521 9321 15555
rect 9355 15552 9367 15555
rect 10045 15555 10103 15561
rect 9355 15524 9904 15552
rect 9355 15521 9367 15524
rect 9309 15515 9367 15521
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15453 6791 15487
rect 6733 15447 6791 15453
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 6880 15456 7389 15484
rect 6880 15444 6886 15456
rect 7377 15453 7389 15456
rect 7423 15453 7435 15487
rect 7377 15447 7435 15453
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15484 8079 15487
rect 8110 15484 8116 15496
rect 8067 15456 8116 15484
rect 8067 15453 8079 15456
rect 8021 15447 8079 15453
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 9398 15484 9404 15496
rect 8352 15456 9404 15484
rect 8352 15444 8358 15456
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 9876 15493 9904 15524
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 10318 15552 10324 15564
rect 10091 15524 10324 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15484 9919 15487
rect 11241 15487 11299 15493
rect 11241 15484 11253 15487
rect 9907 15456 11253 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 11241 15453 11253 15456
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 1412 15388 2774 15416
rect 6638 15376 6644 15428
rect 6696 15416 6702 15428
rect 7837 15419 7895 15425
rect 7837 15416 7849 15419
rect 6696 15388 7849 15416
rect 6696 15376 6702 15388
rect 7837 15385 7849 15388
rect 7883 15385 7895 15419
rect 9784 15416 9812 15444
rect 7837 15379 7895 15385
rect 8588 15388 9812 15416
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 6730 15348 6736 15360
rect 6595 15320 6736 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 7193 15351 7251 15357
rect 7193 15317 7205 15351
rect 7239 15348 7251 15351
rect 8588 15348 8616 15388
rect 7239 15320 8616 15348
rect 7239 15317 7251 15320
rect 7193 15311 7251 15317
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 8938 15348 8944 15360
rect 8720 15320 8944 15348
rect 8720 15308 8726 15320
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 9398 15348 9404 15360
rect 9359 15320 9404 15348
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 9766 15348 9772 15360
rect 9727 15320 9772 15348
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 1104 15258 10856 15280
rect 1104 15206 4213 15258
rect 4265 15206 4277 15258
rect 4329 15206 4341 15258
rect 4393 15206 4405 15258
rect 4457 15206 4469 15258
rect 4521 15206 7477 15258
rect 7529 15206 7541 15258
rect 7593 15206 7605 15258
rect 7657 15206 7669 15258
rect 7721 15206 7733 15258
rect 7785 15206 10856 15258
rect 1104 15184 10856 15206
rect 6825 15147 6883 15153
rect 6825 15113 6837 15147
rect 6871 15144 6883 15147
rect 7926 15144 7932 15156
rect 6871 15116 7932 15144
rect 6871 15113 6883 15116
rect 6825 15107 6883 15113
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8662 15144 8668 15156
rect 8623 15116 8668 15144
rect 8662 15104 8668 15116
rect 8720 15104 8726 15156
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 9766 15144 9772 15156
rect 8904 15116 9772 15144
rect 8904 15104 8910 15116
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 9861 15147 9919 15153
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 11514 15144 11520 15156
rect 9907 15116 11520 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 8294 15076 8300 15088
rect 1412 15048 8300 15076
rect 1412 15017 1440 15048
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 8573 15079 8631 15085
rect 8573 15045 8585 15079
rect 8619 15045 8631 15079
rect 9876 15076 9904 15107
rect 11514 15104 11520 15116
rect 11572 15104 11578 15156
rect 8573 15039 8631 15045
rect 9692 15048 9904 15076
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 15008 7067 15011
rect 7466 15008 7472 15020
rect 7055 14980 7472 15008
rect 7055 14977 7067 14980
rect 7009 14971 7067 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 15008 7619 15011
rect 8478 15008 8484 15020
rect 7607 14980 8484 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 5684 14912 8340 14940
rect 5684 14900 5690 14912
rect 7745 14875 7803 14881
rect 7745 14841 7757 14875
rect 7791 14872 7803 14875
rect 7834 14872 7840 14884
rect 7791 14844 7840 14872
rect 7791 14841 7803 14844
rect 7745 14835 7803 14841
rect 7834 14832 7840 14844
rect 7892 14832 7898 14884
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7374 14804 7380 14816
rect 7156 14776 7380 14804
rect 7156 14764 7162 14776
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 7708 14776 8217 14804
rect 7708 14764 7714 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8312 14804 8340 14912
rect 8386 14900 8392 14952
rect 8444 14940 8450 14952
rect 8588 14940 8616 15039
rect 9030 15008 9036 15020
rect 8772 14980 9036 15008
rect 8772 14949 8800 14980
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 9309 15011 9367 15017
rect 9309 14977 9321 15011
rect 9355 15008 9367 15011
rect 9692 15008 9720 15048
rect 9355 14980 9720 15008
rect 9769 15011 9827 15017
rect 9355 14977 9367 14980
rect 9309 14971 9367 14977
rect 9769 14977 9781 15011
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 8444 14912 8616 14940
rect 8757 14943 8815 14949
rect 8444 14900 8450 14912
rect 8757 14909 8769 14943
rect 8803 14909 8815 14943
rect 9784 14940 9812 14971
rect 8757 14903 8815 14909
rect 8864 14912 9812 14940
rect 9953 14943 10011 14949
rect 8864 14804 8892 14912
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 10318 14940 10324 14952
rect 9999 14912 10324 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 8312 14776 8892 14804
rect 8205 14767 8263 14773
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9401 14807 9459 14813
rect 9401 14804 9413 14807
rect 8996 14776 9413 14804
rect 8996 14764 9002 14776
rect 9401 14773 9413 14776
rect 9447 14773 9459 14807
rect 9401 14767 9459 14773
rect 1104 14714 10856 14736
rect 1104 14662 2582 14714
rect 2634 14662 2646 14714
rect 2698 14662 2710 14714
rect 2762 14662 2774 14714
rect 2826 14662 2838 14714
rect 2890 14662 5845 14714
rect 5897 14662 5909 14714
rect 5961 14662 5973 14714
rect 6025 14662 6037 14714
rect 6089 14662 6101 14714
rect 6153 14662 9109 14714
rect 9161 14662 9173 14714
rect 9225 14662 9237 14714
rect 9289 14662 9301 14714
rect 9353 14662 9365 14714
rect 9417 14662 10856 14714
rect 1104 14640 10856 14662
rect 8938 14600 8944 14612
rect 2746 14572 8944 14600
rect 2746 14532 2774 14572
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 5258 14532 5264 14544
rect 1412 14504 2774 14532
rect 5219 14504 5264 14532
rect 1412 14405 1440 14504
rect 5258 14492 5264 14504
rect 5316 14492 5322 14544
rect 6914 14532 6920 14544
rect 5460 14504 6920 14532
rect 5460 14405 5488 14504
rect 6914 14492 6920 14504
rect 6972 14492 6978 14544
rect 7208 14504 7696 14532
rect 7208 14464 7236 14504
rect 6656 14436 7236 14464
rect 6656 14405 6684 14436
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 7668 14464 7696 14504
rect 7742 14492 7748 14544
rect 7800 14532 7806 14544
rect 8110 14532 8116 14544
rect 7800 14504 8116 14532
rect 7800 14492 7806 14504
rect 8110 14492 8116 14504
rect 8168 14492 8174 14544
rect 8938 14464 8944 14476
rect 7340 14436 7385 14464
rect 7668 14436 8944 14464
rect 7340 14424 7346 14436
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 9858 14464 9864 14476
rect 9819 14436 9864 14464
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 9953 14467 10011 14473
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 10318 14464 10324 14476
rect 9999 14436 10324 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6914 14396 6920 14408
rect 6641 14359 6699 14365
rect 6748 14368 6920 14396
rect 6104 14328 6132 14359
rect 6748 14328 6776 14368
rect 6914 14356 6920 14368
rect 6972 14356 6978 14408
rect 7650 14396 7656 14408
rect 7611 14368 7656 14396
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 7770 14399 7828 14405
rect 7770 14365 7782 14399
rect 7816 14396 7828 14399
rect 7926 14396 7932 14408
rect 7816 14368 7932 14396
rect 7816 14365 7828 14368
rect 7770 14359 7828 14365
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 9968 14396 9996 14427
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 9180 14368 9996 14396
rect 9180 14356 9186 14368
rect 6104 14300 6776 14328
rect 6825 14331 6883 14337
rect 6825 14297 6837 14331
rect 6871 14328 6883 14331
rect 7374 14328 7380 14340
rect 6871 14300 7380 14328
rect 6871 14297 6883 14300
rect 6825 14291 6883 14297
rect 7374 14288 7380 14300
rect 7432 14288 7438 14340
rect 8294 14288 8300 14340
rect 8352 14328 8358 14340
rect 9769 14331 9827 14337
rect 9769 14328 9781 14331
rect 8352 14300 9781 14328
rect 8352 14288 8358 14300
rect 9769 14297 9781 14300
rect 9815 14297 9827 14331
rect 9769 14291 9827 14297
rect 1578 14260 1584 14272
rect 1539 14232 1584 14260
rect 1578 14220 1584 14232
rect 1636 14220 1642 14272
rect 5905 14263 5963 14269
rect 5905 14229 5917 14263
rect 5951 14260 5963 14263
rect 6270 14260 6276 14272
rect 5951 14232 6276 14260
rect 5951 14229 5963 14232
rect 5905 14223 5963 14229
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 7561 14263 7619 14269
rect 7561 14260 7573 14263
rect 7340 14232 7573 14260
rect 7340 14220 7346 14232
rect 7561 14229 7573 14232
rect 7607 14229 7619 14263
rect 7561 14223 7619 14229
rect 7929 14263 7987 14269
rect 7929 14229 7941 14263
rect 7975 14260 7987 14263
rect 8846 14260 8852 14272
rect 7975 14232 8852 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9398 14260 9404 14272
rect 9359 14232 9404 14260
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 1104 14170 10856 14192
rect 1104 14118 4213 14170
rect 4265 14118 4277 14170
rect 4329 14118 4341 14170
rect 4393 14118 4405 14170
rect 4457 14118 4469 14170
rect 4521 14118 7477 14170
rect 7529 14118 7541 14170
rect 7593 14118 7605 14170
rect 7657 14118 7669 14170
rect 7721 14118 7733 14170
rect 7785 14118 10856 14170
rect 1104 14096 10856 14118
rect 5626 14056 5632 14068
rect 5587 14028 5632 14056
rect 5626 14016 5632 14028
rect 5684 14016 5690 14068
rect 6362 14056 6368 14068
rect 6323 14028 6368 14056
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 7469 14059 7527 14065
rect 7469 14056 7481 14059
rect 7156 14028 7481 14056
rect 7156 14016 7162 14028
rect 7469 14025 7481 14028
rect 7515 14025 7527 14059
rect 7469 14019 7527 14025
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 8076 14028 8217 14056
rect 8076 14016 8082 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8205 14019 8263 14025
rect 8386 14016 8392 14068
rect 8444 14056 8450 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8444 14028 8585 14056
rect 8444 14016 8450 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 8573 14019 8631 14025
rect 9861 14059 9919 14065
rect 9861 14025 9873 14059
rect 9907 14056 9919 14059
rect 9950 14056 9956 14068
rect 9907 14028 9956 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 7650 13948 7656 14000
rect 7708 13988 7714 14000
rect 9398 13988 9404 14000
rect 7708 13960 9404 13988
rect 7708 13948 7714 13960
rect 9398 13948 9404 13960
rect 9456 13948 9462 14000
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 6549 13924 6607 13929
rect 6730 13924 6736 13932
rect 6549 13923 6736 13924
rect 6549 13889 6561 13923
rect 6595 13896 6736 13923
rect 6595 13889 6607 13896
rect 6549 13883 6607 13889
rect 1412 13784 1440 13883
rect 5828 13852 5856 13883
rect 6730 13880 6736 13896
rect 6788 13880 6794 13932
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 8665 13923 8723 13929
rect 7423 13892 8432 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7190 13852 7196 13864
rect 5828 13824 7196 13852
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 8404 13852 8432 13892
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 9030 13920 9036 13932
rect 8711 13892 9036 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 8680 13852 8708 13883
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9732 13892 9781 13920
rect 9732 13880 9738 13892
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 7616 13824 7788 13852
rect 8404 13824 8708 13852
rect 8849 13855 8907 13861
rect 7616 13812 7622 13824
rect 7650 13784 7656 13796
rect 1412 13756 7656 13784
rect 7650 13744 7656 13756
rect 7708 13744 7714 13796
rect 7760 13784 7788 13824
rect 8849 13821 8861 13855
rect 8895 13852 8907 13855
rect 9122 13852 9128 13864
rect 8895 13824 9128 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 8864 13784 8892 13815
rect 9122 13812 9128 13824
rect 9180 13852 9186 13864
rect 9950 13852 9956 13864
rect 9180 13824 9956 13852
rect 9180 13812 9186 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 7760 13756 8892 13784
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 7009 13719 7067 13725
rect 7009 13716 7021 13719
rect 5684 13688 7021 13716
rect 5684 13676 5690 13688
rect 7009 13685 7021 13688
rect 7055 13716 7067 13719
rect 7282 13716 7288 13728
rect 7055 13688 7288 13716
rect 7055 13685 7067 13688
rect 7009 13679 7067 13685
rect 7282 13676 7288 13688
rect 7340 13676 7346 13728
rect 8294 13676 8300 13728
rect 8352 13716 8358 13728
rect 9401 13719 9459 13725
rect 9401 13716 9413 13719
rect 8352 13688 9413 13716
rect 8352 13676 8358 13688
rect 9401 13685 9413 13688
rect 9447 13685 9459 13719
rect 9401 13679 9459 13685
rect 1104 13626 10856 13648
rect 1104 13574 2582 13626
rect 2634 13574 2646 13626
rect 2698 13574 2710 13626
rect 2762 13574 2774 13626
rect 2826 13574 2838 13626
rect 2890 13574 5845 13626
rect 5897 13574 5909 13626
rect 5961 13574 5973 13626
rect 6025 13574 6037 13626
rect 6089 13574 6101 13626
rect 6153 13574 9109 13626
rect 9161 13574 9173 13626
rect 9225 13574 9237 13626
rect 9289 13574 9301 13626
rect 9353 13574 9365 13626
rect 9417 13574 10856 13626
rect 1104 13552 10856 13574
rect 5997 13515 6055 13521
rect 5997 13481 6009 13515
rect 6043 13512 6055 13515
rect 6822 13512 6828 13524
rect 6043 13484 6828 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7650 13512 7656 13524
rect 7611 13484 7656 13512
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 8294 13444 8300 13456
rect 1412 13416 8300 13444
rect 1412 13317 1440 13416
rect 8294 13404 8300 13416
rect 8352 13404 8358 13456
rect 9582 13444 9588 13456
rect 8956 13416 9588 13444
rect 5350 13376 5356 13388
rect 5311 13348 5356 13376
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 5626 13376 5632 13388
rect 5587 13348 5632 13376
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7558 13376 7564 13388
rect 7147 13348 7564 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7558 13336 7564 13348
rect 7616 13376 7622 13388
rect 8205 13379 8263 13385
rect 8205 13376 8217 13379
rect 7616 13348 8217 13376
rect 7616 13336 7622 13348
rect 8205 13345 8217 13348
rect 8251 13345 8263 13379
rect 8205 13339 8263 13345
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13308 5779 13311
rect 6086 13308 6092 13320
rect 5767 13280 6092 13308
rect 5767 13277 5779 13280
rect 5721 13271 5779 13277
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6236 13280 6837 13308
rect 6236 13268 6242 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 8018 13308 8024 13320
rect 6825 13271 6883 13277
rect 7576 13280 8024 13308
rect 5838 13243 5896 13249
rect 5838 13209 5850 13243
rect 5884 13240 5896 13243
rect 5884 13212 6684 13240
rect 5884 13209 5896 13212
rect 5838 13203 5896 13209
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 6546 13172 6552 13184
rect 6503 13144 6552 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 6656 13172 6684 13212
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 6917 13243 6975 13249
rect 6917 13240 6929 13243
rect 6788 13212 6929 13240
rect 6788 13200 6794 13212
rect 6917 13209 6929 13212
rect 6963 13209 6975 13243
rect 6917 13203 6975 13209
rect 7576 13172 7604 13280
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8662 13240 8668 13252
rect 8036 13212 8668 13240
rect 8036 13181 8064 13212
rect 8662 13200 8668 13212
rect 8720 13240 8726 13252
rect 8956 13240 8984 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 11149 13447 11207 13453
rect 11149 13444 11161 13447
rect 9876 13416 11161 13444
rect 9876 13376 9904 13416
rect 11149 13413 11161 13416
rect 11195 13413 11207 13447
rect 11149 13407 11207 13413
rect 8720 13212 8984 13240
rect 9232 13348 9904 13376
rect 8720 13200 8726 13212
rect 6656 13144 7604 13172
rect 8021 13175 8079 13181
rect 8021 13141 8033 13175
rect 8067 13141 8079 13175
rect 8021 13135 8079 13141
rect 8113 13175 8171 13181
rect 8113 13141 8125 13175
rect 8159 13172 8171 13175
rect 9232 13172 9260 13348
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 10008 13348 10053 13376
rect 10008 13336 10014 13348
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9861 13311 9919 13317
rect 9861 13308 9873 13311
rect 9355 13280 9873 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9861 13277 9873 13280
rect 9907 13308 9919 13311
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 9907 13280 11897 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 8159 13144 9260 13172
rect 9401 13175 9459 13181
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 9401 13141 9413 13175
rect 9447 13172 9459 13175
rect 9490 13172 9496 13184
rect 9447 13144 9496 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 9766 13172 9772 13184
rect 9727 13144 9772 13172
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 1104 13082 10856 13104
rect 1104 13030 4213 13082
rect 4265 13030 4277 13082
rect 4329 13030 4341 13082
rect 4393 13030 4405 13082
rect 4457 13030 4469 13082
rect 4521 13030 7477 13082
rect 7529 13030 7541 13082
rect 7593 13030 7605 13082
rect 7657 13030 7669 13082
rect 7721 13030 7733 13082
rect 7785 13030 10856 13082
rect 1104 13008 10856 13030
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 7064 12940 7205 12968
rect 7064 12928 7070 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 7193 12931 7251 12937
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7561 12971 7619 12977
rect 7561 12968 7573 12971
rect 7432 12940 7573 12968
rect 7432 12928 7438 12940
rect 7561 12937 7573 12940
rect 7607 12937 7619 12971
rect 7561 12931 7619 12937
rect 7653 12971 7711 12977
rect 7653 12937 7665 12971
rect 7699 12968 7711 12971
rect 7834 12968 7840 12980
rect 7699 12940 7840 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 9582 12968 9588 12980
rect 8996 12940 9588 12968
rect 8996 12928 9002 12940
rect 9582 12928 9588 12940
rect 9640 12968 9646 12980
rect 9677 12971 9735 12977
rect 9677 12968 9689 12971
rect 9640 12940 9689 12968
rect 9640 12928 9646 12940
rect 9677 12937 9689 12940
rect 9723 12937 9735 12971
rect 9677 12931 9735 12937
rect 8202 12860 8208 12912
rect 8260 12900 8266 12912
rect 8389 12903 8447 12909
rect 8389 12900 8401 12903
rect 8260 12872 8401 12900
rect 8260 12860 8266 12872
rect 8389 12869 8401 12872
rect 8435 12869 8447 12903
rect 8389 12863 8447 12869
rect 8846 12860 8852 12912
rect 8904 12860 8910 12912
rect 5626 12832 5632 12844
rect 5587 12804 5632 12832
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12832 6607 12835
rect 7098 12832 7104 12844
rect 6595 12804 7104 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 7098 12792 7104 12804
rect 7156 12792 7162 12844
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 8864 12832 8892 12860
rect 7432 12804 8892 12832
rect 7432 12792 7438 12804
rect 8938 12792 8944 12844
rect 8996 12832 9002 12844
rect 9398 12832 9404 12844
rect 8996 12804 9404 12832
rect 8996 12792 9002 12804
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 8846 12764 8852 12776
rect 7883 12736 8852 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 5813 12699 5871 12705
rect 5813 12665 5825 12699
rect 5859 12696 5871 12699
rect 7006 12696 7012 12708
rect 5859 12668 7012 12696
rect 5859 12665 5871 12668
rect 5813 12659 5871 12665
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 6638 12628 6644 12640
rect 6599 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 1104 12538 10856 12560
rect 1104 12486 2582 12538
rect 2634 12486 2646 12538
rect 2698 12486 2710 12538
rect 2762 12486 2774 12538
rect 2826 12486 2838 12538
rect 2890 12486 5845 12538
rect 5897 12486 5909 12538
rect 5961 12486 5973 12538
rect 6025 12486 6037 12538
rect 6089 12486 6101 12538
rect 6153 12486 9109 12538
rect 9161 12486 9173 12538
rect 9225 12486 9237 12538
rect 9289 12486 9301 12538
rect 9353 12486 9365 12538
rect 9417 12486 10856 12538
rect 1104 12464 10856 12486
rect 934 12384 940 12436
rect 992 12424 998 12436
rect 6178 12424 6184 12436
rect 992 12396 6184 12424
rect 992 12384 998 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 6512 12396 7972 12424
rect 6512 12384 6518 12396
rect 5721 12359 5779 12365
rect 5721 12325 5733 12359
rect 5767 12356 5779 12359
rect 7944 12356 7972 12396
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 8076 12396 8401 12424
rect 8076 12384 8082 12396
rect 8389 12393 8401 12396
rect 8435 12393 8447 12427
rect 8389 12387 8447 12393
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 8904 12396 9996 12424
rect 8904 12384 8910 12396
rect 5767 12328 6868 12356
rect 7944 12328 9904 12356
rect 5767 12325 5779 12328
rect 5721 12319 5779 12325
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 5810 12220 5816 12232
rect 1443 12192 5816 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6362 12220 6368 12232
rect 5960 12192 6005 12220
rect 6323 12192 6368 12220
rect 5960 12180 5966 12192
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 6840 12220 6868 12328
rect 7006 12288 7012 12300
rect 6967 12260 7012 12288
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 9876 12297 9904 12328
rect 9968 12300 9996 12396
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10008 12260 10053 12288
rect 10008 12248 10014 12260
rect 9674 12220 9680 12232
rect 6604 12192 6649 12220
rect 6840 12192 9680 12220
rect 6604 12180 6610 12192
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 7254 12155 7312 12161
rect 7254 12152 7266 12155
rect 6656 12124 7266 12152
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 6457 12087 6515 12093
rect 6457 12053 6469 12087
rect 6503 12084 6515 12087
rect 6656 12084 6684 12124
rect 7254 12121 7266 12124
rect 7300 12121 7312 12155
rect 7254 12115 7312 12121
rect 8386 12112 8392 12164
rect 8444 12152 8450 12164
rect 9490 12152 9496 12164
rect 8444 12124 9496 12152
rect 8444 12112 8450 12124
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 9398 12084 9404 12096
rect 6503 12056 6684 12084
rect 9359 12056 9404 12084
rect 6503 12053 6515 12056
rect 6457 12047 6515 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 9769 12087 9827 12093
rect 9769 12084 9781 12087
rect 9732 12056 9781 12084
rect 9732 12044 9738 12056
rect 9769 12053 9781 12056
rect 9815 12053 9827 12087
rect 9769 12047 9827 12053
rect 1104 11994 10856 12016
rect 1104 11942 4213 11994
rect 4265 11942 4277 11994
rect 4329 11942 4341 11994
rect 4393 11942 4405 11994
rect 4457 11942 4469 11994
rect 4521 11942 7477 11994
rect 7529 11942 7541 11994
rect 7593 11942 7605 11994
rect 7657 11942 7669 11994
rect 7721 11942 7733 11994
rect 7785 11942 10856 11994
rect 1104 11920 10856 11942
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 8386 11880 8392 11892
rect 5868 11852 8392 11880
rect 5868 11840 5874 11852
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 9677 11883 9735 11889
rect 9677 11880 9689 11883
rect 8536 11852 9689 11880
rect 8536 11840 8542 11852
rect 9677 11849 9689 11852
rect 9723 11849 9735 11883
rect 9677 11843 9735 11849
rect 9398 11812 9404 11824
rect 1412 11784 9404 11812
rect 1412 11753 1440 11784
rect 9398 11772 9404 11784
rect 9456 11772 9462 11824
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 6638 11744 6644 11756
rect 6595 11716 6644 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6822 11753 6828 11756
rect 6816 11707 6828 11753
rect 6880 11744 6886 11756
rect 6880 11716 6916 11744
rect 6822 11704 6828 11707
rect 6880 11704 6886 11716
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 8389 11747 8447 11753
rect 8389 11744 8401 11747
rect 8260 11716 8401 11744
rect 8260 11704 8266 11716
rect 8389 11713 8401 11716
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 1394 11568 1400 11620
rect 1452 11608 1458 11620
rect 6546 11608 6552 11620
rect 1452 11580 6552 11608
rect 1452 11568 1458 11580
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 7929 11543 7987 11549
rect 7929 11509 7941 11543
rect 7975 11540 7987 11543
rect 8110 11540 8116 11552
rect 7975 11512 8116 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5845 11450
rect 5897 11398 5909 11450
rect 5961 11398 5973 11450
rect 6025 11398 6037 11450
rect 6089 11398 6101 11450
rect 6153 11398 9109 11450
rect 9161 11398 9173 11450
rect 9225 11398 9237 11450
rect 9289 11398 9301 11450
rect 9353 11398 9365 11450
rect 9417 11398 10856 11450
rect 1104 11376 10856 11398
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6822 11336 6828 11348
rect 6503 11308 6828 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7926 11336 7932 11348
rect 6932 11308 7932 11336
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 6932 11268 6960 11308
rect 7926 11296 7932 11308
rect 7984 11336 7990 11348
rect 8205 11339 8263 11345
rect 8205 11336 8217 11339
rect 7984 11308 8217 11336
rect 7984 11296 7990 11308
rect 8205 11305 8217 11308
rect 8251 11305 8263 11339
rect 8205 11299 8263 11305
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 8996 11308 9229 11336
rect 8996 11296 9002 11308
rect 9217 11305 9229 11308
rect 9263 11336 9275 11339
rect 9858 11336 9864 11348
rect 9263 11308 9864 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 9858 11296 9864 11308
rect 9916 11336 9922 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 9916 11308 10241 11336
rect 9916 11296 9922 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 10229 11299 10287 11305
rect 6604 11240 6960 11268
rect 7101 11271 7159 11277
rect 6604 11228 6610 11240
rect 7101 11237 7113 11271
rect 7147 11268 7159 11271
rect 9766 11268 9772 11280
rect 7147 11240 9772 11268
rect 7147 11237 7159 11240
rect 7101 11231 7159 11237
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 9398 11200 9404 11212
rect 1412 11172 9404 11200
rect 1412 11141 1440 11172
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 7282 11132 7288 11144
rect 7243 11104 7288 11132
rect 6641 11095 6699 11101
rect 6656 11064 6684 11095
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 7374 11064 7380 11076
rect 6656 11036 7380 11064
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 1104 10906 10856 10928
rect 1104 10854 4213 10906
rect 4265 10854 4277 10906
rect 4329 10854 4341 10906
rect 4393 10854 4405 10906
rect 4457 10854 4469 10906
rect 4521 10854 7477 10906
rect 7529 10854 7541 10906
rect 7593 10854 7605 10906
rect 7657 10854 7669 10906
rect 7721 10854 7733 10906
rect 7785 10854 10856 10906
rect 1104 10832 10856 10854
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 5684 10764 7113 10792
rect 5684 10752 5690 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 7837 10795 7895 10801
rect 7837 10761 7849 10795
rect 7883 10792 7895 10795
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 7883 10764 9781 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 9769 10761 9781 10764
rect 9815 10761 9827 10795
rect 9769 10755 9827 10761
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 9916 10764 9961 10792
rect 9916 10752 9922 10764
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 9490 10724 9496 10736
rect 8812 10696 9496 10724
rect 8812 10684 8818 10696
rect 9490 10684 9496 10696
rect 9548 10684 9554 10736
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7190 10656 7196 10668
rect 6963 10628 7196 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 1412 10588 1440 10619
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 8018 10656 8024 10668
rect 7979 10628 8024 10656
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8846 10656 8852 10668
rect 8807 10628 8852 10656
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 10410 10656 10416 10668
rect 10371 10628 10416 10656
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 8754 10588 8760 10600
rect 1412 10560 8760 10588
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 8938 10588 8944 10600
rect 8899 10560 8944 10588
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9950 10588 9956 10600
rect 9171 10560 9956 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 8481 10523 8539 10529
rect 8481 10520 8493 10523
rect 7156 10492 8493 10520
rect 7156 10480 7162 10492
rect 8481 10489 8493 10492
rect 8527 10489 8539 10523
rect 9398 10520 9404 10532
rect 9359 10492 9404 10520
rect 8481 10483 8539 10489
rect 9398 10480 9404 10492
rect 9456 10480 9462 10532
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9824 10424 10241 10452
rect 9824 10412 9830 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5845 10362
rect 5897 10310 5909 10362
rect 5961 10310 5973 10362
rect 6025 10310 6037 10362
rect 6089 10310 6101 10362
rect 6153 10310 9109 10362
rect 9161 10310 9173 10362
rect 9225 10310 9237 10362
rect 9289 10310 9301 10362
rect 9353 10310 9365 10362
rect 9417 10310 10856 10362
rect 1104 10288 10856 10310
rect 7190 10248 7196 10260
rect 7151 10220 7196 10248
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 8812 10220 9413 10248
rect 8812 10208 8818 10220
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9401 10211 9459 10217
rect 8205 10183 8263 10189
rect 8205 10149 8217 10183
rect 8251 10180 8263 10183
rect 9674 10180 9680 10192
rect 8251 10152 9680 10180
rect 8251 10149 8263 10152
rect 8205 10143 8263 10149
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 11609 10183 11667 10189
rect 11609 10180 11621 10183
rect 9784 10152 11621 10180
rect 9784 10112 9812 10152
rect 11609 10149 11621 10152
rect 11655 10149 11667 10183
rect 11609 10143 11667 10149
rect 9950 10112 9956 10124
rect 2746 10084 9812 10112
rect 9911 10084 9956 10112
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2746 10044 2774 10084
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 7098 10044 7104 10056
rect 1443 10016 2774 10044
rect 7059 10016 7104 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 8386 10044 8392 10056
rect 8347 10016 8392 10044
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 9766 10044 9772 10056
rect 9727 10016 9772 10044
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 9861 9979 9919 9985
rect 9861 9976 9873 9979
rect 4764 9948 9873 9976
rect 4764 9936 4770 9948
rect 9861 9945 9873 9948
rect 9907 9945 9919 9979
rect 9861 9939 9919 9945
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 1104 9818 10856 9840
rect 1104 9766 4213 9818
rect 4265 9766 4277 9818
rect 4329 9766 4341 9818
rect 4393 9766 4405 9818
rect 4457 9766 4469 9818
rect 4521 9766 7477 9818
rect 7529 9766 7541 9818
rect 7593 9766 7605 9818
rect 7657 9766 7669 9818
rect 7721 9766 7733 9818
rect 7785 9766 10856 9818
rect 1104 9744 10856 9766
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 8665 9639 8723 9645
rect 8665 9636 8677 9639
rect 8536 9608 8677 9636
rect 8536 9596 8542 9608
rect 8665 9605 8677 9608
rect 8711 9605 8723 9639
rect 8846 9636 8852 9648
rect 8807 9608 8852 9636
rect 8665 9599 8723 9605
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 7834 9568 7840 9580
rect 7795 9540 7840 9568
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 9766 9568 9772 9580
rect 9727 9540 9772 9568
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 8021 9435 8079 9441
rect 8021 9432 8033 9435
rect 1912 9404 8033 9432
rect 1912 9392 1918 9404
rect 8021 9401 8033 9404
rect 8067 9401 8079 9435
rect 8021 9395 8079 9401
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 9214 9432 9220 9444
rect 8904 9404 9220 9432
rect 8904 9392 8910 9404
rect 9214 9392 9220 9404
rect 9272 9392 9278 9444
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 5592 9336 9873 9364
rect 5592 9324 5598 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5845 9274
rect 5897 9222 5909 9274
rect 5961 9222 5973 9274
rect 6025 9222 6037 9274
rect 6089 9222 6101 9274
rect 6153 9222 9109 9274
rect 9161 9222 9173 9274
rect 9225 9222 9237 9274
rect 9289 9222 9301 9274
rect 9353 9222 9365 9274
rect 9417 9222 10856 9274
rect 1104 9200 10856 9222
rect 5442 9120 5448 9172
rect 5500 9160 5506 9172
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 5500 9132 9321 9160
rect 5500 9120 5506 9132
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 9309 9123 9367 9129
rect 10045 9163 10103 9169
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 11701 9163 11759 9169
rect 11701 9160 11713 9163
rect 10091 9132 11713 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 11701 9129 11713 9132
rect 11747 9129 11759 9163
rect 11701 9123 11759 9129
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 2746 8996 11529 9024
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 2746 8956 2774 8996
rect 11517 8993 11529 8996
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 9122 8956 9128 8968
rect 1443 8928 2774 8956
rect 9083 8928 9128 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9858 8956 9864 8968
rect 9819 8928 9864 8956
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 1104 8730 10856 8752
rect 1104 8678 4213 8730
rect 4265 8678 4277 8730
rect 4329 8678 4341 8730
rect 4393 8678 4405 8730
rect 4457 8678 4469 8730
rect 4521 8678 7477 8730
rect 7529 8678 7541 8730
rect 7593 8678 7605 8730
rect 7657 8678 7669 8730
rect 7721 8678 7733 8730
rect 7785 8678 10856 8730
rect 1104 8656 10856 8678
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8996 8588 9229 8616
rect 8996 8576 9002 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9217 8579 9275 8585
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 10459 8588 11805 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 9125 8551 9183 8557
rect 9125 8517 9137 8551
rect 9171 8548 9183 8551
rect 9582 8548 9588 8560
rect 9171 8520 9588 8548
rect 9171 8517 9183 8520
rect 9125 8511 9183 8517
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 10965 8551 11023 8557
rect 10965 8548 10977 8551
rect 9815 8520 10977 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10965 8517 10977 8520
rect 11011 8517 11023 8551
rect 10965 8511 11023 8517
rect 750 8440 756 8492
rect 808 8480 814 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 808 8452 1409 8480
rect 808 8440 814 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 10226 8480 10232 8492
rect 10187 8452 10232 8480
rect 1397 8443 1455 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 10091 8384 11437 8412
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 1578 8344 1584 8356
rect 1539 8316 1584 8344
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5845 8186
rect 5897 8134 5909 8186
rect 5961 8134 5973 8186
rect 6025 8134 6037 8186
rect 6089 8134 6101 8186
rect 6153 8134 9109 8186
rect 9161 8134 9173 8186
rect 9225 8134 9237 8186
rect 9289 8134 9301 8186
rect 9353 8134 9365 8186
rect 9417 8134 10856 8186
rect 1104 8112 10856 8134
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 10091 8044 11345 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 11333 8041 11345 8044
rect 11379 8041 11391 8075
rect 11333 8035 11391 8041
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 1670 7868 1676 7880
rect 1443 7840 1676 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 9766 7800 9772 7812
rect 9727 7772 9772 7800
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 1104 7642 10856 7664
rect 1104 7590 4213 7642
rect 4265 7590 4277 7642
rect 4329 7590 4341 7642
rect 4393 7590 4405 7642
rect 4457 7590 4469 7642
rect 4521 7590 7477 7642
rect 7529 7590 7541 7642
rect 7593 7590 7605 7642
rect 7657 7590 7669 7642
rect 7721 7590 7733 7642
rect 7785 7590 10856 7642
rect 1104 7568 10856 7590
rect 5166 7488 5172 7540
rect 5224 7528 5230 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 5224 7500 9137 7528
rect 5224 7488 5230 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 11057 7531 11115 7537
rect 11057 7528 11069 7531
rect 9907 7500 11069 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 11057 7497 11069 7500
rect 11103 7497 11115 7531
rect 11057 7491 11115 7497
rect 1210 7352 1216 7404
rect 1268 7392 1274 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 1268 7364 1409 7392
rect 1268 7352 1274 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 8938 7392 8944 7404
rect 8899 7364 8944 7392
rect 1397 7355 1455 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 9769 7395 9827 7401
rect 9769 7392 9781 7395
rect 9732 7364 9781 7392
rect 9732 7352 9738 7364
rect 9769 7361 9781 7364
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 8386 7216 8392 7268
rect 8444 7256 8450 7268
rect 9401 7259 9459 7265
rect 9401 7256 9413 7259
rect 8444 7228 9413 7256
rect 8444 7216 8450 7228
rect 9401 7225 9413 7228
rect 9447 7225 9459 7259
rect 9401 7219 9459 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 8754 7188 8760 7200
rect 8628 7160 8760 7188
rect 8628 7148 8634 7160
rect 8754 7148 8760 7160
rect 8812 7148 8818 7200
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5845 7098
rect 5897 7046 5909 7098
rect 5961 7046 5973 7098
rect 6025 7046 6037 7098
rect 6089 7046 6101 7098
rect 6153 7046 9109 7098
rect 9161 7046 9173 7098
rect 9225 7046 9237 7098
rect 9289 7046 9301 7098
rect 9353 7046 9365 7098
rect 9417 7046 10856 7098
rect 1104 7024 10856 7046
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 8904 6820 9873 6848
rect 8904 6808 8910 6820
rect 9861 6817 9873 6820
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10008 6820 10053 6848
rect 10008 6808 10014 6820
rect 10962 6780 10968 6792
rect 10923 6752 10968 6780
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 9030 6672 9036 6724
rect 9088 6712 9094 6724
rect 9769 6715 9827 6721
rect 9769 6712 9781 6715
rect 9088 6684 9781 6712
rect 9088 6672 9094 6684
rect 9769 6681 9781 6684
rect 9815 6681 9827 6715
rect 9769 6675 9827 6681
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 8720 6616 9413 6644
rect 8720 6604 8726 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 1104 6554 10856 6576
rect 1104 6502 4213 6554
rect 4265 6502 4277 6554
rect 4329 6502 4341 6554
rect 4393 6502 4405 6554
rect 4457 6502 4469 6554
rect 4521 6502 7477 6554
rect 7529 6502 7541 6554
rect 7593 6502 7605 6554
rect 7657 6502 7669 6554
rect 7721 6502 7733 6554
rect 7785 6502 10856 6554
rect 1104 6480 10856 6502
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 8904 6412 9229 6440
rect 8904 6400 8910 6412
rect 9217 6409 9229 6412
rect 9263 6440 9275 6443
rect 10229 6443 10287 6449
rect 10229 6440 10241 6443
rect 9263 6412 10241 6440
rect 9263 6409 9275 6412
rect 9217 6403 9275 6409
rect 10229 6409 10241 6412
rect 10275 6409 10287 6443
rect 10229 6403 10287 6409
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1486 6304 1492 6316
rect 1443 6276 1492 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1486 6264 1492 6276
rect 1544 6264 1550 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 6236 6276 8769 6304
rect 6236 6264 6242 6276
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 1578 6168 1584 6180
rect 1539 6140 1584 6168
rect 1578 6128 1584 6140
rect 1636 6128 1642 6180
rect 8846 6100 8852 6112
rect 8807 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5845 6010
rect 5897 5958 5909 6010
rect 5961 5958 5973 6010
rect 6025 5958 6037 6010
rect 6089 5958 6101 6010
rect 6153 5958 9109 6010
rect 9161 5958 9173 6010
rect 9225 5958 9237 6010
rect 9289 5958 9301 6010
rect 9353 5958 9365 6010
rect 9417 5958 10856 6010
rect 1104 5936 10856 5958
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 8904 5732 9413 5760
rect 8904 5720 8910 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9585 5763 9643 5769
rect 9585 5729 9597 5763
rect 9631 5760 9643 5763
rect 9950 5760 9956 5772
rect 9631 5732 9956 5760
rect 9631 5729 9643 5732
rect 9585 5723 9643 5729
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 5718 5692 5724 5704
rect 1443 5664 5724 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 8018 5692 8024 5704
rect 6788 5664 8024 5692
rect 6788 5652 6794 5664
rect 8018 5652 8024 5664
rect 8076 5692 8082 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 8076 5664 8125 5692
rect 8076 5652 8082 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8435 5596 9321 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9309 5587 9367 5593
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 8628 5528 8953 5556
rect 8628 5516 8634 5528
rect 8941 5525 8953 5528
rect 8987 5525 8999 5559
rect 8941 5519 8999 5525
rect 1104 5466 10856 5488
rect 1104 5414 4213 5466
rect 4265 5414 4277 5466
rect 4329 5414 4341 5466
rect 4393 5414 4405 5466
rect 4457 5414 4469 5466
rect 4521 5414 7477 5466
rect 7529 5414 7541 5466
rect 7593 5414 7605 5466
rect 7657 5414 7669 5466
rect 7721 5414 7733 5466
rect 7785 5414 10856 5466
rect 1104 5392 10856 5414
rect 8113 5355 8171 5361
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 9674 5352 9680 5364
rect 8159 5324 9680 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 11149 5355 11207 5361
rect 11149 5352 11161 5355
rect 9907 5324 11161 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 11149 5321 11161 5324
rect 11195 5321 11207 5355
rect 11149 5315 11207 5321
rect 9309 5287 9367 5293
rect 9309 5253 9321 5287
rect 9355 5284 9367 5287
rect 9876 5284 9904 5315
rect 9355 5256 9904 5284
rect 9355 5253 9367 5256
rect 9309 5247 9367 5253
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1762 5216 1768 5228
rect 1443 5188 1768 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8168 5188 8309 5216
rect 8168 5176 8174 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8938 5216 8944 5228
rect 8899 5188 8944 5216
rect 8297 5179 8355 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 8754 5108 8760 5160
rect 8812 5148 8818 5160
rect 9582 5148 9588 5160
rect 8812 5120 9588 5148
rect 8812 5108 8818 5120
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9950 5148 9956 5160
rect 9911 5120 9956 5148
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 9401 5083 9459 5089
rect 9401 5080 9413 5083
rect 5592 5052 9413 5080
rect 5592 5040 5598 5052
rect 9401 5049 9413 5052
rect 9447 5049 9459 5083
rect 9401 5043 9459 5049
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 8754 5012 8760 5024
rect 8715 4984 8760 5012
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5845 4922
rect 5897 4870 5909 4922
rect 5961 4870 5973 4922
rect 6025 4870 6037 4922
rect 6089 4870 6101 4922
rect 6153 4870 9109 4922
rect 9161 4870 9173 4922
rect 9225 4870 9237 4922
rect 9289 4870 9301 4922
rect 9353 4870 9365 4922
rect 9417 4870 10856 4922
rect 1104 4848 10856 4870
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 9582 4808 9588 4820
rect 9355 4780 9588 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 9600 4672 9628 4768
rect 9861 4675 9919 4681
rect 9861 4672 9873 4675
rect 9600 4644 9873 4672
rect 9861 4641 9873 4644
rect 9907 4641 9919 4675
rect 9861 4635 9919 4641
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10008 4644 10053 4672
rect 10008 4632 10014 4644
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 8386 4604 8392 4616
rect 1443 4576 8392 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 8812 4576 9781 4604
rect 8812 4564 8818 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 9398 4468 9404 4480
rect 9359 4440 9404 4468
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 1104 4378 10856 4400
rect 1104 4326 4213 4378
rect 4265 4326 4277 4378
rect 4329 4326 4341 4378
rect 4393 4326 4405 4378
rect 4457 4326 4469 4378
rect 4521 4326 7477 4378
rect 7529 4326 7541 4378
rect 7593 4326 7605 4378
rect 7657 4326 7669 4378
rect 7721 4326 7733 4378
rect 7785 4326 10856 4378
rect 1104 4304 10856 4326
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 8076 4236 9536 4264
rect 8076 4224 8082 4236
rect 9398 4196 9404 4208
rect 8312 4168 9404 4196
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 8312 4128 8340 4168
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 9508 4196 9536 4236
rect 9508 4168 9628 4196
rect 1443 4100 8340 4128
rect 8849 4131 8907 4137
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9122 4128 9128 4140
rect 8895 4100 9128 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 9490 4128 9496 4140
rect 9355 4100 9496 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 9600 4137 9628 4168
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4097 9643 4131
rect 9585 4091 9643 4097
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 9214 4060 9220 4072
rect 8996 4032 9220 4060
rect 8996 4020 9002 4032
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 8665 3995 8723 4001
rect 8665 3961 8677 3995
rect 8711 3992 8723 3995
rect 9030 3992 9036 4004
rect 8711 3964 9036 3992
rect 8711 3961 8723 3964
rect 8665 3955 8723 3961
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5845 3834
rect 5897 3782 5909 3834
rect 5961 3782 5973 3834
rect 6025 3782 6037 3834
rect 6089 3782 6101 3834
rect 6153 3782 9109 3834
rect 9161 3782 9173 3834
rect 9225 3782 9237 3834
rect 9289 3782 9301 3834
rect 9353 3782 9365 3834
rect 9417 3782 10856 3834
rect 1104 3760 10856 3782
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 9766 3720 9772 3732
rect 8251 3692 9772 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 8662 3584 8668 3596
rect 2746 3556 8668 3584
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3516 1455 3519
rect 2746 3516 2774 3556
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 8904 3556 9597 3584
rect 8904 3544 8910 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 1443 3488 2774 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8168 3488 8401 3516
rect 8168 3476 8174 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9490 3516 9496 3528
rect 9355 3488 9496 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 1104 3290 10856 3312
rect 1104 3238 4213 3290
rect 4265 3238 4277 3290
rect 4329 3238 4341 3290
rect 4393 3238 4405 3290
rect 4457 3238 4469 3290
rect 4521 3238 7477 3290
rect 7529 3238 7541 3290
rect 7593 3238 7605 3290
rect 7657 3238 7669 3290
rect 7721 3238 7733 3290
rect 7785 3238 10856 3290
rect 1104 3216 10856 3238
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 9950 3176 9956 3188
rect 9907 3148 9956 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 8570 3108 8576 3120
rect 2746 3080 8576 3108
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 2746 3040 2774 3080
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 1443 3012 2774 3040
rect 7653 3043 7711 3049
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 7653 3009 7665 3043
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 7668 2972 7696 3003
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 8389 3043 8447 3049
rect 8389 3040 8401 3043
rect 8168 3012 8401 3040
rect 8168 3000 8174 3012
rect 8389 3009 8401 3012
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8938 2972 8944 2984
rect 7668 2944 8944 2972
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 7834 2904 7840 2916
rect 7795 2876 7840 2904
rect 7834 2864 7840 2876
rect 7892 2864 7898 2916
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8570 2904 8576 2916
rect 8352 2876 8576 2904
rect 8352 2864 8358 2876
rect 8570 2864 8576 2876
rect 8628 2864 8634 2916
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1452 2808 1593 2836
rect 1452 2796 1458 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5845 2746
rect 5897 2694 5909 2746
rect 5961 2694 5973 2746
rect 6025 2694 6037 2746
rect 6089 2694 6101 2746
rect 6153 2694 9109 2746
rect 9161 2694 9173 2746
rect 9225 2694 9237 2746
rect 9289 2694 9301 2746
rect 9353 2694 9365 2746
rect 9417 2694 10856 2746
rect 1104 2672 10856 2694
rect 5534 2496 5540 2508
rect 2148 2468 5540 2496
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2428 1455 2431
rect 1486 2428 1492 2440
rect 1443 2400 1492 2428
rect 1443 2397 1455 2400
rect 1397 2391 1455 2397
rect 1486 2388 1492 2400
rect 1544 2388 1550 2440
rect 2148 2437 2176 2468
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 7561 2499 7619 2505
rect 7561 2465 7573 2499
rect 7607 2496 7619 2499
rect 7926 2496 7932 2508
rect 7607 2468 7932 2496
rect 7607 2465 7619 2468
rect 7561 2459 7619 2465
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 8536 2468 9597 2496
rect 8536 2456 8542 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 7098 2428 7104 2440
rect 3099 2400 7104 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8570 2428 8576 2440
rect 7883 2400 8576 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 2314 2292 2320 2304
rect 2275 2264 2320 2292
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 1104 2202 10856 2224
rect 1104 2150 4213 2202
rect 4265 2150 4277 2202
rect 4329 2150 4341 2202
rect 4393 2150 4405 2202
rect 4457 2150 4469 2202
rect 4521 2150 7477 2202
rect 7529 2150 7541 2202
rect 7593 2150 7605 2202
rect 7657 2150 7669 2202
rect 7721 2150 7733 2202
rect 7785 2150 10856 2202
rect 1104 2128 10856 2150
<< via1 >>
rect 2582 77766 2634 77818
rect 2646 77766 2698 77818
rect 2710 77766 2762 77818
rect 2774 77766 2826 77818
rect 2838 77766 2890 77818
rect 5845 77766 5897 77818
rect 5909 77766 5961 77818
rect 5973 77766 6025 77818
rect 6037 77766 6089 77818
rect 6101 77766 6153 77818
rect 9109 77766 9161 77818
rect 9173 77766 9225 77818
rect 9237 77766 9289 77818
rect 9301 77766 9353 77818
rect 9365 77766 9417 77818
rect 7564 77707 7616 77716
rect 7564 77673 7573 77707
rect 7573 77673 7607 77707
rect 7607 77673 7616 77707
rect 7564 77664 7616 77673
rect 8208 77664 8260 77716
rect 1400 77571 1452 77580
rect 1400 77537 1409 77571
rect 1409 77537 1443 77571
rect 1443 77537 1452 77571
rect 1400 77528 1452 77537
rect 2872 77503 2924 77512
rect 2872 77469 2881 77503
rect 2881 77469 2915 77503
rect 2915 77469 2924 77503
rect 2872 77460 2924 77469
rect 6184 77460 6236 77512
rect 3148 77392 3200 77444
rect 8944 77460 8996 77512
rect 3056 77324 3108 77376
rect 9312 77367 9364 77376
rect 9312 77333 9321 77367
rect 9321 77333 9355 77367
rect 9355 77333 9364 77367
rect 9312 77324 9364 77333
rect 10140 77324 10192 77376
rect 4213 77222 4265 77274
rect 4277 77222 4329 77274
rect 4341 77222 4393 77274
rect 4405 77222 4457 77274
rect 4469 77222 4521 77274
rect 7477 77222 7529 77274
rect 7541 77222 7593 77274
rect 7605 77222 7657 77274
rect 7669 77222 7721 77274
rect 7733 77222 7785 77274
rect 3700 77120 3752 77172
rect 8576 77163 8628 77172
rect 8576 77129 8585 77163
rect 8585 77129 8619 77163
rect 8619 77129 8628 77163
rect 8576 77120 8628 77129
rect 9588 77120 9640 77172
rect 1584 77027 1636 77036
rect 1584 76993 1593 77027
rect 1593 76993 1627 77027
rect 1627 76993 1636 77027
rect 1584 76984 1636 76993
rect 2964 77052 3016 77104
rect 3240 76984 3292 77036
rect 8392 77027 8444 77036
rect 8392 76993 8401 77027
rect 8401 76993 8435 77027
rect 8435 76993 8444 77027
rect 8392 76984 8444 76993
rect 3332 76916 3384 76968
rect 2964 76848 3016 76900
rect 6460 76780 6512 76832
rect 10048 76823 10100 76832
rect 10048 76789 10057 76823
rect 10057 76789 10091 76823
rect 10091 76789 10100 76823
rect 10048 76780 10100 76789
rect 2582 76678 2634 76730
rect 2646 76678 2698 76730
rect 2710 76678 2762 76730
rect 2774 76678 2826 76730
rect 2838 76678 2890 76730
rect 5845 76678 5897 76730
rect 5909 76678 5961 76730
rect 5973 76678 6025 76730
rect 6037 76678 6089 76730
rect 6101 76678 6153 76730
rect 9109 76678 9161 76730
rect 9173 76678 9225 76730
rect 9237 76678 9289 76730
rect 9301 76678 9353 76730
rect 9365 76678 9417 76730
rect 9496 76576 9548 76628
rect 1584 76415 1636 76424
rect 1584 76381 1593 76415
rect 1593 76381 1627 76415
rect 1627 76381 1636 76415
rect 1584 76372 1636 76381
rect 8300 76372 8352 76424
rect 2136 76236 2188 76288
rect 10048 76279 10100 76288
rect 10048 76245 10057 76279
rect 10057 76245 10091 76279
rect 10091 76245 10100 76279
rect 10048 76236 10100 76245
rect 4213 76134 4265 76186
rect 4277 76134 4329 76186
rect 4341 76134 4393 76186
rect 4405 76134 4457 76186
rect 4469 76134 4521 76186
rect 7477 76134 7529 76186
rect 7541 76134 7593 76186
rect 7605 76134 7657 76186
rect 7669 76134 7721 76186
rect 7733 76134 7785 76186
rect 9312 76075 9364 76084
rect 9312 76041 9321 76075
rect 9321 76041 9355 76075
rect 9355 76041 9364 76075
rect 9312 76032 9364 76041
rect 1768 75896 1820 75948
rect 8484 75896 8536 75948
rect 9864 75939 9916 75948
rect 9864 75905 9873 75939
rect 9873 75905 9907 75939
rect 9907 75905 9916 75939
rect 9864 75896 9916 75905
rect 1400 75871 1452 75880
rect 1400 75837 1409 75871
rect 1409 75837 1443 75871
rect 1443 75837 1452 75871
rect 1400 75828 1452 75837
rect 2582 75590 2634 75642
rect 2646 75590 2698 75642
rect 2710 75590 2762 75642
rect 2774 75590 2826 75642
rect 2838 75590 2890 75642
rect 5845 75590 5897 75642
rect 5909 75590 5961 75642
rect 5973 75590 6025 75642
rect 6037 75590 6089 75642
rect 6101 75590 6153 75642
rect 9109 75590 9161 75642
rect 9173 75590 9225 75642
rect 9237 75590 9289 75642
rect 9301 75590 9353 75642
rect 9365 75590 9417 75642
rect 1860 75259 1912 75268
rect 1860 75225 1869 75259
rect 1869 75225 1903 75259
rect 1903 75225 1912 75259
rect 1860 75216 1912 75225
rect 1952 75191 2004 75200
rect 1952 75157 1961 75191
rect 1961 75157 1995 75191
rect 1995 75157 2004 75191
rect 1952 75148 2004 75157
rect 10140 75148 10192 75200
rect 4213 75046 4265 75098
rect 4277 75046 4329 75098
rect 4341 75046 4393 75098
rect 4405 75046 4457 75098
rect 4469 75046 4521 75098
rect 7477 75046 7529 75098
rect 7541 75046 7593 75098
rect 7605 75046 7657 75098
rect 7669 75046 7721 75098
rect 7733 75046 7785 75098
rect 3056 74987 3108 74996
rect 3056 74953 3065 74987
rect 3065 74953 3099 74987
rect 3099 74953 3108 74987
rect 3056 74944 3108 74953
rect 3148 74876 3200 74928
rect 10968 74919 11020 74928
rect 10968 74885 10977 74919
rect 10977 74885 11011 74919
rect 11011 74885 11020 74919
rect 10968 74876 11020 74885
rect 1584 74851 1636 74860
rect 1584 74817 1593 74851
rect 1593 74817 1627 74851
rect 1627 74817 1636 74851
rect 1584 74808 1636 74817
rect 2228 74851 2280 74860
rect 2228 74817 2237 74851
rect 2237 74817 2271 74851
rect 2271 74817 2280 74851
rect 2228 74808 2280 74817
rect 2504 74740 2556 74792
rect 3148 74783 3200 74792
rect 3148 74749 3157 74783
rect 3157 74749 3191 74783
rect 3191 74749 3200 74783
rect 3148 74740 3200 74749
rect 2044 74647 2096 74656
rect 2044 74613 2053 74647
rect 2053 74613 2087 74647
rect 2087 74613 2096 74647
rect 2044 74604 2096 74613
rect 4620 74604 4672 74656
rect 10048 74647 10100 74656
rect 10048 74613 10057 74647
rect 10057 74613 10091 74647
rect 10091 74613 10100 74647
rect 10048 74604 10100 74613
rect 2582 74502 2634 74554
rect 2646 74502 2698 74554
rect 2710 74502 2762 74554
rect 2774 74502 2826 74554
rect 2838 74502 2890 74554
rect 5845 74502 5897 74554
rect 5909 74502 5961 74554
rect 5973 74502 6025 74554
rect 6037 74502 6089 74554
rect 6101 74502 6153 74554
rect 9109 74502 9161 74554
rect 9173 74502 9225 74554
rect 9237 74502 9289 74554
rect 9301 74502 9353 74554
rect 9365 74502 9417 74554
rect 6184 74400 6236 74452
rect 8392 74400 8444 74452
rect 8944 74332 8996 74384
rect 2504 74307 2556 74316
rect 2504 74273 2513 74307
rect 2513 74273 2547 74307
rect 2547 74273 2556 74307
rect 2504 74264 2556 74273
rect 6828 74264 6880 74316
rect 10232 74264 10284 74316
rect 2320 74196 2372 74248
rect 6460 74171 6512 74180
rect 6460 74137 6469 74171
rect 6469 74137 6503 74171
rect 6503 74137 6512 74171
rect 6460 74128 6512 74137
rect 6644 74128 6696 74180
rect 9956 74128 10008 74180
rect 2136 74060 2188 74112
rect 6368 74060 6420 74112
rect 10140 74060 10192 74112
rect 4213 73958 4265 74010
rect 4277 73958 4329 74010
rect 4341 73958 4393 74010
rect 4405 73958 4457 74010
rect 4469 73958 4521 74010
rect 7477 73958 7529 74010
rect 7541 73958 7593 74010
rect 7605 73958 7657 74010
rect 7669 73958 7721 74010
rect 7733 73958 7785 74010
rect 3332 73899 3384 73908
rect 3332 73865 3341 73899
rect 3341 73865 3375 73899
rect 3375 73865 3384 73899
rect 3332 73856 3384 73865
rect 1952 73763 2004 73772
rect 1952 73729 1961 73763
rect 1961 73729 1995 73763
rect 1995 73729 2004 73763
rect 1952 73720 2004 73729
rect 2412 73720 2464 73772
rect 3700 73763 3752 73772
rect 3700 73729 3709 73763
rect 3709 73729 3743 73763
rect 3743 73729 3752 73763
rect 3700 73720 3752 73729
rect 4068 73720 4120 73772
rect 8668 73720 8720 73772
rect 2504 73652 2556 73704
rect 6828 73652 6880 73704
rect 1952 73584 2004 73636
rect 9496 73516 9548 73568
rect 10048 73559 10100 73568
rect 10048 73525 10057 73559
rect 10057 73525 10091 73559
rect 10091 73525 10100 73559
rect 10048 73516 10100 73525
rect 2582 73414 2634 73466
rect 2646 73414 2698 73466
rect 2710 73414 2762 73466
rect 2774 73414 2826 73466
rect 2838 73414 2890 73466
rect 5845 73414 5897 73466
rect 5909 73414 5961 73466
rect 5973 73414 6025 73466
rect 6037 73414 6089 73466
rect 6101 73414 6153 73466
rect 9109 73414 9161 73466
rect 9173 73414 9225 73466
rect 9237 73414 9289 73466
rect 9301 73414 9353 73466
rect 9365 73414 9417 73466
rect 2136 73312 2188 73364
rect 2596 73244 2648 73296
rect 2504 73176 2556 73228
rect 6828 73176 6880 73228
rect 10140 73176 10192 73228
rect 1676 73108 1728 73160
rect 2872 73151 2924 73160
rect 2872 73117 2881 73151
rect 2881 73117 2915 73151
rect 2915 73117 2924 73151
rect 2872 73108 2924 73117
rect 6920 73040 6972 73092
rect 1768 72972 1820 73024
rect 2136 72972 2188 73024
rect 7012 72972 7064 73024
rect 9864 73108 9916 73160
rect 10232 73108 10284 73160
rect 7380 73040 7432 73092
rect 9956 73083 10008 73092
rect 9956 73049 9965 73083
rect 9965 73049 9999 73083
rect 9999 73049 10008 73083
rect 9956 73040 10008 73049
rect 7288 72972 7340 73024
rect 8576 72972 8628 73024
rect 4213 72870 4265 72922
rect 4277 72870 4329 72922
rect 4341 72870 4393 72922
rect 4405 72870 4457 72922
rect 4469 72870 4521 72922
rect 7477 72870 7529 72922
rect 7541 72870 7593 72922
rect 7605 72870 7657 72922
rect 7669 72870 7721 72922
rect 7733 72870 7785 72922
rect 1768 72811 1820 72820
rect 1768 72777 1777 72811
rect 1777 72777 1811 72811
rect 1811 72777 1820 72811
rect 1768 72768 1820 72777
rect 2044 72768 2096 72820
rect 8300 72768 8352 72820
rect 2228 72700 2280 72752
rect 2504 72700 2556 72752
rect 940 72632 992 72684
rect 2964 72675 3016 72684
rect 1860 72607 1912 72616
rect 1860 72573 1869 72607
rect 1869 72573 1903 72607
rect 1903 72573 1912 72607
rect 1860 72564 1912 72573
rect 2228 72564 2280 72616
rect 2964 72641 2973 72675
rect 2973 72641 3007 72675
rect 3007 72641 3016 72675
rect 2964 72632 3016 72641
rect 6920 72700 6972 72752
rect 9036 72632 9088 72684
rect 9312 72539 9364 72548
rect 9312 72505 9321 72539
rect 9321 72505 9355 72539
rect 9355 72505 9364 72539
rect 9312 72496 9364 72505
rect 8484 72428 8536 72480
rect 10140 72428 10192 72480
rect 2582 72326 2634 72378
rect 2646 72326 2698 72378
rect 2710 72326 2762 72378
rect 2774 72326 2826 72378
rect 2838 72326 2890 72378
rect 5845 72326 5897 72378
rect 5909 72326 5961 72378
rect 5973 72326 6025 72378
rect 6037 72326 6089 72378
rect 6101 72326 6153 72378
rect 9109 72326 9161 72378
rect 9173 72326 9225 72378
rect 9237 72326 9289 72378
rect 9301 72326 9353 72378
rect 9365 72326 9417 72378
rect 3148 72156 3200 72208
rect 6184 72199 6236 72208
rect 6184 72165 6193 72199
rect 6193 72165 6227 72199
rect 6227 72165 6236 72199
rect 6184 72156 6236 72165
rect 3700 72088 3752 72140
rect 1584 72063 1636 72072
rect 1584 72029 1593 72063
rect 1593 72029 1627 72063
rect 1627 72029 1636 72063
rect 1584 72020 1636 72029
rect 2228 72063 2280 72072
rect 2228 72029 2237 72063
rect 2237 72029 2271 72063
rect 2271 72029 2280 72063
rect 2228 72020 2280 72029
rect 4068 72063 4120 72072
rect 4068 72029 4077 72063
rect 4077 72029 4111 72063
rect 4111 72029 4120 72063
rect 4068 72020 4120 72029
rect 4804 71995 4856 72004
rect 4804 71961 4813 71995
rect 4813 71961 4847 71995
rect 4847 71961 4856 71995
rect 4804 71952 4856 71961
rect 5724 71952 5776 72004
rect 6368 71952 6420 72004
rect 6644 71995 6696 72004
rect 6644 71961 6653 71995
rect 6653 71961 6687 71995
rect 6687 71961 6696 71995
rect 6644 71952 6696 71961
rect 6828 72020 6880 72072
rect 6920 71952 6972 72004
rect 2044 71927 2096 71936
rect 2044 71893 2053 71927
rect 2053 71893 2087 71927
rect 2087 71893 2096 71927
rect 2044 71884 2096 71893
rect 9312 71927 9364 71936
rect 9312 71893 9321 71927
rect 9321 71893 9355 71927
rect 9355 71893 9364 71927
rect 9312 71884 9364 71893
rect 10048 71927 10100 71936
rect 10048 71893 10057 71927
rect 10057 71893 10091 71927
rect 10091 71893 10100 71927
rect 10048 71884 10100 71893
rect 4213 71782 4265 71834
rect 4277 71782 4329 71834
rect 4341 71782 4393 71834
rect 4405 71782 4457 71834
rect 4469 71782 4521 71834
rect 7477 71782 7529 71834
rect 7541 71782 7593 71834
rect 7605 71782 7657 71834
rect 7669 71782 7721 71834
rect 7733 71782 7785 71834
rect 1492 71544 1544 71596
rect 2136 71476 2188 71528
rect 2320 71476 2372 71528
rect 9772 71340 9824 71392
rect 10140 71340 10192 71392
rect 2582 71238 2634 71290
rect 2646 71238 2698 71290
rect 2710 71238 2762 71290
rect 2774 71238 2826 71290
rect 2838 71238 2890 71290
rect 5845 71238 5897 71290
rect 5909 71238 5961 71290
rect 5973 71238 6025 71290
rect 6037 71238 6089 71290
rect 6101 71238 6153 71290
rect 9109 71238 9161 71290
rect 9173 71238 9225 71290
rect 9237 71238 9289 71290
rect 9301 71238 9353 71290
rect 9365 71238 9417 71290
rect 7104 71068 7156 71120
rect 2136 71000 2188 71052
rect 2596 71000 2648 71052
rect 6920 71000 6972 71052
rect 7932 71000 7984 71052
rect 1400 70975 1452 70984
rect 1400 70941 1409 70975
rect 1409 70941 1443 70975
rect 1443 70941 1452 70975
rect 1400 70932 1452 70941
rect 4620 70932 4672 70984
rect 3884 70796 3936 70848
rect 10048 70839 10100 70848
rect 10048 70805 10057 70839
rect 10057 70805 10091 70839
rect 10091 70805 10100 70839
rect 10048 70796 10100 70805
rect 4213 70694 4265 70746
rect 4277 70694 4329 70746
rect 4341 70694 4393 70746
rect 4405 70694 4457 70746
rect 4469 70694 4521 70746
rect 7477 70694 7529 70746
rect 7541 70694 7593 70746
rect 7605 70694 7657 70746
rect 7669 70694 7721 70746
rect 7733 70694 7785 70746
rect 2504 70592 2556 70644
rect 2228 70499 2280 70508
rect 2228 70465 2237 70499
rect 2237 70465 2271 70499
rect 2271 70465 2280 70499
rect 2228 70456 2280 70465
rect 2596 70456 2648 70508
rect 5080 70456 5132 70508
rect 7288 70456 7340 70508
rect 7932 70456 7984 70508
rect 4896 70388 4948 70440
rect 7380 70431 7432 70440
rect 7380 70397 7389 70431
rect 7389 70397 7423 70431
rect 7423 70397 7432 70431
rect 7380 70388 7432 70397
rect 7840 70388 7892 70440
rect 9864 70388 9916 70440
rect 2582 70150 2634 70202
rect 2646 70150 2698 70202
rect 2710 70150 2762 70202
rect 2774 70150 2826 70202
rect 2838 70150 2890 70202
rect 5845 70150 5897 70202
rect 5909 70150 5961 70202
rect 5973 70150 6025 70202
rect 6037 70150 6089 70202
rect 6101 70150 6153 70202
rect 9109 70150 9161 70202
rect 9173 70150 9225 70202
rect 9237 70150 9289 70202
rect 9301 70150 9353 70202
rect 9365 70150 9417 70202
rect 9036 70048 9088 70100
rect 7196 69980 7248 70032
rect 1124 69844 1176 69896
rect 1860 69912 1912 69964
rect 10232 69912 10284 69964
rect 1768 69887 1820 69896
rect 1768 69853 1777 69887
rect 1777 69853 1811 69887
rect 1811 69853 1820 69887
rect 1768 69844 1820 69853
rect 2136 69844 2188 69896
rect 2872 69844 2924 69896
rect 3976 69887 4028 69896
rect 3976 69853 3985 69887
rect 3985 69853 4019 69887
rect 4019 69853 4028 69887
rect 3976 69844 4028 69853
rect 3516 69776 3568 69828
rect 9956 69776 10008 69828
rect 8852 69708 8904 69760
rect 9864 69751 9916 69760
rect 9864 69717 9873 69751
rect 9873 69717 9907 69751
rect 9907 69717 9916 69751
rect 9864 69708 9916 69717
rect 4213 69606 4265 69658
rect 4277 69606 4329 69658
rect 4341 69606 4393 69658
rect 4405 69606 4457 69658
rect 4469 69606 4521 69658
rect 7477 69606 7529 69658
rect 7541 69606 7593 69658
rect 7605 69606 7657 69658
rect 7669 69606 7721 69658
rect 7733 69606 7785 69658
rect 2044 69504 2096 69556
rect 1216 69368 1268 69420
rect 3332 69436 3384 69488
rect 9588 69504 9640 69556
rect 10416 69547 10468 69556
rect 10416 69513 10425 69547
rect 10425 69513 10459 69547
rect 10459 69513 10468 69547
rect 10416 69504 10468 69513
rect 3056 69411 3108 69420
rect 2136 69343 2188 69352
rect 2136 69309 2145 69343
rect 2145 69309 2179 69343
rect 2179 69309 2188 69343
rect 2136 69300 2188 69309
rect 3056 69377 3065 69411
rect 3065 69377 3099 69411
rect 3099 69377 3108 69411
rect 3056 69368 3108 69377
rect 8392 69411 8444 69420
rect 2504 69232 2556 69284
rect 8392 69377 8401 69411
rect 8401 69377 8435 69411
rect 8435 69377 8444 69411
rect 8392 69368 8444 69377
rect 9036 69411 9088 69420
rect 9036 69377 9045 69411
rect 9045 69377 9079 69411
rect 9079 69377 9088 69411
rect 9036 69368 9088 69377
rect 9772 69411 9824 69420
rect 9772 69377 9781 69411
rect 9781 69377 9815 69411
rect 9815 69377 9824 69411
rect 9772 69368 9824 69377
rect 3792 69300 3844 69352
rect 8852 69300 8904 69352
rect 10140 69300 10192 69352
rect 9496 69232 9548 69284
rect 3424 69164 3476 69216
rect 2582 69062 2634 69114
rect 2646 69062 2698 69114
rect 2710 69062 2762 69114
rect 2774 69062 2826 69114
rect 2838 69062 2890 69114
rect 5845 69062 5897 69114
rect 5909 69062 5961 69114
rect 5973 69062 6025 69114
rect 6037 69062 6089 69114
rect 6101 69062 6153 69114
rect 9109 69062 9161 69114
rect 9173 69062 9225 69114
rect 9237 69062 9289 69114
rect 9301 69062 9353 69114
rect 9365 69062 9417 69114
rect 6828 69003 6880 69012
rect 6828 68969 6837 69003
rect 6837 68969 6871 69003
rect 6871 68969 6880 69003
rect 6828 68960 6880 68969
rect 940 68824 992 68876
rect 1584 68799 1636 68808
rect 1584 68765 1593 68799
rect 1593 68765 1627 68799
rect 1627 68765 1636 68799
rect 1584 68756 1636 68765
rect 2964 68824 3016 68876
rect 7932 68824 7984 68876
rect 7196 68799 7248 68808
rect 2504 68688 2556 68740
rect 7196 68765 7205 68799
rect 7205 68765 7239 68799
rect 7239 68765 7248 68799
rect 7196 68756 7248 68765
rect 3240 68731 3292 68740
rect 3240 68697 3249 68731
rect 3249 68697 3283 68731
rect 3283 68697 3292 68731
rect 3240 68688 3292 68697
rect 7012 68688 7064 68740
rect 7932 68688 7984 68740
rect 2320 68620 2372 68672
rect 8208 68620 8260 68672
rect 8576 68620 8628 68672
rect 9496 68620 9548 68672
rect 9864 68620 9916 68672
rect 4213 68518 4265 68570
rect 4277 68518 4329 68570
rect 4341 68518 4393 68570
rect 4405 68518 4457 68570
rect 4469 68518 4521 68570
rect 7477 68518 7529 68570
rect 7541 68518 7593 68570
rect 7605 68518 7657 68570
rect 7669 68518 7721 68570
rect 7733 68518 7785 68570
rect 1492 68280 1544 68332
rect 3884 68416 3936 68468
rect 9956 68459 10008 68468
rect 9956 68425 9965 68459
rect 9965 68425 9999 68459
rect 9999 68425 10008 68459
rect 9956 68416 10008 68425
rect 4620 68348 4672 68400
rect 9496 68348 9548 68400
rect 10140 68348 10192 68400
rect 1308 68212 1360 68264
rect 1584 68144 1636 68196
rect 1952 68144 2004 68196
rect 2504 68144 2556 68196
rect 8208 68280 8260 68332
rect 4620 68212 4672 68264
rect 1768 68076 1820 68128
rect 8760 68119 8812 68128
rect 8760 68085 8769 68119
rect 8769 68085 8803 68119
rect 8803 68085 8812 68119
rect 8760 68076 8812 68085
rect 8852 68076 8904 68128
rect 2582 67974 2634 68026
rect 2646 67974 2698 68026
rect 2710 67974 2762 68026
rect 2774 67974 2826 68026
rect 2838 67974 2890 68026
rect 5845 67974 5897 68026
rect 5909 67974 5961 68026
rect 5973 67974 6025 68026
rect 6037 67974 6089 68026
rect 6101 67974 6153 68026
rect 9109 67974 9161 68026
rect 9173 67974 9225 68026
rect 9237 67974 9289 68026
rect 9301 67974 9353 68026
rect 9365 67974 9417 68026
rect 9404 67847 9456 67856
rect 9404 67813 9413 67847
rect 9413 67813 9447 67847
rect 9447 67813 9456 67847
rect 9404 67804 9456 67813
rect 10140 67736 10192 67788
rect 1400 67711 1452 67720
rect 1400 67677 1409 67711
rect 1409 67677 1443 67711
rect 1443 67677 1452 67711
rect 1400 67668 1452 67677
rect 1952 67668 2004 67720
rect 6920 67668 6972 67720
rect 8852 67600 8904 67652
rect 9772 67600 9824 67652
rect 8300 67575 8352 67584
rect 8300 67541 8309 67575
rect 8309 67541 8343 67575
rect 8343 67541 8352 67575
rect 8300 67532 8352 67541
rect 4213 67430 4265 67482
rect 4277 67430 4329 67482
rect 4341 67430 4393 67482
rect 4405 67430 4457 67482
rect 4469 67430 4521 67482
rect 7477 67430 7529 67482
rect 7541 67430 7593 67482
rect 7605 67430 7657 67482
rect 7669 67430 7721 67482
rect 7733 67430 7785 67482
rect 1768 67371 1820 67380
rect 1768 67337 1777 67371
rect 1777 67337 1811 67371
rect 1811 67337 1820 67371
rect 1768 67328 1820 67337
rect 8392 67328 8444 67380
rect 10140 67328 10192 67380
rect 2964 67192 3016 67244
rect 1860 67167 1912 67176
rect 1860 67133 1869 67167
rect 1869 67133 1903 67167
rect 1903 67133 1912 67167
rect 1860 67124 1912 67133
rect 2504 67124 2556 67176
rect 8300 67235 8352 67244
rect 8300 67201 8309 67235
rect 8309 67201 8343 67235
rect 8343 67201 8352 67235
rect 8300 67192 8352 67201
rect 8944 67192 8996 67244
rect 9128 67167 9180 67176
rect 9128 67133 9137 67167
rect 9137 67133 9171 67167
rect 9171 67133 9180 67167
rect 9128 67124 9180 67133
rect 9680 67124 9732 67176
rect 9496 67056 9548 67108
rect 7380 66988 7432 67040
rect 10048 67031 10100 67040
rect 10048 66997 10057 67031
rect 10057 66997 10091 67031
rect 10091 66997 10100 67031
rect 10048 66988 10100 66997
rect 2582 66886 2634 66938
rect 2646 66886 2698 66938
rect 2710 66886 2762 66938
rect 2774 66886 2826 66938
rect 2838 66886 2890 66938
rect 5845 66886 5897 66938
rect 5909 66886 5961 66938
rect 5973 66886 6025 66938
rect 6037 66886 6089 66938
rect 6101 66886 6153 66938
rect 9109 66886 9161 66938
rect 9173 66886 9225 66938
rect 9237 66886 9289 66938
rect 9301 66886 9353 66938
rect 9365 66886 9417 66938
rect 3424 66648 3476 66700
rect 3608 66648 3660 66700
rect 2136 66623 2188 66632
rect 2136 66589 2145 66623
rect 2145 66589 2179 66623
rect 2179 66589 2188 66623
rect 2136 66580 2188 66589
rect 2504 66580 2556 66632
rect 7012 66580 7064 66632
rect 7196 66623 7248 66632
rect 7196 66589 7205 66623
rect 7205 66589 7239 66623
rect 7239 66589 7248 66623
rect 7196 66580 7248 66589
rect 9036 66580 9088 66632
rect 9404 66623 9456 66632
rect 9404 66589 9413 66623
rect 9413 66589 9447 66623
rect 9447 66589 9456 66623
rect 9404 66580 9456 66589
rect 9680 66623 9732 66632
rect 6276 66512 6328 66564
rect 8024 66512 8076 66564
rect 8944 66512 8996 66564
rect 9680 66589 9689 66623
rect 9689 66589 9723 66623
rect 9723 66589 9732 66623
rect 9680 66580 9732 66589
rect 10140 66555 10192 66564
rect 10140 66521 10149 66555
rect 10149 66521 10183 66555
rect 10183 66521 10192 66555
rect 10140 66512 10192 66521
rect 4213 66342 4265 66394
rect 4277 66342 4329 66394
rect 4341 66342 4393 66394
rect 4405 66342 4457 66394
rect 4469 66342 4521 66394
rect 7477 66342 7529 66394
rect 7541 66342 7593 66394
rect 7605 66342 7657 66394
rect 7669 66342 7721 66394
rect 7733 66342 7785 66394
rect 3056 66172 3108 66224
rect 3148 66172 3200 66224
rect 1768 66147 1820 66156
rect 1768 66113 1777 66147
rect 1777 66113 1811 66147
rect 1811 66113 1820 66147
rect 1768 66104 1820 66113
rect 2504 66104 2556 66156
rect 5632 66104 5684 66156
rect 11704 66104 11756 66156
rect 1860 66036 1912 66088
rect 2964 66036 3016 66088
rect 3608 66036 3660 66088
rect 5172 65968 5224 66020
rect 9496 65900 9548 65952
rect 10048 65943 10100 65952
rect 10048 65909 10057 65943
rect 10057 65909 10091 65943
rect 10091 65909 10100 65943
rect 10048 65900 10100 65909
rect 2582 65798 2634 65850
rect 2646 65798 2698 65850
rect 2710 65798 2762 65850
rect 2774 65798 2826 65850
rect 2838 65798 2890 65850
rect 5845 65798 5897 65850
rect 5909 65798 5961 65850
rect 5973 65798 6025 65850
rect 6037 65798 6089 65850
rect 6101 65798 6153 65850
rect 9109 65798 9161 65850
rect 9173 65798 9225 65850
rect 9237 65798 9289 65850
rect 9301 65798 9353 65850
rect 9365 65798 9417 65850
rect 3056 65696 3108 65748
rect 9036 65628 9088 65680
rect 9588 65560 9640 65612
rect 1584 65535 1636 65544
rect 1584 65501 1593 65535
rect 1593 65501 1627 65535
rect 1627 65501 1636 65535
rect 1584 65492 1636 65501
rect 2228 65535 2280 65544
rect 2228 65501 2237 65535
rect 2237 65501 2271 65535
rect 2271 65501 2280 65535
rect 2228 65492 2280 65501
rect 6736 65492 6788 65544
rect 9496 65535 9548 65544
rect 9496 65501 9505 65535
rect 9505 65501 9539 65535
rect 9539 65501 9548 65535
rect 9496 65492 9548 65501
rect 6552 65424 6604 65476
rect 9864 65424 9916 65476
rect 10600 65424 10652 65476
rect 8944 65356 8996 65408
rect 4213 65254 4265 65306
rect 4277 65254 4329 65306
rect 4341 65254 4393 65306
rect 4405 65254 4457 65306
rect 4469 65254 4521 65306
rect 7477 65254 7529 65306
rect 7541 65254 7593 65306
rect 7605 65254 7657 65306
rect 7669 65254 7721 65306
rect 7733 65254 7785 65306
rect 7380 65152 7432 65204
rect 9496 65152 9548 65204
rect 1860 65059 1912 65068
rect 1860 65025 1869 65059
rect 1869 65025 1903 65059
rect 1903 65025 1912 65059
rect 1860 65016 1912 65025
rect 8116 65016 8168 65068
rect 8760 65059 8812 65068
rect 8760 65025 8769 65059
rect 8769 65025 8803 65059
rect 8803 65025 8812 65059
rect 8760 65016 8812 65025
rect 9588 65016 9640 65068
rect 9864 65059 9916 65068
rect 9864 65025 9873 65059
rect 9873 65025 9907 65059
rect 9907 65025 9916 65059
rect 9864 65016 9916 65025
rect 9680 64880 9732 64932
rect 10048 64923 10100 64932
rect 10048 64889 10057 64923
rect 10057 64889 10091 64923
rect 10091 64889 10100 64923
rect 10048 64880 10100 64889
rect 9496 64812 9548 64864
rect 2582 64710 2634 64762
rect 2646 64710 2698 64762
rect 2710 64710 2762 64762
rect 2774 64710 2826 64762
rect 2838 64710 2890 64762
rect 5845 64710 5897 64762
rect 5909 64710 5961 64762
rect 5973 64710 6025 64762
rect 6037 64710 6089 64762
rect 6101 64710 6153 64762
rect 9109 64710 9161 64762
rect 9173 64710 9225 64762
rect 9237 64710 9289 64762
rect 9301 64710 9353 64762
rect 9365 64710 9417 64762
rect 1400 64447 1452 64456
rect 1400 64413 1409 64447
rect 1409 64413 1443 64447
rect 1443 64413 1452 64447
rect 1400 64404 1452 64413
rect 8392 64404 8444 64456
rect 9496 64447 9548 64456
rect 9496 64413 9505 64447
rect 9505 64413 9539 64447
rect 9539 64413 9548 64447
rect 9496 64404 9548 64413
rect 9680 64447 9732 64456
rect 9680 64413 9689 64447
rect 9689 64413 9723 64447
rect 9723 64413 9732 64447
rect 9680 64404 9732 64413
rect 10416 64336 10468 64388
rect 8852 64268 8904 64320
rect 9496 64268 9548 64320
rect 4213 64166 4265 64218
rect 4277 64166 4329 64218
rect 4341 64166 4393 64218
rect 4405 64166 4457 64218
rect 4469 64166 4521 64218
rect 7477 64166 7529 64218
rect 7541 64166 7593 64218
rect 7605 64166 7657 64218
rect 7669 64166 7721 64218
rect 7733 64166 7785 64218
rect 9036 64064 9088 64116
rect 1032 63928 1084 63980
rect 10140 63971 10192 63980
rect 10140 63937 10149 63971
rect 10149 63937 10183 63971
rect 10183 63937 10192 63971
rect 10140 63928 10192 63937
rect 9588 63860 9640 63912
rect 1768 63724 1820 63776
rect 2582 63622 2634 63674
rect 2646 63622 2698 63674
rect 2710 63622 2762 63674
rect 2774 63622 2826 63674
rect 2838 63622 2890 63674
rect 5845 63622 5897 63674
rect 5909 63622 5961 63674
rect 5973 63622 6025 63674
rect 6037 63622 6089 63674
rect 6101 63622 6153 63674
rect 9109 63622 9161 63674
rect 9173 63622 9225 63674
rect 9237 63622 9289 63674
rect 9301 63622 9353 63674
rect 9365 63622 9417 63674
rect 2596 63495 2648 63504
rect 2596 63461 2605 63495
rect 2605 63461 2639 63495
rect 2639 63461 2648 63495
rect 2596 63452 2648 63461
rect 2964 63427 3016 63436
rect 2964 63393 2973 63427
rect 2973 63393 3007 63427
rect 3007 63393 3016 63427
rect 2964 63384 3016 63393
rect 1400 63359 1452 63368
rect 1400 63325 1409 63359
rect 1409 63325 1443 63359
rect 1443 63325 1452 63359
rect 1400 63316 1452 63325
rect 2504 63316 2556 63368
rect 3608 63384 3660 63436
rect 9496 63359 9548 63368
rect 9496 63325 9505 63359
rect 9505 63325 9539 63359
rect 9539 63325 9548 63359
rect 9496 63316 9548 63325
rect 10232 63316 10284 63368
rect 6460 63248 6512 63300
rect 3148 63180 3200 63232
rect 9496 63180 9548 63232
rect 4213 63078 4265 63130
rect 4277 63078 4329 63130
rect 4341 63078 4393 63130
rect 4405 63078 4457 63130
rect 4469 63078 4521 63130
rect 7477 63078 7529 63130
rect 7541 63078 7593 63130
rect 7605 63078 7657 63130
rect 7669 63078 7721 63130
rect 7733 63078 7785 63130
rect 2320 63019 2372 63028
rect 2320 62985 2329 63019
rect 2329 62985 2363 63019
rect 2363 62985 2372 63019
rect 2320 62976 2372 62985
rect 7380 62976 7432 63028
rect 9036 62976 9088 63028
rect 2228 62772 2280 62824
rect 2504 62815 2556 62824
rect 2504 62781 2513 62815
rect 2513 62781 2547 62815
rect 2547 62781 2556 62815
rect 2504 62772 2556 62781
rect 9588 62840 9640 62892
rect 10140 62883 10192 62892
rect 10140 62849 10149 62883
rect 10149 62849 10183 62883
rect 10183 62849 10192 62883
rect 10140 62840 10192 62849
rect 6184 62704 6236 62756
rect 8484 62772 8536 62824
rect 11428 62772 11480 62824
rect 7380 62679 7432 62688
rect 7380 62645 7389 62679
rect 7389 62645 7423 62679
rect 7423 62645 7432 62679
rect 7380 62636 7432 62645
rect 8116 62704 8168 62756
rect 2582 62534 2634 62586
rect 2646 62534 2698 62586
rect 2710 62534 2762 62586
rect 2774 62534 2826 62586
rect 2838 62534 2890 62586
rect 5845 62534 5897 62586
rect 5909 62534 5961 62586
rect 5973 62534 6025 62586
rect 6037 62534 6089 62586
rect 6101 62534 6153 62586
rect 9109 62534 9161 62586
rect 9173 62534 9225 62586
rect 9237 62534 9289 62586
rect 9301 62534 9353 62586
rect 9365 62534 9417 62586
rect 8668 62432 8720 62484
rect 11244 62364 11296 62416
rect 8484 62296 8536 62348
rect 7104 62228 7156 62280
rect 9312 62271 9364 62280
rect 9312 62237 9321 62271
rect 9321 62237 9355 62271
rect 9355 62237 9364 62271
rect 9312 62228 9364 62237
rect 1860 62203 1912 62212
rect 1860 62169 1869 62203
rect 1869 62169 1903 62203
rect 1903 62169 1912 62203
rect 1860 62160 1912 62169
rect 3516 62160 3568 62212
rect 8208 62092 8260 62144
rect 4213 61990 4265 62042
rect 4277 61990 4329 62042
rect 4341 61990 4393 62042
rect 4405 61990 4457 62042
rect 4469 61990 4521 62042
rect 7477 61990 7529 62042
rect 7541 61990 7593 62042
rect 7605 61990 7657 62042
rect 7669 61990 7721 62042
rect 7733 61990 7785 62042
rect 1400 61752 1452 61804
rect 3608 61616 3660 61668
rect 9588 61548 9640 61600
rect 2582 61446 2634 61498
rect 2646 61446 2698 61498
rect 2710 61446 2762 61498
rect 2774 61446 2826 61498
rect 2838 61446 2890 61498
rect 5845 61446 5897 61498
rect 5909 61446 5961 61498
rect 5973 61446 6025 61498
rect 6037 61446 6089 61498
rect 6101 61446 6153 61498
rect 9109 61446 9161 61498
rect 9173 61446 9225 61498
rect 9237 61446 9289 61498
rect 9301 61446 9353 61498
rect 9365 61446 9417 61498
rect 2228 61251 2280 61260
rect 2228 61217 2237 61251
rect 2237 61217 2271 61251
rect 2271 61217 2280 61251
rect 2228 61208 2280 61217
rect 5356 61208 5408 61260
rect 2320 61183 2372 61192
rect 2320 61149 2329 61183
rect 2329 61149 2363 61183
rect 2363 61149 2372 61183
rect 2320 61140 2372 61149
rect 2504 61183 2556 61192
rect 2504 61149 2513 61183
rect 2513 61149 2547 61183
rect 2547 61149 2556 61183
rect 9404 61183 9456 61192
rect 2504 61140 2556 61149
rect 9404 61149 9413 61183
rect 9413 61149 9447 61183
rect 9447 61149 9456 61183
rect 9404 61140 9456 61149
rect 9496 61183 9548 61192
rect 9496 61149 9505 61183
rect 9505 61149 9539 61183
rect 9539 61149 9548 61183
rect 9496 61140 9548 61149
rect 9680 61183 9732 61192
rect 9680 61149 9689 61183
rect 9689 61149 9723 61183
rect 9723 61149 9732 61183
rect 9680 61140 9732 61149
rect 4988 61072 5040 61124
rect 10508 61072 10560 61124
rect 11336 61047 11388 61056
rect 11336 61013 11345 61047
rect 11345 61013 11379 61047
rect 11379 61013 11388 61047
rect 11336 61004 11388 61013
rect 4213 60902 4265 60954
rect 4277 60902 4329 60954
rect 4341 60902 4393 60954
rect 4405 60902 4457 60954
rect 4469 60902 4521 60954
rect 7477 60902 7529 60954
rect 7541 60902 7593 60954
rect 7605 60902 7657 60954
rect 7669 60902 7721 60954
rect 7733 60902 7785 60954
rect 10968 60936 11020 60988
rect 2044 60843 2096 60852
rect 2044 60809 2053 60843
rect 2053 60809 2087 60843
rect 2087 60809 2096 60843
rect 2044 60800 2096 60809
rect 8116 60800 8168 60852
rect 8300 60800 8352 60852
rect 2504 60732 2556 60784
rect 8668 60775 8720 60784
rect 8668 60741 8677 60775
rect 8677 60741 8711 60775
rect 8711 60741 8720 60775
rect 8668 60732 8720 60741
rect 2780 60707 2832 60716
rect 2780 60673 2789 60707
rect 2789 60673 2823 60707
rect 2823 60673 2832 60707
rect 9312 60707 9364 60716
rect 2780 60664 2832 60673
rect 9312 60673 9321 60707
rect 9321 60673 9355 60707
rect 9355 60673 9364 60707
rect 9312 60664 9364 60673
rect 11428 60843 11480 60852
rect 11428 60809 11437 60843
rect 11437 60809 11471 60843
rect 11471 60809 11480 60843
rect 11428 60800 11480 60809
rect 11796 60843 11848 60852
rect 11244 60775 11296 60784
rect 11244 60741 11253 60775
rect 11253 60741 11287 60775
rect 11287 60741 11296 60775
rect 11796 60809 11805 60843
rect 11805 60809 11839 60843
rect 11839 60809 11848 60843
rect 11796 60800 11848 60809
rect 11244 60732 11296 60741
rect 1676 60596 1728 60648
rect 2044 60639 2096 60648
rect 2044 60605 2053 60639
rect 2053 60605 2087 60639
rect 2087 60605 2096 60639
rect 2044 60596 2096 60605
rect 10232 60596 10284 60648
rect 10968 60596 11020 60648
rect 3976 60528 4028 60580
rect 1584 60503 1636 60512
rect 1584 60469 1593 60503
rect 1593 60469 1627 60503
rect 1627 60469 1636 60503
rect 1584 60460 1636 60469
rect 8760 60503 8812 60512
rect 8760 60469 8769 60503
rect 8769 60469 8803 60503
rect 8803 60469 8812 60503
rect 8760 60460 8812 60469
rect 2582 60358 2634 60410
rect 2646 60358 2698 60410
rect 2710 60358 2762 60410
rect 2774 60358 2826 60410
rect 2838 60358 2890 60410
rect 5845 60358 5897 60410
rect 5909 60358 5961 60410
rect 5973 60358 6025 60410
rect 6037 60358 6089 60410
rect 6101 60358 6153 60410
rect 9109 60358 9161 60410
rect 9173 60358 9225 60410
rect 9237 60358 9289 60410
rect 9301 60358 9353 60410
rect 9365 60358 9417 60410
rect 11520 60299 11572 60308
rect 11520 60265 11529 60299
rect 11529 60265 11563 60299
rect 11563 60265 11572 60299
rect 11520 60256 11572 60265
rect 7104 60188 7156 60240
rect 8208 60163 8260 60172
rect 8208 60129 8217 60163
rect 8217 60129 8251 60163
rect 8251 60129 8260 60163
rect 8208 60120 8260 60129
rect 8484 60120 8536 60172
rect 10048 60052 10100 60104
rect 1860 60027 1912 60036
rect 1860 59993 1869 60027
rect 1869 59993 1903 60027
rect 1903 59993 1912 60027
rect 1860 59984 1912 59993
rect 848 59916 900 59968
rect 7196 59916 7248 59968
rect 4213 59814 4265 59866
rect 4277 59814 4329 59866
rect 4341 59814 4393 59866
rect 4405 59814 4457 59866
rect 4469 59814 4521 59866
rect 7477 59814 7529 59866
rect 7541 59814 7593 59866
rect 7605 59814 7657 59866
rect 7669 59814 7721 59866
rect 7733 59814 7785 59866
rect 7196 59712 7248 59764
rect 8208 59712 8260 59764
rect 9220 59687 9272 59696
rect 9220 59653 9229 59687
rect 9229 59653 9263 59687
rect 9263 59653 9272 59687
rect 9220 59644 9272 59653
rect 1860 59619 1912 59628
rect 1860 59585 1869 59619
rect 1869 59585 1903 59619
rect 1903 59585 1912 59619
rect 1860 59576 1912 59585
rect 9956 59619 10008 59628
rect 9956 59585 9965 59619
rect 9965 59585 9999 59619
rect 9999 59585 10008 59619
rect 9956 59576 10008 59585
rect 10784 59440 10836 59492
rect 664 59372 716 59424
rect 8484 59372 8536 59424
rect 2582 59270 2634 59322
rect 2646 59270 2698 59322
rect 2710 59270 2762 59322
rect 2774 59270 2826 59322
rect 2838 59270 2890 59322
rect 5845 59270 5897 59322
rect 5909 59270 5961 59322
rect 5973 59270 6025 59322
rect 6037 59270 6089 59322
rect 6101 59270 6153 59322
rect 9109 59270 9161 59322
rect 9173 59270 9225 59322
rect 9237 59270 9289 59322
rect 9301 59270 9353 59322
rect 9365 59270 9417 59322
rect 10232 58896 10284 58948
rect 4213 58726 4265 58778
rect 4277 58726 4329 58778
rect 4341 58726 4393 58778
rect 4405 58726 4457 58778
rect 4469 58726 4521 58778
rect 7477 58726 7529 58778
rect 7541 58726 7593 58778
rect 7605 58726 7657 58778
rect 7669 58726 7721 58778
rect 7733 58726 7785 58778
rect 3608 58624 3660 58676
rect 3884 58624 3936 58676
rect 8300 58624 8352 58676
rect 8852 58624 8904 58676
rect 8852 58488 8904 58540
rect 9956 58531 10008 58540
rect 9956 58497 9965 58531
rect 9965 58497 9999 58531
rect 9999 58497 10008 58531
rect 9956 58488 10008 58497
rect 1584 58395 1636 58404
rect 1584 58361 1593 58395
rect 1593 58361 1627 58395
rect 1627 58361 1636 58395
rect 1584 58352 1636 58361
rect 11888 58352 11940 58404
rect 2582 58182 2634 58234
rect 2646 58182 2698 58234
rect 2710 58182 2762 58234
rect 2774 58182 2826 58234
rect 2838 58182 2890 58234
rect 5845 58182 5897 58234
rect 5909 58182 5961 58234
rect 5973 58182 6025 58234
rect 6037 58182 6089 58234
rect 6101 58182 6153 58234
rect 9109 58182 9161 58234
rect 9173 58182 9225 58234
rect 9237 58182 9289 58234
rect 9301 58182 9353 58234
rect 9365 58182 9417 58234
rect 8668 57876 8720 57928
rect 5264 57808 5316 57860
rect 11704 57876 11756 57928
rect 10324 57808 10376 57860
rect 1584 57783 1636 57792
rect 1584 57749 1593 57783
rect 1593 57749 1627 57783
rect 1627 57749 1636 57783
rect 1584 57740 1636 57749
rect 11244 57740 11296 57792
rect 4213 57638 4265 57690
rect 4277 57638 4329 57690
rect 4341 57638 4393 57690
rect 4405 57638 4457 57690
rect 4469 57638 4521 57690
rect 7477 57638 7529 57690
rect 7541 57638 7593 57690
rect 7605 57638 7657 57690
rect 7669 57638 7721 57690
rect 7733 57638 7785 57690
rect 1676 57468 1728 57520
rect 11336 57468 11388 57520
rect 9036 57400 9088 57452
rect 9220 57443 9272 57452
rect 9220 57409 9229 57443
rect 9229 57409 9263 57443
rect 9263 57409 9272 57443
rect 9220 57400 9272 57409
rect 9588 57400 9640 57452
rect 1860 57332 1912 57384
rect 5724 57332 5776 57384
rect 1584 57239 1636 57248
rect 1584 57205 1593 57239
rect 1593 57205 1627 57239
rect 1627 57205 1636 57239
rect 1584 57196 1636 57205
rect 5724 57196 5776 57248
rect 11152 57196 11204 57248
rect 2582 57094 2634 57146
rect 2646 57094 2698 57146
rect 2710 57094 2762 57146
rect 2774 57094 2826 57146
rect 2838 57094 2890 57146
rect 5845 57094 5897 57146
rect 5909 57094 5961 57146
rect 5973 57094 6025 57146
rect 6037 57094 6089 57146
rect 6101 57094 6153 57146
rect 9109 57094 9161 57146
rect 9173 57094 9225 57146
rect 9237 57094 9289 57146
rect 9301 57094 9353 57146
rect 9365 57094 9417 57146
rect 1032 56992 1084 57044
rect 5724 56992 5776 57044
rect 3240 56924 3292 56976
rect 3608 56924 3660 56976
rect 5448 56924 5500 56976
rect 11704 56967 11756 56976
rect 11704 56933 11713 56967
rect 11713 56933 11747 56967
rect 11747 56933 11756 56967
rect 11704 56924 11756 56933
rect 10232 56856 10284 56908
rect 3792 56788 3844 56840
rect 6644 56788 6696 56840
rect 11796 56788 11848 56840
rect 10048 56763 10100 56772
rect 10048 56729 10057 56763
rect 10057 56729 10091 56763
rect 10091 56729 10100 56763
rect 10048 56720 10100 56729
rect 1584 56695 1636 56704
rect 1584 56661 1593 56695
rect 1593 56661 1627 56695
rect 1627 56661 1636 56695
rect 1584 56652 1636 56661
rect 4213 56550 4265 56602
rect 4277 56550 4329 56602
rect 4341 56550 4393 56602
rect 4405 56550 4457 56602
rect 4469 56550 4521 56602
rect 7477 56550 7529 56602
rect 7541 56550 7593 56602
rect 7605 56550 7657 56602
rect 7669 56550 7721 56602
rect 7733 56550 7785 56602
rect 2964 56312 3016 56364
rect 9864 56355 9916 56364
rect 9864 56321 9873 56355
rect 9873 56321 9907 56355
rect 9907 56321 9916 56355
rect 9864 56312 9916 56321
rect 1584 56151 1636 56160
rect 1584 56117 1593 56151
rect 1593 56117 1627 56151
rect 1627 56117 1636 56151
rect 1584 56108 1636 56117
rect 7748 56108 7800 56160
rect 8024 56108 8076 56160
rect 10692 56108 10744 56160
rect 2582 56006 2634 56058
rect 2646 56006 2698 56058
rect 2710 56006 2762 56058
rect 2774 56006 2826 56058
rect 2838 56006 2890 56058
rect 5845 56006 5897 56058
rect 5909 56006 5961 56058
rect 5973 56006 6025 56058
rect 6037 56006 6089 56058
rect 6101 56006 6153 56058
rect 9109 56006 9161 56058
rect 9173 56006 9225 56058
rect 9237 56006 9289 56058
rect 9301 56006 9353 56058
rect 9365 56006 9417 56058
rect 10968 56040 11020 56092
rect 11796 55879 11848 55888
rect 5540 55700 5592 55752
rect 9864 55743 9916 55752
rect 9864 55709 9873 55743
rect 9873 55709 9907 55743
rect 9907 55709 9916 55743
rect 9864 55700 9916 55709
rect 11796 55845 11805 55879
rect 11805 55845 11839 55879
rect 11839 55845 11848 55879
rect 11796 55836 11848 55845
rect 1584 55607 1636 55616
rect 1584 55573 1593 55607
rect 1593 55573 1627 55607
rect 1627 55573 1636 55607
rect 1584 55564 1636 55573
rect 4213 55462 4265 55514
rect 4277 55462 4329 55514
rect 4341 55462 4393 55514
rect 4405 55462 4457 55514
rect 4469 55462 4521 55514
rect 7477 55462 7529 55514
rect 7541 55462 7593 55514
rect 7605 55462 7657 55514
rect 7669 55462 7721 55514
rect 7733 55462 7785 55514
rect 2228 55224 2280 55276
rect 9864 55267 9916 55276
rect 9864 55233 9873 55267
rect 9873 55233 9907 55267
rect 9907 55233 9916 55267
rect 9864 55224 9916 55233
rect 10876 55156 10928 55208
rect 1584 55063 1636 55072
rect 1584 55029 1593 55063
rect 1593 55029 1627 55063
rect 1627 55029 1636 55063
rect 1584 55020 1636 55029
rect 2582 54918 2634 54970
rect 2646 54918 2698 54970
rect 2710 54918 2762 54970
rect 2774 54918 2826 54970
rect 2838 54918 2890 54970
rect 5845 54918 5897 54970
rect 5909 54918 5961 54970
rect 5973 54918 6025 54970
rect 6037 54918 6089 54970
rect 6101 54918 6153 54970
rect 9109 54918 9161 54970
rect 9173 54918 9225 54970
rect 9237 54918 9289 54970
rect 9301 54918 9353 54970
rect 9365 54918 9417 54970
rect 1676 54859 1728 54868
rect 1676 54825 1685 54859
rect 1685 54825 1719 54859
rect 1719 54825 1728 54859
rect 1676 54816 1728 54825
rect 1952 54680 2004 54732
rect 2136 54723 2188 54732
rect 2136 54689 2145 54723
rect 2145 54689 2179 54723
rect 2179 54689 2188 54723
rect 2136 54680 2188 54689
rect 2320 54544 2372 54596
rect 2504 54544 2556 54596
rect 9956 54587 10008 54596
rect 9956 54553 9965 54587
rect 9965 54553 9999 54587
rect 9999 54553 10008 54587
rect 9956 54544 10008 54553
rect 1676 54476 1728 54528
rect 4213 54374 4265 54426
rect 4277 54374 4329 54426
rect 4341 54374 4393 54426
rect 4405 54374 4457 54426
rect 4469 54374 4521 54426
rect 7477 54374 7529 54426
rect 7541 54374 7593 54426
rect 7605 54374 7657 54426
rect 7669 54374 7721 54426
rect 7733 54374 7785 54426
rect 2412 54315 2464 54324
rect 2412 54281 2421 54315
rect 2421 54281 2455 54315
rect 2455 54281 2464 54315
rect 2412 54272 2464 54281
rect 1492 54136 1544 54188
rect 1952 54136 2004 54188
rect 9496 54136 9548 54188
rect 9956 54136 10008 54188
rect 2412 54068 2464 54120
rect 388 53932 440 53984
rect 3056 53932 3108 53984
rect 6552 53932 6604 53984
rect 8668 53932 8720 53984
rect 10232 53932 10284 53984
rect 10416 53932 10468 53984
rect 2582 53830 2634 53882
rect 2646 53830 2698 53882
rect 2710 53830 2762 53882
rect 2774 53830 2826 53882
rect 2838 53830 2890 53882
rect 5845 53830 5897 53882
rect 5909 53830 5961 53882
rect 5973 53830 6025 53882
rect 6037 53830 6089 53882
rect 6101 53830 6153 53882
rect 9109 53830 9161 53882
rect 9173 53830 9225 53882
rect 9237 53830 9289 53882
rect 9301 53830 9353 53882
rect 9365 53830 9417 53882
rect 1584 53771 1636 53780
rect 1584 53737 1593 53771
rect 1593 53737 1627 53771
rect 1627 53737 1636 53771
rect 1584 53728 1636 53737
rect 10140 53592 10192 53644
rect 1492 53524 1544 53576
rect 9588 53524 9640 53576
rect 9864 53567 9916 53576
rect 9864 53533 9873 53567
rect 9873 53533 9907 53567
rect 9907 53533 9916 53567
rect 9864 53524 9916 53533
rect 8576 53388 8628 53440
rect 10048 53431 10100 53440
rect 10048 53397 10057 53431
rect 10057 53397 10091 53431
rect 10091 53397 10100 53431
rect 10048 53388 10100 53397
rect 10140 53388 10192 53440
rect 4213 53286 4265 53338
rect 4277 53286 4329 53338
rect 4341 53286 4393 53338
rect 4405 53286 4457 53338
rect 4469 53286 4521 53338
rect 7477 53286 7529 53338
rect 7541 53286 7593 53338
rect 7605 53286 7657 53338
rect 7669 53286 7721 53338
rect 7733 53286 7785 53338
rect 1584 53227 1636 53236
rect 1584 53193 1593 53227
rect 1593 53193 1627 53227
rect 1627 53193 1636 53227
rect 1584 53184 1636 53193
rect 11520 53184 11572 53236
rect 10968 53116 11020 53168
rect 2504 53048 2556 53100
rect 9772 53091 9824 53100
rect 9772 53057 9781 53091
rect 9781 53057 9815 53091
rect 9815 53057 9824 53091
rect 9772 53048 9824 53057
rect 11520 53048 11572 53100
rect 10232 52980 10284 53032
rect 11888 53023 11940 53032
rect 11888 52989 11897 53023
rect 11897 52989 11931 53023
rect 11931 52989 11940 53023
rect 11888 52980 11940 52989
rect 11244 52844 11296 52896
rect 2582 52742 2634 52794
rect 2646 52742 2698 52794
rect 2710 52742 2762 52794
rect 2774 52742 2826 52794
rect 2838 52742 2890 52794
rect 5845 52742 5897 52794
rect 5909 52742 5961 52794
rect 5973 52742 6025 52794
rect 6037 52742 6089 52794
rect 6101 52742 6153 52794
rect 9109 52742 9161 52794
rect 9173 52742 9225 52794
rect 9237 52742 9289 52794
rect 9301 52742 9353 52794
rect 9365 52742 9417 52794
rect 11428 52640 11480 52692
rect 2780 52615 2832 52624
rect 2780 52581 2789 52615
rect 2789 52581 2823 52615
rect 2823 52581 2832 52615
rect 2780 52572 2832 52581
rect 4712 52572 4764 52624
rect 1676 52436 1728 52488
rect 2412 52436 2464 52488
rect 2964 52479 3016 52488
rect 2964 52445 2973 52479
rect 2973 52445 3007 52479
rect 3007 52445 3016 52479
rect 2964 52436 3016 52445
rect 9128 52479 9180 52488
rect 9128 52445 9137 52479
rect 9137 52445 9171 52479
rect 9171 52445 9180 52479
rect 9128 52436 9180 52445
rect 2136 52411 2188 52420
rect 2136 52377 2145 52411
rect 2145 52377 2179 52411
rect 2179 52377 2188 52411
rect 2136 52368 2188 52377
rect 10692 52300 10744 52352
rect 4213 52198 4265 52250
rect 4277 52198 4329 52250
rect 4341 52198 4393 52250
rect 4405 52198 4457 52250
rect 4469 52198 4521 52250
rect 7477 52198 7529 52250
rect 7541 52198 7593 52250
rect 7605 52198 7657 52250
rect 7669 52198 7721 52250
rect 7733 52198 7785 52250
rect 1860 52096 1912 52148
rect 1860 52003 1912 52012
rect 1860 51969 1869 52003
rect 1869 51969 1903 52003
rect 1903 51969 1912 52003
rect 1860 51960 1912 51969
rect 9496 51960 9548 52012
rect 9864 52003 9916 52012
rect 9864 51969 9873 52003
rect 9873 51969 9907 52003
rect 9907 51969 9916 52003
rect 9864 51960 9916 51969
rect 6828 51756 6880 51808
rect 10048 51799 10100 51808
rect 10048 51765 10057 51799
rect 10057 51765 10091 51799
rect 10091 51765 10100 51799
rect 10048 51756 10100 51765
rect 2582 51654 2634 51706
rect 2646 51654 2698 51706
rect 2710 51654 2762 51706
rect 2774 51654 2826 51706
rect 2838 51654 2890 51706
rect 5845 51654 5897 51706
rect 5909 51654 5961 51706
rect 5973 51654 6025 51706
rect 6037 51654 6089 51706
rect 6101 51654 6153 51706
rect 9109 51654 9161 51706
rect 9173 51654 9225 51706
rect 9237 51654 9289 51706
rect 9301 51654 9353 51706
rect 9365 51654 9417 51706
rect 6644 51552 6696 51604
rect 8852 51552 8904 51604
rect 10876 51595 10928 51604
rect 10876 51561 10885 51595
rect 10885 51561 10919 51595
rect 10919 51561 10928 51595
rect 10876 51552 10928 51561
rect 2596 51484 2648 51536
rect 9588 51484 9640 51536
rect 2412 51416 2464 51468
rect 10232 51416 10284 51468
rect 10876 51416 10928 51468
rect 1400 51391 1452 51400
rect 1400 51357 1409 51391
rect 1409 51357 1443 51391
rect 1443 51357 1452 51391
rect 1400 51348 1452 51357
rect 10968 51391 11020 51400
rect 10968 51357 10977 51391
rect 10977 51357 11011 51391
rect 11011 51357 11020 51391
rect 10968 51348 11020 51357
rect 11060 51391 11112 51400
rect 11060 51357 11069 51391
rect 11069 51357 11103 51391
rect 11103 51357 11112 51391
rect 11060 51348 11112 51357
rect 9496 51280 9548 51332
rect 6644 51212 6696 51264
rect 8208 51212 8260 51264
rect 9680 51212 9732 51264
rect 10784 51212 10836 51264
rect 4213 51110 4265 51162
rect 4277 51110 4329 51162
rect 4341 51110 4393 51162
rect 4405 51110 4457 51162
rect 4469 51110 4521 51162
rect 7477 51110 7529 51162
rect 7541 51110 7593 51162
rect 7605 51110 7657 51162
rect 7669 51110 7721 51162
rect 7733 51110 7785 51162
rect 10968 51144 11020 51196
rect 11336 51416 11388 51468
rect 11796 51391 11848 51400
rect 11796 51357 11805 51391
rect 11805 51357 11839 51391
rect 11839 51357 11848 51391
rect 11796 51348 11848 51357
rect 11336 51076 11388 51128
rect 940 51008 992 51060
rect 2504 51051 2556 51060
rect 2504 51017 2513 51051
rect 2513 51017 2547 51051
rect 2547 51017 2556 51051
rect 2504 51008 2556 51017
rect 3148 51008 3200 51060
rect 7012 51008 7064 51060
rect 1860 50915 1912 50924
rect 1860 50881 1869 50915
rect 1869 50881 1903 50915
rect 1903 50881 1912 50915
rect 1860 50872 1912 50881
rect 480 50804 532 50856
rect 7288 51008 7340 51060
rect 7380 51008 7432 51060
rect 8300 51008 8352 51060
rect 10968 51008 11020 51060
rect 9772 50940 9824 50992
rect 10692 50940 10744 50992
rect 8300 50872 8352 50924
rect 8944 50872 8996 50924
rect 11704 50983 11756 50992
rect 11704 50949 11713 50983
rect 11713 50949 11747 50983
rect 11747 50949 11756 50983
rect 11704 50940 11756 50949
rect 3608 50804 3660 50856
rect 7196 50804 7248 50856
rect 7288 50804 7340 50856
rect 7380 50804 7432 50856
rect 8852 50804 8904 50856
rect 10232 50804 10284 50856
rect 11152 50804 11204 50856
rect 9496 50668 9548 50720
rect 9588 50668 9640 50720
rect 10784 50668 10836 50720
rect 11428 50668 11480 50720
rect 2582 50566 2634 50618
rect 2646 50566 2698 50618
rect 2710 50566 2762 50618
rect 2774 50566 2826 50618
rect 2838 50566 2890 50618
rect 5845 50566 5897 50618
rect 5909 50566 5961 50618
rect 5973 50566 6025 50618
rect 6037 50566 6089 50618
rect 6101 50566 6153 50618
rect 9109 50566 9161 50618
rect 9173 50566 9225 50618
rect 9237 50566 9289 50618
rect 9301 50566 9353 50618
rect 9365 50566 9417 50618
rect 11336 50600 11388 50652
rect 1216 50464 1268 50516
rect 9036 50464 9088 50516
rect 9956 50396 10008 50448
rect 11888 50396 11940 50448
rect 9496 50328 9548 50380
rect 9864 50328 9916 50380
rect 11796 50328 11848 50380
rect 8116 50303 8168 50312
rect 8116 50269 8125 50303
rect 8125 50269 8159 50303
rect 8159 50269 8168 50303
rect 8116 50260 8168 50269
rect 1860 50235 1912 50244
rect 1860 50201 1869 50235
rect 1869 50201 1903 50235
rect 1903 50201 1912 50235
rect 1860 50192 1912 50201
rect 3056 50192 3108 50244
rect 5264 50192 5316 50244
rect 8392 50124 8444 50176
rect 8760 50124 8812 50176
rect 9036 50124 9088 50176
rect 9496 50167 9548 50176
rect 9496 50133 9505 50167
rect 9505 50133 9539 50167
rect 9539 50133 9548 50167
rect 9496 50124 9548 50133
rect 9680 50124 9732 50176
rect 4213 50022 4265 50074
rect 4277 50022 4329 50074
rect 4341 50022 4393 50074
rect 4405 50022 4457 50074
rect 4469 50022 4521 50074
rect 7477 50022 7529 50074
rect 7541 50022 7593 50074
rect 7605 50022 7657 50074
rect 7669 50022 7721 50074
rect 7733 50022 7785 50074
rect 5264 49920 5316 49972
rect 9956 49963 10008 49972
rect 9956 49929 9965 49963
rect 9965 49929 9999 49963
rect 9999 49929 10008 49963
rect 9956 49920 10008 49929
rect 6552 49852 6604 49904
rect 6828 49852 6880 49904
rect 8668 49827 8720 49836
rect 8668 49793 8677 49827
rect 8677 49793 8711 49827
rect 8711 49793 8720 49827
rect 8668 49784 8720 49793
rect 9864 49784 9916 49836
rect 11244 49784 11296 49836
rect 3608 49716 3660 49768
rect 4160 49716 4212 49768
rect 6828 49716 6880 49768
rect 2412 49648 2464 49700
rect 7012 49648 7064 49700
rect 8668 49648 8720 49700
rect 9128 49648 9180 49700
rect 11796 49716 11848 49768
rect 2320 49580 2372 49632
rect 7196 49580 7248 49632
rect 2582 49478 2634 49530
rect 2646 49478 2698 49530
rect 2710 49478 2762 49530
rect 2774 49478 2826 49530
rect 2838 49478 2890 49530
rect 5845 49478 5897 49530
rect 5909 49478 5961 49530
rect 5973 49478 6025 49530
rect 6037 49478 6089 49530
rect 6101 49478 6153 49530
rect 9109 49478 9161 49530
rect 9173 49478 9225 49530
rect 9237 49478 9289 49530
rect 9301 49478 9353 49530
rect 9365 49478 9417 49530
rect 3792 49376 3844 49428
rect 6644 49376 6696 49428
rect 8944 49376 8996 49428
rect 4068 49308 4120 49360
rect 7196 49240 7248 49292
rect 9772 49308 9824 49360
rect 10968 49351 11020 49360
rect 10968 49317 10977 49351
rect 10977 49317 11011 49351
rect 11011 49317 11020 49351
rect 10968 49308 11020 49317
rect 1860 49215 1912 49224
rect 1860 49181 1869 49215
rect 1869 49181 1903 49215
rect 1903 49181 1912 49215
rect 1860 49172 1912 49181
rect 8208 49172 8260 49224
rect 9588 49240 9640 49292
rect 9404 49172 9456 49224
rect 572 49036 624 49088
rect 11152 49036 11204 49088
rect 4213 48934 4265 48986
rect 4277 48934 4329 48986
rect 4341 48934 4393 48986
rect 4405 48934 4457 48986
rect 4469 48934 4521 48986
rect 7477 48934 7529 48986
rect 7541 48934 7593 48986
rect 7605 48934 7657 48986
rect 7669 48934 7721 48986
rect 7733 48934 7785 48986
rect 9496 48832 9548 48884
rect 5080 48764 5132 48816
rect 1860 48739 1912 48748
rect 1860 48705 1869 48739
rect 1869 48705 1903 48739
rect 1903 48705 1912 48739
rect 1860 48696 1912 48705
rect 8208 48696 8260 48748
rect 8944 48696 8996 48748
rect 9404 48696 9456 48748
rect 9956 48696 10008 48748
rect 1584 48628 1636 48680
rect 8852 48628 8904 48680
rect 10784 48628 10836 48680
rect 2582 48390 2634 48442
rect 2646 48390 2698 48442
rect 2710 48390 2762 48442
rect 2774 48390 2826 48442
rect 2838 48390 2890 48442
rect 5845 48390 5897 48442
rect 5909 48390 5961 48442
rect 5973 48390 6025 48442
rect 6037 48390 6089 48442
rect 6101 48390 6153 48442
rect 9109 48390 9161 48442
rect 9173 48390 9225 48442
rect 9237 48390 9289 48442
rect 9301 48390 9353 48442
rect 9365 48390 9417 48442
rect 5356 48288 5408 48340
rect 8852 48288 8904 48340
rect 9036 48288 9088 48340
rect 2044 48263 2096 48272
rect 2044 48229 2053 48263
rect 2053 48229 2087 48263
rect 2087 48229 2096 48263
rect 2044 48220 2096 48229
rect 2136 48220 2188 48272
rect 4712 48152 4764 48204
rect 8760 48152 8812 48204
rect 9036 48152 9088 48204
rect 5264 48084 5316 48136
rect 8208 48084 8260 48136
rect 8852 48084 8904 48136
rect 9588 48220 9640 48272
rect 9496 48084 9548 48136
rect 9956 48084 10008 48136
rect 11244 48084 11296 48136
rect 11612 48084 11664 48136
rect 1860 48059 1912 48068
rect 1860 48025 1869 48059
rect 1869 48025 1903 48059
rect 1903 48025 1912 48059
rect 1860 48016 1912 48025
rect 4712 48016 4764 48068
rect 9680 47948 9732 48000
rect 11612 47991 11664 48000
rect 11612 47957 11621 47991
rect 11621 47957 11655 47991
rect 11655 47957 11664 47991
rect 11612 47948 11664 47957
rect 4213 47846 4265 47898
rect 4277 47846 4329 47898
rect 4341 47846 4393 47898
rect 4405 47846 4457 47898
rect 4469 47846 4521 47898
rect 7477 47846 7529 47898
rect 7541 47846 7593 47898
rect 7605 47846 7657 47898
rect 7669 47846 7721 47898
rect 7733 47846 7785 47898
rect 1952 47787 2004 47796
rect 1952 47753 1961 47787
rect 1961 47753 1995 47787
rect 1995 47753 2004 47787
rect 1952 47744 2004 47753
rect 2228 47744 2280 47796
rect 5080 47787 5132 47796
rect 5080 47753 5089 47787
rect 5089 47753 5123 47787
rect 5123 47753 5132 47787
rect 5080 47744 5132 47753
rect 9220 47744 9272 47796
rect 10048 47744 10100 47796
rect 3608 47676 3660 47728
rect 9680 47719 9732 47728
rect 1860 47651 1912 47660
rect 1860 47617 1869 47651
rect 1869 47617 1903 47651
rect 1903 47617 1912 47651
rect 1860 47608 1912 47617
rect 756 47540 808 47592
rect 4712 47540 4764 47592
rect 2872 47472 2924 47524
rect 3608 47472 3660 47524
rect 4712 47404 4764 47456
rect 9680 47685 9689 47719
rect 9689 47685 9723 47719
rect 9723 47685 9732 47719
rect 9680 47676 9732 47685
rect 9588 47608 9640 47660
rect 9864 47608 9916 47660
rect 10232 47608 10284 47660
rect 9496 47540 9548 47592
rect 9956 47583 10008 47592
rect 9956 47549 9965 47583
rect 9965 47549 9999 47583
rect 9999 47549 10008 47583
rect 9956 47540 10008 47549
rect 5724 47404 5776 47456
rect 8668 47447 8720 47456
rect 8668 47413 8677 47447
rect 8677 47413 8711 47447
rect 8711 47413 8720 47447
rect 8668 47404 8720 47413
rect 10048 47404 10100 47456
rect 2582 47302 2634 47354
rect 2646 47302 2698 47354
rect 2710 47302 2762 47354
rect 2774 47302 2826 47354
rect 2838 47302 2890 47354
rect 5845 47302 5897 47354
rect 5909 47302 5961 47354
rect 5973 47302 6025 47354
rect 6037 47302 6089 47354
rect 6101 47302 6153 47354
rect 9109 47302 9161 47354
rect 9173 47302 9225 47354
rect 9237 47302 9289 47354
rect 9301 47302 9353 47354
rect 9365 47302 9417 47354
rect 1124 47200 1176 47252
rect 4068 47200 4120 47252
rect 10876 47200 10928 47252
rect 9772 47132 9824 47184
rect 6644 47064 6696 47116
rect 8852 47064 8904 47116
rect 9404 47064 9456 47116
rect 9956 47107 10008 47116
rect 9956 47073 9965 47107
rect 9965 47073 9999 47107
rect 9999 47073 10008 47107
rect 9956 47064 10008 47073
rect 8208 46996 8260 47048
rect 1860 46971 1912 46980
rect 1860 46937 1869 46971
rect 1869 46937 1903 46971
rect 1903 46937 1912 46971
rect 1860 46928 1912 46937
rect 8668 46928 8720 46980
rect 9680 46860 9732 46912
rect 4213 46758 4265 46810
rect 4277 46758 4329 46810
rect 4341 46758 4393 46810
rect 4405 46758 4457 46810
rect 4469 46758 4521 46810
rect 7477 46758 7529 46810
rect 7541 46758 7593 46810
rect 7605 46758 7657 46810
rect 7669 46758 7721 46810
rect 7733 46758 7785 46810
rect 5540 46656 5592 46708
rect 9772 46699 9824 46708
rect 9772 46665 9781 46699
rect 9781 46665 9815 46699
rect 9815 46665 9824 46699
rect 9772 46656 9824 46665
rect 4068 46588 4120 46640
rect 5080 46563 5132 46572
rect 5080 46529 5089 46563
rect 5089 46529 5123 46563
rect 5123 46529 5132 46563
rect 5080 46520 5132 46529
rect 5724 46588 5776 46640
rect 8116 46588 8168 46640
rect 11244 46520 11296 46572
rect 4712 46452 4764 46504
rect 5724 46495 5776 46504
rect 5724 46461 5733 46495
rect 5733 46461 5767 46495
rect 5767 46461 5776 46495
rect 5724 46452 5776 46461
rect 9404 46452 9456 46504
rect 9496 46452 9548 46504
rect 8024 46384 8076 46436
rect 8576 46384 8628 46436
rect 8852 46384 8904 46436
rect 9588 46384 9640 46436
rect 9956 46316 10008 46368
rect 2582 46214 2634 46266
rect 2646 46214 2698 46266
rect 2710 46214 2762 46266
rect 2774 46214 2826 46266
rect 2838 46214 2890 46266
rect 5845 46214 5897 46266
rect 5909 46214 5961 46266
rect 5973 46214 6025 46266
rect 6037 46214 6089 46266
rect 6101 46214 6153 46266
rect 9109 46214 9161 46266
rect 9173 46214 9225 46266
rect 9237 46214 9289 46266
rect 9301 46214 9353 46266
rect 9365 46214 9417 46266
rect 1308 46112 1360 46164
rect 7012 46112 7064 46164
rect 10232 46112 10284 46164
rect 10416 46112 10468 46164
rect 8668 46044 8720 46096
rect 9588 45976 9640 46028
rect 1860 45951 1912 45960
rect 1860 45917 1869 45951
rect 1869 45917 1903 45951
rect 1903 45917 1912 45951
rect 1860 45908 1912 45917
rect 6920 45908 6972 45960
rect 7012 45908 7064 45960
rect 8208 45908 8260 45960
rect 9588 45840 9640 45892
rect 10416 45840 10468 45892
rect 9956 45815 10008 45824
rect 9956 45781 9965 45815
rect 9965 45781 9999 45815
rect 9999 45781 10008 45815
rect 9956 45772 10008 45781
rect 4213 45670 4265 45722
rect 4277 45670 4329 45722
rect 4341 45670 4393 45722
rect 4405 45670 4457 45722
rect 4469 45670 4521 45722
rect 7477 45670 7529 45722
rect 7541 45670 7593 45722
rect 7605 45670 7657 45722
rect 7669 45670 7721 45722
rect 7733 45670 7785 45722
rect 3884 45568 3936 45620
rect 5172 45568 5224 45620
rect 9956 45568 10008 45620
rect 11704 45568 11756 45620
rect 1952 45500 2004 45552
rect 2320 45500 2372 45552
rect 4712 45500 4764 45552
rect 10048 45500 10100 45552
rect 1400 45475 1452 45484
rect 1400 45441 1409 45475
rect 1409 45441 1443 45475
rect 1443 45441 1452 45475
rect 1400 45432 1452 45441
rect 4068 45432 4120 45484
rect 8208 45432 8260 45484
rect 10968 45432 11020 45484
rect 11704 45432 11756 45484
rect 1768 45364 1820 45416
rect 2228 45364 2280 45416
rect 4160 45364 4212 45416
rect 1492 45296 1544 45348
rect 8760 45296 8812 45348
rect 9588 45296 9640 45348
rect 7288 45228 7340 45280
rect 11244 45228 11296 45280
rect 2582 45126 2634 45178
rect 2646 45126 2698 45178
rect 2710 45126 2762 45178
rect 2774 45126 2826 45178
rect 2838 45126 2890 45178
rect 5845 45126 5897 45178
rect 5909 45126 5961 45178
rect 5973 45126 6025 45178
rect 6037 45126 6089 45178
rect 6101 45126 6153 45178
rect 9109 45126 9161 45178
rect 9173 45126 9225 45178
rect 9237 45126 9289 45178
rect 9301 45126 9353 45178
rect 9365 45126 9417 45178
rect 1584 45024 1636 45076
rect 1768 45024 1820 45076
rect 9588 45024 9640 45076
rect 9864 45024 9916 45076
rect 3332 44956 3384 45008
rect 3332 44820 3384 44872
rect 4160 44820 4212 44872
rect 9404 44863 9456 44872
rect 9404 44829 9413 44863
rect 9413 44829 9447 44863
rect 9447 44829 9456 44863
rect 9404 44820 9456 44829
rect 9772 44888 9824 44940
rect 9956 44820 10008 44872
rect 10416 44820 10468 44872
rect 1860 44795 1912 44804
rect 1860 44761 1869 44795
rect 1869 44761 1903 44795
rect 1903 44761 1912 44795
rect 1860 44752 1912 44761
rect 10140 44795 10192 44804
rect 10140 44761 10149 44795
rect 10149 44761 10183 44795
rect 10183 44761 10192 44795
rect 10140 44752 10192 44761
rect 5632 44684 5684 44736
rect 6368 44684 6420 44736
rect 7288 44684 7340 44736
rect 8392 44684 8444 44736
rect 4213 44582 4265 44634
rect 4277 44582 4329 44634
rect 4341 44582 4393 44634
rect 4405 44582 4457 44634
rect 4469 44582 4521 44634
rect 7477 44582 7529 44634
rect 7541 44582 7593 44634
rect 7605 44582 7657 44634
rect 7669 44582 7721 44634
rect 7733 44582 7785 44634
rect 9588 44480 9640 44532
rect 10140 44480 10192 44532
rect 3240 44412 3292 44464
rect 8208 44412 8260 44464
rect 1860 44387 1912 44396
rect 1860 44353 1869 44387
rect 1869 44353 1903 44387
rect 1903 44353 1912 44387
rect 1860 44344 1912 44353
rect 1584 44276 1636 44328
rect 2504 44276 2556 44328
rect 2044 44208 2096 44260
rect 5080 44208 5132 44260
rect 9220 44344 9272 44396
rect 9404 44319 9456 44328
rect 9404 44285 9414 44319
rect 9414 44285 9448 44319
rect 9448 44285 9456 44319
rect 9956 44344 10008 44396
rect 9404 44276 9456 44285
rect 10048 44276 10100 44328
rect 2320 44140 2372 44192
rect 3976 44140 4028 44192
rect 8392 44140 8444 44192
rect 2582 44038 2634 44090
rect 2646 44038 2698 44090
rect 2710 44038 2762 44090
rect 2774 44038 2826 44090
rect 2838 44038 2890 44090
rect 5845 44038 5897 44090
rect 5909 44038 5961 44090
rect 5973 44038 6025 44090
rect 6037 44038 6089 44090
rect 6101 44038 6153 44090
rect 9109 44038 9161 44090
rect 9173 44038 9225 44090
rect 9237 44038 9289 44090
rect 9301 44038 9353 44090
rect 9365 44038 9417 44090
rect 388 43936 440 43988
rect 1492 43936 1544 43988
rect 7564 43936 7616 43988
rect 11152 43936 11204 43988
rect 848 43868 900 43920
rect 2504 43868 2556 43920
rect 4068 43775 4120 43784
rect 4068 43741 4077 43775
rect 4077 43741 4111 43775
rect 4111 43741 4120 43775
rect 4068 43732 4120 43741
rect 4712 43800 4764 43852
rect 8208 43843 8260 43852
rect 8208 43809 8217 43843
rect 8217 43809 8251 43843
rect 8251 43809 8260 43843
rect 8208 43800 8260 43809
rect 5080 43732 5132 43784
rect 8116 43732 8168 43784
rect 1216 43664 1268 43716
rect 4712 43596 4764 43648
rect 5356 43596 5408 43648
rect 7288 43596 7340 43648
rect 11612 43732 11664 43784
rect 10140 43707 10192 43716
rect 10140 43673 10149 43707
rect 10149 43673 10183 43707
rect 10183 43673 10192 43707
rect 10140 43664 10192 43673
rect 11336 43664 11388 43716
rect 9680 43596 9732 43648
rect 10416 43596 10468 43648
rect 11612 43596 11664 43648
rect 4213 43494 4265 43546
rect 4277 43494 4329 43546
rect 4341 43494 4393 43546
rect 4405 43494 4457 43546
rect 4469 43494 4521 43546
rect 7477 43494 7529 43546
rect 7541 43494 7593 43546
rect 7605 43494 7657 43546
rect 7669 43494 7721 43546
rect 7733 43494 7785 43546
rect 6920 43392 6972 43444
rect 8300 43392 8352 43444
rect 9680 43392 9732 43444
rect 9864 43392 9916 43444
rect 3608 43324 3660 43376
rect 3976 43324 4028 43376
rect 5356 43324 5408 43376
rect 6644 43324 6696 43376
rect 1860 43299 1912 43308
rect 1860 43265 1869 43299
rect 1869 43265 1903 43299
rect 1903 43265 1912 43299
rect 1860 43256 1912 43265
rect 6368 43256 6420 43308
rect 8576 43324 8628 43376
rect 9128 43299 9180 43308
rect 9128 43265 9137 43299
rect 9137 43265 9171 43299
rect 9171 43265 9180 43299
rect 9128 43256 9180 43265
rect 9864 43299 9916 43308
rect 9864 43265 9873 43299
rect 9873 43265 9907 43299
rect 9907 43265 9916 43299
rect 9864 43256 9916 43265
rect 9956 43256 10008 43308
rect 10692 43256 10744 43308
rect 10968 43188 11020 43240
rect 11060 43188 11112 43240
rect 11336 43188 11388 43240
rect 1124 43120 1176 43172
rect 10140 43120 10192 43172
rect 8576 43095 8628 43104
rect 8576 43061 8585 43095
rect 8585 43061 8619 43095
rect 8619 43061 8628 43095
rect 8576 43052 8628 43061
rect 11060 43052 11112 43104
rect 2582 42950 2634 43002
rect 2646 42950 2698 43002
rect 2710 42950 2762 43002
rect 2774 42950 2826 43002
rect 2838 42950 2890 43002
rect 5845 42950 5897 43002
rect 5909 42950 5961 43002
rect 5973 42950 6025 43002
rect 6037 42950 6089 43002
rect 6101 42950 6153 43002
rect 9109 42950 9161 43002
rect 9173 42950 9225 43002
rect 9237 42950 9289 43002
rect 9301 42950 9353 43002
rect 9365 42950 9417 43002
rect 4068 42848 4120 42900
rect 6828 42848 6880 42900
rect 10692 42848 10744 42900
rect 1400 42687 1452 42696
rect 1400 42653 1409 42687
rect 1409 42653 1443 42687
rect 1443 42653 1452 42687
rect 1400 42644 1452 42653
rect 6368 42712 6420 42764
rect 10140 42780 10192 42832
rect 6828 42712 6880 42764
rect 6920 42712 6972 42764
rect 3608 42644 3660 42696
rect 3976 42576 4028 42628
rect 6552 42576 6604 42628
rect 3516 42508 3568 42560
rect 6368 42508 6420 42560
rect 8208 42576 8260 42628
rect 8576 42576 8628 42628
rect 9956 42619 10008 42628
rect 9956 42585 9965 42619
rect 9965 42585 9999 42619
rect 9999 42585 10008 42619
rect 9956 42576 10008 42585
rect 6920 42508 6972 42560
rect 11152 42712 11204 42764
rect 11704 42712 11756 42764
rect 11704 42508 11756 42560
rect 4213 42406 4265 42458
rect 4277 42406 4329 42458
rect 4341 42406 4393 42458
rect 4405 42406 4457 42458
rect 4469 42406 4521 42458
rect 7477 42406 7529 42458
rect 7541 42406 7593 42458
rect 7605 42406 7657 42458
rect 7669 42406 7721 42458
rect 7733 42406 7785 42458
rect 1584 42347 1636 42356
rect 1584 42313 1593 42347
rect 1593 42313 1627 42347
rect 1627 42313 1636 42347
rect 1584 42304 1636 42313
rect 5080 42236 5132 42288
rect 6368 42236 6420 42288
rect 6552 42236 6604 42288
rect 6920 42236 6972 42288
rect 11152 42236 11204 42288
rect 1400 42211 1452 42220
rect 1400 42177 1409 42211
rect 1409 42177 1443 42211
rect 1443 42177 1452 42211
rect 1400 42168 1452 42177
rect 3240 42168 3292 42220
rect 6092 42168 6144 42220
rect 9128 42211 9180 42220
rect 9128 42177 9137 42211
rect 9137 42177 9171 42211
rect 9171 42177 9180 42211
rect 9128 42168 9180 42177
rect 9956 42211 10008 42220
rect 9956 42177 9965 42211
rect 9965 42177 9999 42211
rect 9999 42177 10008 42211
rect 9956 42168 10008 42177
rect 10140 42168 10192 42220
rect 5172 42143 5224 42152
rect 5172 42109 5181 42143
rect 5181 42109 5215 42143
rect 5215 42109 5224 42143
rect 5172 42100 5224 42109
rect 8208 42032 8260 42084
rect 6368 41964 6420 42016
rect 2582 41862 2634 41914
rect 2646 41862 2698 41914
rect 2710 41862 2762 41914
rect 2774 41862 2826 41914
rect 2838 41862 2890 41914
rect 5845 41862 5897 41914
rect 5909 41862 5961 41914
rect 5973 41862 6025 41914
rect 6037 41862 6089 41914
rect 6101 41862 6153 41914
rect 9109 41862 9161 41914
rect 9173 41862 9225 41914
rect 9237 41862 9289 41914
rect 9301 41862 9353 41914
rect 9365 41862 9417 41914
rect 2412 41760 2464 41812
rect 940 41692 992 41744
rect 6368 41692 6420 41744
rect 8944 41692 8996 41744
rect 9404 41692 9456 41744
rect 3516 41624 3568 41676
rect 10140 41624 10192 41676
rect 1400 41599 1452 41608
rect 1400 41565 1409 41599
rect 1409 41565 1443 41599
rect 1443 41565 1452 41599
rect 1400 41556 1452 41565
rect 3792 41556 3844 41608
rect 9864 41556 9916 41608
rect 10692 41556 10744 41608
rect 11336 41828 11388 41880
rect 11336 41692 11388 41744
rect 11612 41828 11664 41880
rect 11888 41964 11940 42016
rect 11152 41556 11204 41608
rect 3332 41488 3384 41540
rect 5448 41488 5500 41540
rect 8576 41488 8628 41540
rect 9956 41531 10008 41540
rect 9956 41497 9965 41531
rect 9965 41497 9999 41531
rect 9999 41497 10008 41531
rect 9956 41488 10008 41497
rect 10140 41488 10192 41540
rect 10784 41488 10836 41540
rect 3792 41420 3844 41472
rect 6920 41420 6972 41472
rect 8760 41420 8812 41472
rect 11888 41488 11940 41540
rect 11244 41420 11296 41472
rect 4213 41318 4265 41370
rect 4277 41318 4329 41370
rect 4341 41318 4393 41370
rect 4405 41318 4457 41370
rect 4469 41318 4521 41370
rect 7477 41318 7529 41370
rect 7541 41318 7593 41370
rect 7605 41318 7657 41370
rect 7669 41318 7721 41370
rect 7733 41318 7785 41370
rect 11060 41284 11112 41336
rect 11152 41284 11204 41336
rect 2504 41216 2556 41268
rect 5540 41216 5592 41268
rect 2136 41148 2188 41200
rect 7472 41148 7524 41200
rect 11060 41148 11112 41200
rect 1860 41123 1912 41132
rect 1860 41089 1869 41123
rect 1869 41089 1903 41123
rect 1903 41089 1912 41123
rect 1860 41080 1912 41089
rect 6460 41080 6512 41132
rect 6828 41080 6880 41132
rect 9956 41123 10008 41132
rect 9956 41089 9965 41123
rect 9965 41089 9999 41123
rect 9999 41089 10008 41123
rect 9956 41080 10008 41089
rect 10968 41123 11020 41132
rect 10968 41089 10977 41123
rect 10977 41089 11011 41123
rect 11011 41089 11020 41123
rect 10968 41080 11020 41089
rect 1308 41012 1360 41064
rect 9496 41012 9548 41064
rect 11520 41012 11572 41064
rect 11796 41012 11848 41064
rect 6828 40944 6880 40996
rect 7196 40944 7248 40996
rect 8852 40944 8904 40996
rect 9404 40944 9456 40996
rect 10968 40944 11020 40996
rect 6920 40876 6972 40928
rect 7840 40876 7892 40928
rect 8576 40876 8628 40928
rect 9496 40876 9548 40928
rect 10876 40876 10928 40928
rect 2582 40774 2634 40826
rect 2646 40774 2698 40826
rect 2710 40774 2762 40826
rect 2774 40774 2826 40826
rect 2838 40774 2890 40826
rect 5845 40774 5897 40826
rect 5909 40774 5961 40826
rect 5973 40774 6025 40826
rect 6037 40774 6089 40826
rect 6101 40774 6153 40826
rect 9109 40774 9161 40826
rect 9173 40774 9225 40826
rect 9237 40774 9289 40826
rect 9301 40774 9353 40826
rect 9365 40774 9417 40826
rect 4988 40672 5040 40724
rect 5448 40672 5500 40724
rect 7196 40672 7248 40724
rect 7932 40672 7984 40724
rect 10876 40672 10928 40724
rect 2044 40647 2096 40656
rect 2044 40613 2053 40647
rect 2053 40613 2087 40647
rect 2087 40613 2096 40647
rect 2044 40604 2096 40613
rect 9128 40604 9180 40656
rect 11612 40604 11664 40656
rect 10140 40536 10192 40588
rect 5632 40468 5684 40520
rect 9864 40511 9916 40520
rect 9864 40477 9873 40511
rect 9873 40477 9907 40511
rect 9907 40477 9916 40511
rect 9864 40468 9916 40477
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 7472 40400 7524 40452
rect 7932 40400 7984 40452
rect 8208 40400 8260 40452
rect 5632 40332 5684 40384
rect 8024 40332 8076 40384
rect 10784 40400 10836 40452
rect 9312 40375 9364 40384
rect 9312 40341 9321 40375
rect 9321 40341 9355 40375
rect 9355 40341 9364 40375
rect 9312 40332 9364 40341
rect 10048 40375 10100 40384
rect 10048 40341 10057 40375
rect 10057 40341 10091 40375
rect 10091 40341 10100 40375
rect 10048 40332 10100 40341
rect 10416 40332 10468 40384
rect 11796 40332 11848 40384
rect 4213 40230 4265 40282
rect 4277 40230 4329 40282
rect 4341 40230 4393 40282
rect 4405 40230 4457 40282
rect 4469 40230 4521 40282
rect 7477 40230 7529 40282
rect 7541 40230 7593 40282
rect 7605 40230 7657 40282
rect 7669 40230 7721 40282
rect 7733 40230 7785 40282
rect 1584 40060 1636 40112
rect 3884 40060 3936 40112
rect 1676 40035 1728 40044
rect 1676 40001 1685 40035
rect 1685 40001 1719 40035
rect 1719 40001 1728 40035
rect 1676 39992 1728 40001
rect 2044 39992 2096 40044
rect 3332 39992 3384 40044
rect 1400 39967 1452 39976
rect 1400 39933 1409 39967
rect 1409 39933 1443 39967
rect 1443 39933 1452 39967
rect 1400 39924 1452 39933
rect 6460 40060 6512 40112
rect 8576 40060 8628 40112
rect 9864 40060 9916 40112
rect 10784 40060 10836 40112
rect 10140 39992 10192 40044
rect 6552 39924 6604 39976
rect 7472 39856 7524 39908
rect 9128 39856 9180 39908
rect 10416 39924 10468 39976
rect 6552 39788 6604 39840
rect 8668 39831 8720 39840
rect 8668 39797 8677 39831
rect 8677 39797 8711 39831
rect 8711 39797 8720 39831
rect 8668 39788 8720 39797
rect 10692 39788 10744 39840
rect 2582 39686 2634 39738
rect 2646 39686 2698 39738
rect 2710 39686 2762 39738
rect 2774 39686 2826 39738
rect 2838 39686 2890 39738
rect 5845 39686 5897 39738
rect 5909 39686 5961 39738
rect 5973 39686 6025 39738
rect 6037 39686 6089 39738
rect 6101 39686 6153 39738
rect 9109 39686 9161 39738
rect 9173 39686 9225 39738
rect 9237 39686 9289 39738
rect 9301 39686 9353 39738
rect 9365 39686 9417 39738
rect 2504 39584 2556 39636
rect 1676 39516 1728 39568
rect 7012 39584 7064 39636
rect 9956 39584 10008 39636
rect 11888 39516 11940 39568
rect 2320 39491 2372 39500
rect 2320 39457 2329 39491
rect 2329 39457 2363 39491
rect 2363 39457 2372 39491
rect 2320 39448 2372 39457
rect 3240 39448 3292 39500
rect 6552 39448 6604 39500
rect 9496 39448 9548 39500
rect 9956 39448 10008 39500
rect 5172 39423 5224 39432
rect 5172 39389 5181 39423
rect 5181 39389 5215 39423
rect 5215 39389 5224 39423
rect 5172 39380 5224 39389
rect 2504 39312 2556 39364
rect 10140 39380 10192 39432
rect 2228 39244 2280 39296
rect 9404 39312 9456 39364
rect 4988 39244 5040 39296
rect 5172 39244 5224 39296
rect 5632 39244 5684 39296
rect 6552 39244 6604 39296
rect 10416 39312 10468 39364
rect 9864 39244 9916 39296
rect 4213 39142 4265 39194
rect 4277 39142 4329 39194
rect 4341 39142 4393 39194
rect 4405 39142 4457 39194
rect 4469 39142 4521 39194
rect 7477 39142 7529 39194
rect 7541 39142 7593 39194
rect 7605 39142 7657 39194
rect 7669 39142 7721 39194
rect 7733 39142 7785 39194
rect 1584 39083 1636 39092
rect 1584 39049 1593 39083
rect 1593 39049 1627 39083
rect 1627 39049 1636 39083
rect 1584 39040 1636 39049
rect 6828 38972 6880 39024
rect 8024 38972 8076 39024
rect 8668 38972 8720 39024
rect 1400 38947 1452 38956
rect 1400 38913 1409 38947
rect 1409 38913 1443 38947
rect 1443 38913 1452 38947
rect 1400 38904 1452 38913
rect 3700 38904 3752 38956
rect 10416 38972 10468 39024
rect 9496 38879 9548 38888
rect 1952 38768 2004 38820
rect 9496 38845 9505 38879
rect 9505 38845 9539 38879
rect 9539 38845 9548 38879
rect 9496 38836 9548 38845
rect 10048 38836 10100 38888
rect 9128 38811 9180 38820
rect 9128 38777 9137 38811
rect 9137 38777 9171 38811
rect 9171 38777 9180 38811
rect 9128 38768 9180 38777
rect 8116 38700 8168 38752
rect 2582 38598 2634 38650
rect 2646 38598 2698 38650
rect 2710 38598 2762 38650
rect 2774 38598 2826 38650
rect 2838 38598 2890 38650
rect 5845 38598 5897 38650
rect 5909 38598 5961 38650
rect 5973 38598 6025 38650
rect 6037 38598 6089 38650
rect 6101 38598 6153 38650
rect 9109 38598 9161 38650
rect 9173 38598 9225 38650
rect 9237 38598 9289 38650
rect 9301 38598 9353 38650
rect 9365 38598 9417 38650
rect 572 38496 624 38548
rect 7104 38496 7156 38548
rect 9588 38496 9640 38548
rect 9312 38428 9364 38480
rect 6368 38360 6420 38412
rect 7748 38360 7800 38412
rect 9588 38403 9640 38412
rect 9588 38369 9597 38403
rect 9597 38369 9631 38403
rect 9631 38369 9640 38403
rect 9588 38360 9640 38369
rect 10048 38360 10100 38412
rect 1400 38335 1452 38344
rect 1400 38301 1409 38335
rect 1409 38301 1443 38335
rect 1443 38301 1452 38335
rect 1400 38292 1452 38301
rect 4804 38292 4856 38344
rect 8116 38156 8168 38208
rect 9220 38156 9272 38208
rect 4213 38054 4265 38106
rect 4277 38054 4329 38106
rect 4341 38054 4393 38106
rect 4405 38054 4457 38106
rect 4469 38054 4521 38106
rect 7477 38054 7529 38106
rect 7541 38054 7593 38106
rect 7605 38054 7657 38106
rect 7669 38054 7721 38106
rect 7733 38054 7785 38106
rect 9496 37995 9548 38004
rect 9496 37961 9505 37995
rect 9505 37961 9539 37995
rect 9539 37961 9548 37995
rect 9496 37952 9548 37961
rect 9956 37884 10008 37936
rect 1308 37816 1360 37868
rect 4896 37816 4948 37868
rect 8668 37816 8720 37868
rect 8024 37748 8076 37800
rect 9588 37791 9640 37800
rect 9588 37757 9597 37791
rect 9597 37757 9631 37791
rect 9631 37757 9640 37791
rect 9588 37748 9640 37757
rect 2688 37680 2740 37732
rect 7748 37680 7800 37732
rect 9128 37680 9180 37732
rect 9588 37612 9640 37664
rect 2582 37510 2634 37562
rect 2646 37510 2698 37562
rect 2710 37510 2762 37562
rect 2774 37510 2826 37562
rect 2838 37510 2890 37562
rect 5845 37510 5897 37562
rect 5909 37510 5961 37562
rect 5973 37510 6025 37562
rect 6037 37510 6089 37562
rect 6101 37510 6153 37562
rect 9109 37510 9161 37562
rect 9173 37510 9225 37562
rect 9237 37510 9289 37562
rect 9301 37510 9353 37562
rect 9365 37510 9417 37562
rect 7748 37408 7800 37460
rect 8116 37340 8168 37392
rect 2504 37272 2556 37324
rect 8392 37408 8444 37460
rect 8576 37408 8628 37460
rect 2228 37204 2280 37256
rect 6920 37204 6972 37256
rect 8116 37247 8168 37256
rect 8116 37213 8125 37247
rect 8125 37213 8159 37247
rect 8159 37213 8168 37247
rect 8116 37204 8168 37213
rect 8300 37204 8352 37256
rect 8484 37204 8536 37256
rect 9680 37315 9732 37324
rect 9680 37281 9689 37315
rect 9689 37281 9723 37315
rect 9723 37281 9732 37315
rect 9680 37272 9732 37281
rect 5632 37136 5684 37188
rect 1768 37111 1820 37120
rect 1768 37077 1777 37111
rect 1777 37077 1811 37111
rect 1811 37077 1820 37111
rect 1768 37068 1820 37077
rect 2320 37068 2372 37120
rect 8116 37068 8168 37120
rect 8484 37068 8536 37120
rect 9864 37068 9916 37120
rect 11336 37068 11388 37120
rect 4213 36966 4265 37018
rect 4277 36966 4329 37018
rect 4341 36966 4393 37018
rect 4405 36966 4457 37018
rect 4469 36966 4521 37018
rect 7477 36966 7529 37018
rect 7541 36966 7593 37018
rect 7605 36966 7657 37018
rect 7669 36966 7721 37018
rect 7733 36966 7785 37018
rect 1768 36864 1820 36916
rect 6276 36864 6328 36916
rect 8852 36864 8904 36916
rect 3424 36796 3476 36848
rect 1584 36728 1636 36780
rect 9588 36796 9640 36848
rect 9680 36796 9732 36848
rect 1400 36703 1452 36712
rect 1400 36669 1409 36703
rect 1409 36669 1443 36703
rect 1443 36669 1452 36703
rect 1400 36660 1452 36669
rect 6920 36660 6972 36712
rect 11336 36932 11388 36984
rect 11612 36932 11664 36984
rect 11612 36796 11664 36848
rect 8116 36635 8168 36644
rect 8116 36601 8125 36635
rect 8125 36601 8159 36635
rect 8159 36601 8168 36635
rect 8116 36592 8168 36601
rect 8852 36567 8904 36576
rect 8852 36533 8861 36567
rect 8861 36533 8895 36567
rect 8895 36533 8904 36567
rect 8852 36524 8904 36533
rect 9496 36567 9548 36576
rect 9496 36533 9505 36567
rect 9505 36533 9539 36567
rect 9539 36533 9548 36567
rect 9496 36524 9548 36533
rect 11612 36524 11664 36576
rect 2582 36422 2634 36474
rect 2646 36422 2698 36474
rect 2710 36422 2762 36474
rect 2774 36422 2826 36474
rect 2838 36422 2890 36474
rect 5845 36422 5897 36474
rect 5909 36422 5961 36474
rect 5973 36422 6025 36474
rect 6037 36422 6089 36474
rect 6101 36422 6153 36474
rect 9109 36422 9161 36474
rect 9173 36422 9225 36474
rect 9237 36422 9289 36474
rect 9301 36422 9353 36474
rect 9365 36422 9417 36474
rect 8024 36320 8076 36372
rect 5540 36252 5592 36304
rect 7840 36252 7892 36304
rect 10232 36252 10284 36304
rect 2320 36227 2372 36236
rect 2320 36193 2329 36227
rect 2329 36193 2363 36227
rect 2363 36193 2372 36227
rect 2320 36184 2372 36193
rect 2504 36184 2556 36236
rect 3056 36227 3108 36236
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 2412 36159 2464 36168
rect 2412 36125 2421 36159
rect 2421 36125 2455 36159
rect 2455 36125 2464 36159
rect 3056 36193 3065 36227
rect 3065 36193 3099 36227
rect 3099 36193 3108 36227
rect 3056 36184 3108 36193
rect 6276 36184 6328 36236
rect 8024 36184 8076 36236
rect 9404 36227 9456 36236
rect 9404 36193 9413 36227
rect 9413 36193 9447 36227
rect 9447 36193 9456 36227
rect 9404 36184 9456 36193
rect 9588 36227 9640 36236
rect 9588 36193 9597 36227
rect 9597 36193 9631 36227
rect 9631 36193 9640 36227
rect 9588 36184 9640 36193
rect 9680 36184 9732 36236
rect 2412 36116 2464 36125
rect 1400 35980 1452 36032
rect 8852 35980 8904 36032
rect 4213 35878 4265 35930
rect 4277 35878 4329 35930
rect 4341 35878 4393 35930
rect 4405 35878 4457 35930
rect 4469 35878 4521 35930
rect 7477 35878 7529 35930
rect 7541 35878 7593 35930
rect 7605 35878 7657 35930
rect 7669 35878 7721 35930
rect 7733 35878 7785 35930
rect 5632 35776 5684 35828
rect 9864 35776 9916 35828
rect 10140 35776 10192 35828
rect 6368 35708 6420 35760
rect 1584 35683 1636 35692
rect 1584 35649 1593 35683
rect 1593 35649 1627 35683
rect 1627 35649 1636 35683
rect 1584 35640 1636 35649
rect 7196 35640 7248 35692
rect 7196 35504 7248 35556
rect 8116 35436 8168 35488
rect 10140 35436 10192 35488
rect 2582 35334 2634 35386
rect 2646 35334 2698 35386
rect 2710 35334 2762 35386
rect 2774 35334 2826 35386
rect 2838 35334 2890 35386
rect 5845 35334 5897 35386
rect 5909 35334 5961 35386
rect 5973 35334 6025 35386
rect 6037 35334 6089 35386
rect 6101 35334 6153 35386
rect 9109 35334 9161 35386
rect 9173 35334 9225 35386
rect 9237 35334 9289 35386
rect 9301 35334 9353 35386
rect 9365 35334 9417 35386
rect 1400 35275 1452 35284
rect 1400 35241 1409 35275
rect 1409 35241 1443 35275
rect 1443 35241 1452 35275
rect 1400 35232 1452 35241
rect 8852 35232 8904 35284
rect 2320 35096 2372 35148
rect 2596 35139 2648 35148
rect 2596 35105 2605 35139
rect 2605 35105 2639 35139
rect 2639 35105 2648 35139
rect 2596 35096 2648 35105
rect 9312 35096 9364 35148
rect 10048 35096 10100 35148
rect 1584 35071 1636 35080
rect 1584 35037 1593 35071
rect 1593 35037 1627 35071
rect 1627 35037 1636 35071
rect 1584 35028 1636 35037
rect 2044 35028 2096 35080
rect 2412 35071 2464 35080
rect 2412 35037 2421 35071
rect 2421 35037 2455 35071
rect 2455 35037 2464 35071
rect 2412 35028 2464 35037
rect 4620 35028 4672 35080
rect 9772 35028 9824 35080
rect 8116 34960 8168 35012
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 4213 34790 4265 34842
rect 4277 34790 4329 34842
rect 4341 34790 4393 34842
rect 4405 34790 4457 34842
rect 4469 34790 4521 34842
rect 7477 34790 7529 34842
rect 7541 34790 7593 34842
rect 7605 34790 7657 34842
rect 7669 34790 7721 34842
rect 7733 34790 7785 34842
rect 4804 34688 4856 34740
rect 3148 34663 3200 34672
rect 3148 34629 3157 34663
rect 3157 34629 3191 34663
rect 3191 34629 3200 34663
rect 3148 34620 3200 34629
rect 9312 34620 9364 34672
rect 2504 34595 2556 34604
rect 2504 34561 2513 34595
rect 2513 34561 2547 34595
rect 2547 34561 2556 34595
rect 2504 34552 2556 34561
rect 2596 34552 2648 34604
rect 8668 34552 8720 34604
rect 8852 34552 8904 34604
rect 664 34484 716 34536
rect 2320 34484 2372 34536
rect 7840 34484 7892 34536
rect 9588 34416 9640 34468
rect 10140 34484 10192 34536
rect 2582 34246 2634 34298
rect 2646 34246 2698 34298
rect 2710 34246 2762 34298
rect 2774 34246 2826 34298
rect 2838 34246 2890 34298
rect 5845 34246 5897 34298
rect 5909 34246 5961 34298
rect 5973 34246 6025 34298
rect 6037 34246 6089 34298
rect 6101 34246 6153 34298
rect 9109 34246 9161 34298
rect 9173 34246 9225 34298
rect 9237 34246 9289 34298
rect 9301 34246 9353 34298
rect 9365 34246 9417 34298
rect 8024 34144 8076 34196
rect 9772 34144 9824 34196
rect 6460 34008 6512 34060
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 7104 33940 7156 33992
rect 10876 33940 10928 33992
rect 9312 33847 9364 33856
rect 9312 33813 9321 33847
rect 9321 33813 9355 33847
rect 9355 33813 9364 33847
rect 9312 33804 9364 33813
rect 10048 33847 10100 33856
rect 10048 33813 10057 33847
rect 10057 33813 10091 33847
rect 10091 33813 10100 33847
rect 10048 33804 10100 33813
rect 4213 33702 4265 33754
rect 4277 33702 4329 33754
rect 4341 33702 4393 33754
rect 4405 33702 4457 33754
rect 4469 33702 4521 33754
rect 7477 33702 7529 33754
rect 7541 33702 7593 33754
rect 7605 33702 7657 33754
rect 7669 33702 7721 33754
rect 7733 33702 7785 33754
rect 3424 33600 3476 33652
rect 10784 33600 10836 33652
rect 4988 33464 5040 33516
rect 8668 33507 8720 33516
rect 8668 33473 8677 33507
rect 8677 33473 8711 33507
rect 8711 33473 8720 33507
rect 8668 33464 8720 33473
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 10140 33396 10192 33448
rect 9588 33328 9640 33380
rect 8024 33260 8076 33312
rect 10692 33260 10744 33312
rect 2582 33158 2634 33210
rect 2646 33158 2698 33210
rect 2710 33158 2762 33210
rect 2774 33158 2826 33210
rect 2838 33158 2890 33210
rect 5845 33158 5897 33210
rect 5909 33158 5961 33210
rect 5973 33158 6025 33210
rect 6037 33158 6089 33210
rect 6101 33158 6153 33210
rect 9109 33158 9161 33210
rect 9173 33158 9225 33210
rect 9237 33158 9289 33210
rect 9301 33158 9353 33210
rect 9365 33158 9417 33210
rect 2228 33056 2280 33108
rect 8116 33056 8168 33108
rect 8484 33056 8536 33108
rect 10600 33056 10652 33108
rect 4896 32988 4948 33040
rect 9680 32988 9732 33040
rect 9864 32988 9916 33040
rect 2504 32920 2556 32972
rect 8116 32920 8168 32972
rect 8852 32920 8904 32972
rect 1584 32895 1636 32904
rect 1584 32861 1593 32895
rect 1593 32861 1627 32895
rect 1627 32861 1636 32895
rect 1584 32852 1636 32861
rect 2320 32852 2372 32904
rect 7012 32852 7064 32904
rect 11336 32988 11388 33040
rect 7104 32784 7156 32836
rect 9496 32784 9548 32836
rect 10140 32920 10192 32972
rect 10600 32920 10652 32972
rect 11520 32920 11572 32972
rect 2136 32759 2188 32768
rect 2136 32725 2145 32759
rect 2145 32725 2179 32759
rect 2179 32725 2188 32759
rect 2136 32716 2188 32725
rect 2504 32759 2556 32768
rect 2504 32725 2513 32759
rect 2513 32725 2547 32759
rect 2547 32725 2556 32759
rect 2504 32716 2556 32725
rect 9220 32759 9272 32768
rect 9220 32725 9229 32759
rect 9229 32725 9263 32759
rect 9263 32725 9272 32759
rect 9220 32716 9272 32725
rect 9404 32716 9456 32768
rect 11704 32716 11756 32768
rect 4213 32614 4265 32666
rect 4277 32614 4329 32666
rect 4341 32614 4393 32666
rect 4405 32614 4457 32666
rect 4469 32614 4521 32666
rect 7477 32614 7529 32666
rect 7541 32614 7593 32666
rect 7605 32614 7657 32666
rect 7669 32614 7721 32666
rect 7733 32614 7785 32666
rect 11336 32648 11388 32700
rect 11888 32691 11940 32700
rect 11888 32657 11897 32691
rect 11897 32657 11931 32691
rect 11931 32657 11940 32691
rect 11888 32648 11940 32657
rect 2044 32512 2096 32564
rect 2136 32512 2188 32564
rect 10048 32512 10100 32564
rect 10140 32444 10192 32496
rect 11060 32444 11112 32496
rect 1584 32419 1636 32428
rect 1584 32385 1593 32419
rect 1593 32385 1627 32419
rect 1627 32385 1636 32419
rect 1584 32376 1636 32385
rect 5448 32376 5500 32428
rect 11428 32376 11480 32428
rect 9404 32308 9456 32360
rect 5172 32240 5224 32292
rect 5448 32240 5500 32292
rect 11152 32240 11204 32292
rect 8852 32215 8904 32224
rect 8852 32181 8861 32215
rect 8861 32181 8895 32215
rect 8895 32181 8904 32215
rect 8852 32172 8904 32181
rect 2582 32070 2634 32122
rect 2646 32070 2698 32122
rect 2710 32070 2762 32122
rect 2774 32070 2826 32122
rect 2838 32070 2890 32122
rect 5845 32070 5897 32122
rect 5909 32070 5961 32122
rect 5973 32070 6025 32122
rect 6037 32070 6089 32122
rect 6101 32070 6153 32122
rect 9109 32070 9161 32122
rect 9173 32070 9225 32122
rect 9237 32070 9289 32122
rect 9301 32070 9353 32122
rect 9365 32070 9417 32122
rect 2504 31968 2556 32020
rect 10784 31968 10836 32020
rect 11796 32036 11848 32088
rect 11244 31968 11296 32020
rect 11336 31968 11388 32020
rect 6184 31832 6236 31884
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 10600 31764 10652 31816
rect 10876 31764 10928 31816
rect 9956 31696 10008 31748
rect 10140 31696 10192 31748
rect 11612 31900 11664 31952
rect 11336 31764 11388 31816
rect 11888 31764 11940 31816
rect 4213 31526 4265 31578
rect 4277 31526 4329 31578
rect 4341 31526 4393 31578
rect 4405 31526 4457 31578
rect 4469 31526 4521 31578
rect 7477 31526 7529 31578
rect 7541 31526 7593 31578
rect 7605 31526 7657 31578
rect 7669 31526 7721 31578
rect 7733 31526 7785 31578
rect 9956 31424 10008 31476
rect 10692 31424 10744 31476
rect 10048 31263 10100 31272
rect 10048 31229 10057 31263
rect 10057 31229 10091 31263
rect 10091 31229 10100 31263
rect 10048 31220 10100 31229
rect 10140 31220 10192 31272
rect 10416 31220 10468 31272
rect 10968 31220 11020 31272
rect 11428 31560 11480 31612
rect 11520 31492 11572 31544
rect 11704 31560 11756 31612
rect 11612 31220 11664 31272
rect 10692 31152 10744 31204
rect 8852 31084 8904 31136
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 2582 30982 2634 31034
rect 2646 30982 2698 31034
rect 2710 30982 2762 31034
rect 2774 30982 2826 31034
rect 2838 30982 2890 31034
rect 5845 30982 5897 31034
rect 5909 30982 5961 31034
rect 5973 30982 6025 31034
rect 6037 30982 6089 31034
rect 6101 30982 6153 31034
rect 9109 30982 9161 31034
rect 9173 30982 9225 31034
rect 9237 30982 9289 31034
rect 9301 30982 9353 31034
rect 9365 30982 9417 31034
rect 10140 30744 10192 30796
rect 7380 30676 7432 30728
rect 10048 30676 10100 30728
rect 10416 30744 10468 30796
rect 10416 30608 10468 30660
rect 1584 30583 1636 30592
rect 1584 30549 1593 30583
rect 1593 30549 1627 30583
rect 1627 30549 1636 30583
rect 1584 30540 1636 30549
rect 10048 30583 10100 30592
rect 10048 30549 10057 30583
rect 10057 30549 10091 30583
rect 10091 30549 10100 30583
rect 10048 30540 10100 30549
rect 4213 30438 4265 30490
rect 4277 30438 4329 30490
rect 4341 30438 4393 30490
rect 4405 30438 4457 30490
rect 4469 30438 4521 30490
rect 7477 30438 7529 30490
rect 7541 30438 7593 30490
rect 7605 30438 7657 30490
rect 7669 30438 7721 30490
rect 7733 30438 7785 30490
rect 10140 30268 10192 30320
rect 10600 30200 10652 30252
rect 1584 30039 1636 30048
rect 1584 30005 1593 30039
rect 1593 30005 1627 30039
rect 1627 30005 1636 30039
rect 1584 29996 1636 30005
rect 10048 30039 10100 30048
rect 10048 30005 10057 30039
rect 10057 30005 10091 30039
rect 10091 30005 10100 30039
rect 10048 29996 10100 30005
rect 2582 29894 2634 29946
rect 2646 29894 2698 29946
rect 2710 29894 2762 29946
rect 2774 29894 2826 29946
rect 2838 29894 2890 29946
rect 5845 29894 5897 29946
rect 5909 29894 5961 29946
rect 5973 29894 6025 29946
rect 6037 29894 6089 29946
rect 6101 29894 6153 29946
rect 9109 29894 9161 29946
rect 9173 29894 9225 29946
rect 9237 29894 9289 29946
rect 9301 29894 9353 29946
rect 9365 29894 9417 29946
rect 10048 29656 10100 29708
rect 11888 29699 11940 29708
rect 11888 29665 11897 29699
rect 11897 29665 11931 29699
rect 11931 29665 11940 29699
rect 11888 29656 11940 29665
rect 9864 29631 9916 29640
rect 9864 29597 9873 29631
rect 9873 29597 9907 29631
rect 9907 29597 9916 29631
rect 9864 29588 9916 29597
rect 10140 29520 10192 29572
rect 1584 29495 1636 29504
rect 1584 29461 1593 29495
rect 1593 29461 1627 29495
rect 1627 29461 1636 29495
rect 1584 29452 1636 29461
rect 9312 29495 9364 29504
rect 9312 29461 9321 29495
rect 9321 29461 9355 29495
rect 9355 29461 9364 29495
rect 9312 29452 9364 29461
rect 10048 29495 10100 29504
rect 10048 29461 10057 29495
rect 10057 29461 10091 29495
rect 10091 29461 10100 29495
rect 10048 29452 10100 29461
rect 4213 29350 4265 29402
rect 4277 29350 4329 29402
rect 4341 29350 4393 29402
rect 4405 29350 4457 29402
rect 4469 29350 4521 29402
rect 7477 29350 7529 29402
rect 7541 29350 7593 29402
rect 7605 29350 7657 29402
rect 7669 29350 7721 29402
rect 7733 29350 7785 29402
rect 7380 29248 7432 29300
rect 9864 29291 9916 29300
rect 9864 29257 9873 29291
rect 9873 29257 9907 29291
rect 9907 29257 9916 29291
rect 9864 29248 9916 29257
rect 1952 29112 2004 29164
rect 7288 29112 7340 29164
rect 9864 29044 9916 29096
rect 10416 29044 10468 29096
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 7288 28976 7340 29028
rect 9128 28976 9180 29028
rect 2582 28806 2634 28858
rect 2646 28806 2698 28858
rect 2710 28806 2762 28858
rect 2774 28806 2826 28858
rect 2838 28806 2890 28858
rect 5845 28806 5897 28858
rect 5909 28806 5961 28858
rect 5973 28806 6025 28858
rect 6037 28806 6089 28858
rect 6101 28806 6153 28858
rect 9109 28806 9161 28858
rect 9173 28806 9225 28858
rect 9237 28806 9289 28858
rect 9301 28806 9353 28858
rect 9365 28806 9417 28858
rect 7196 28500 7248 28552
rect 8668 28500 8720 28552
rect 10232 28500 10284 28552
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 9312 28407 9364 28416
rect 9312 28373 9321 28407
rect 9321 28373 9355 28407
rect 9355 28373 9364 28407
rect 9312 28364 9364 28373
rect 10140 28364 10192 28416
rect 4213 28262 4265 28314
rect 4277 28262 4329 28314
rect 4341 28262 4393 28314
rect 4405 28262 4457 28314
rect 4469 28262 4521 28314
rect 7477 28262 7529 28314
rect 7541 28262 7593 28314
rect 7605 28262 7657 28314
rect 7669 28262 7721 28314
rect 7733 28262 7785 28314
rect 10232 28160 10284 28212
rect 11244 28160 11296 28212
rect 11888 28160 11940 28212
rect 10048 27863 10100 27872
rect 10048 27829 10057 27863
rect 10057 27829 10091 27863
rect 10091 27829 10100 27863
rect 10048 27820 10100 27829
rect 2582 27718 2634 27770
rect 2646 27718 2698 27770
rect 2710 27718 2762 27770
rect 2774 27718 2826 27770
rect 2838 27718 2890 27770
rect 5845 27718 5897 27770
rect 5909 27718 5961 27770
rect 5973 27718 6025 27770
rect 6037 27718 6089 27770
rect 6101 27718 6153 27770
rect 9109 27718 9161 27770
rect 9173 27718 9225 27770
rect 9237 27718 9289 27770
rect 9301 27718 9353 27770
rect 9365 27718 9417 27770
rect 7012 27412 7064 27464
rect 9680 27412 9732 27464
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 10140 27276 10192 27328
rect 4213 27174 4265 27226
rect 4277 27174 4329 27226
rect 4341 27174 4393 27226
rect 4405 27174 4457 27226
rect 4469 27174 4521 27226
rect 7477 27174 7529 27226
rect 7541 27174 7593 27226
rect 7605 27174 7657 27226
rect 7669 27174 7721 27226
rect 7733 27174 7785 27226
rect 8116 27004 8168 27056
rect 8852 27004 8904 27056
rect 7196 26936 7248 26988
rect 7932 26936 7984 26988
rect 8668 26936 8720 26988
rect 8944 26936 8996 26988
rect 9772 26936 9824 26988
rect 1584 26775 1636 26784
rect 1584 26741 1593 26775
rect 1593 26741 1627 26775
rect 1627 26741 1636 26775
rect 1584 26732 1636 26741
rect 9036 26732 9088 26784
rect 10048 26775 10100 26784
rect 10048 26741 10057 26775
rect 10057 26741 10091 26775
rect 10091 26741 10100 26775
rect 10048 26732 10100 26741
rect 2582 26630 2634 26682
rect 2646 26630 2698 26682
rect 2710 26630 2762 26682
rect 2774 26630 2826 26682
rect 2838 26630 2890 26682
rect 5845 26630 5897 26682
rect 5909 26630 5961 26682
rect 5973 26630 6025 26682
rect 6037 26630 6089 26682
rect 6101 26630 6153 26682
rect 9109 26630 9161 26682
rect 9173 26630 9225 26682
rect 9237 26630 9289 26682
rect 9301 26630 9353 26682
rect 9365 26630 9417 26682
rect 8944 26528 8996 26580
rect 9496 26528 9548 26580
rect 7932 26460 7984 26512
rect 8116 26460 8168 26512
rect 3608 26324 3660 26376
rect 9956 26324 10008 26376
rect 10600 26324 10652 26376
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 4213 26086 4265 26138
rect 4277 26086 4329 26138
rect 4341 26086 4393 26138
rect 4405 26086 4457 26138
rect 4469 26086 4521 26138
rect 7477 26086 7529 26138
rect 7541 26086 7593 26138
rect 7605 26086 7657 26138
rect 7669 26086 7721 26138
rect 7733 26086 7785 26138
rect 6736 25984 6788 26036
rect 11612 25916 11664 25968
rect 8484 25848 8536 25900
rect 9864 25891 9916 25900
rect 9864 25857 9873 25891
rect 9873 25857 9907 25891
rect 9907 25857 9916 25891
rect 9864 25848 9916 25857
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 9496 25644 9548 25696
rect 2582 25542 2634 25594
rect 2646 25542 2698 25594
rect 2710 25542 2762 25594
rect 2774 25542 2826 25594
rect 2838 25542 2890 25594
rect 5845 25542 5897 25594
rect 5909 25542 5961 25594
rect 5973 25542 6025 25594
rect 6037 25542 6089 25594
rect 6101 25542 6153 25594
rect 9109 25542 9161 25594
rect 9173 25542 9225 25594
rect 9237 25542 9289 25594
rect 9301 25542 9353 25594
rect 9365 25542 9417 25594
rect 10416 25372 10468 25424
rect 10968 25372 11020 25424
rect 9956 25347 10008 25356
rect 9956 25313 9965 25347
rect 9965 25313 9999 25347
rect 9999 25313 10008 25347
rect 9956 25304 10008 25313
rect 10968 25279 11020 25288
rect 10968 25245 10977 25279
rect 10977 25245 11011 25279
rect 11011 25245 11020 25279
rect 10968 25236 11020 25245
rect 1032 25168 1084 25220
rect 8484 25100 8536 25152
rect 9772 25143 9824 25152
rect 9772 25109 9781 25143
rect 9781 25109 9815 25143
rect 9815 25109 9824 25143
rect 9772 25100 9824 25109
rect 4213 24998 4265 25050
rect 4277 24998 4329 25050
rect 4341 24998 4393 25050
rect 4405 24998 4457 25050
rect 4469 24998 4521 25050
rect 7477 24998 7529 25050
rect 7541 24998 7593 25050
rect 7605 24998 7657 25050
rect 7669 24998 7721 25050
rect 7733 24998 7785 25050
rect 7104 24760 7156 24812
rect 9496 24760 9548 24812
rect 9956 24803 10008 24812
rect 9956 24769 9965 24803
rect 9965 24769 9999 24803
rect 9999 24769 10008 24803
rect 9956 24760 10008 24769
rect 10324 24760 10376 24812
rect 1584 24667 1636 24676
rect 1584 24633 1593 24667
rect 1593 24633 1627 24667
rect 1627 24633 1636 24667
rect 1584 24624 1636 24633
rect 11796 24624 11848 24676
rect 2582 24454 2634 24506
rect 2646 24454 2698 24506
rect 2710 24454 2762 24506
rect 2774 24454 2826 24506
rect 2838 24454 2890 24506
rect 5845 24454 5897 24506
rect 5909 24454 5961 24506
rect 5973 24454 6025 24506
rect 6037 24454 6089 24506
rect 6101 24454 6153 24506
rect 9109 24454 9161 24506
rect 9173 24454 9225 24506
rect 9237 24454 9289 24506
rect 9301 24454 9353 24506
rect 9365 24454 9417 24506
rect 4068 24352 4120 24404
rect 10508 24284 10560 24336
rect 4804 24148 4856 24200
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 10048 24148 10100 24200
rect 11796 24148 11848 24200
rect 9496 24080 9548 24132
rect 11704 24080 11756 24132
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 4213 23910 4265 23962
rect 4277 23910 4329 23962
rect 4341 23910 4393 23962
rect 4405 23910 4457 23962
rect 4469 23910 4521 23962
rect 7477 23910 7529 23962
rect 7541 23910 7593 23962
rect 7605 23910 7657 23962
rect 7669 23910 7721 23962
rect 7733 23910 7785 23962
rect 8760 23808 8812 23860
rect 11520 23808 11572 23860
rect 3424 23672 3476 23724
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 8760 23672 8812 23681
rect 9680 23672 9732 23724
rect 10140 23604 10192 23656
rect 6736 23536 6788 23588
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 2582 23366 2634 23418
rect 2646 23366 2698 23418
rect 2710 23366 2762 23418
rect 2774 23366 2826 23418
rect 2838 23366 2890 23418
rect 5845 23366 5897 23418
rect 5909 23366 5961 23418
rect 5973 23366 6025 23418
rect 6037 23366 6089 23418
rect 6101 23366 6153 23418
rect 9109 23366 9161 23418
rect 9173 23366 9225 23418
rect 9237 23366 9289 23418
rect 9301 23366 9353 23418
rect 9365 23366 9417 23418
rect 5448 23128 5500 23180
rect 10140 23128 10192 23180
rect 9036 23060 9088 23112
rect 10140 22992 10192 23044
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 5632 22924 5684 22976
rect 4213 22822 4265 22874
rect 4277 22822 4329 22874
rect 4341 22822 4393 22874
rect 4405 22822 4457 22874
rect 4469 22822 4521 22874
rect 7477 22822 7529 22874
rect 7541 22822 7593 22874
rect 7605 22822 7657 22874
rect 7669 22822 7721 22874
rect 7733 22822 7785 22874
rect 3792 22720 3844 22772
rect 11152 22720 11204 22772
rect 6552 22652 6604 22704
rect 10324 22652 10376 22704
rect 4896 22584 4948 22636
rect 7104 22584 7156 22636
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 8760 22516 8812 22568
rect 10232 22516 10284 22568
rect 6184 22448 6236 22500
rect 10784 22448 10836 22500
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 7840 22380 7892 22432
rect 2582 22278 2634 22330
rect 2646 22278 2698 22330
rect 2710 22278 2762 22330
rect 2774 22278 2826 22330
rect 2838 22278 2890 22330
rect 5845 22278 5897 22330
rect 5909 22278 5961 22330
rect 5973 22278 6025 22330
rect 6037 22278 6089 22330
rect 6101 22278 6153 22330
rect 9109 22278 9161 22330
rect 9173 22278 9225 22330
rect 9237 22278 9289 22330
rect 9301 22278 9353 22330
rect 9365 22278 9417 22330
rect 11244 22380 11296 22432
rect 11060 22244 11112 22296
rect 11336 22244 11388 22296
rect 11704 22244 11756 22296
rect 10968 22108 11020 22160
rect 8300 22040 8352 22092
rect 10324 22040 10376 22092
rect 11520 22083 11572 22092
rect 11520 22049 11529 22083
rect 11529 22049 11563 22083
rect 11563 22049 11572 22083
rect 11520 22040 11572 22049
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 10416 21972 10468 22024
rect 8116 21904 8168 21956
rect 11244 21904 11296 21956
rect 5264 21836 5316 21888
rect 9772 21836 9824 21888
rect 11796 21904 11848 21956
rect 11612 21836 11664 21888
rect 4213 21734 4265 21786
rect 4277 21734 4329 21786
rect 4341 21734 4393 21786
rect 4405 21734 4457 21786
rect 4469 21734 4521 21786
rect 7477 21734 7529 21786
rect 7541 21734 7593 21786
rect 7605 21734 7657 21786
rect 7669 21734 7721 21786
rect 7733 21734 7785 21786
rect 11060 21700 11112 21752
rect 11704 21700 11756 21752
rect 3516 21632 3568 21684
rect 10232 21564 10284 21616
rect 7380 21496 7432 21548
rect 10784 21496 10836 21548
rect 8760 21471 8812 21480
rect 8760 21437 8769 21471
rect 8769 21437 8803 21471
rect 8803 21437 8812 21471
rect 8760 21428 8812 21437
rect 9496 21428 9548 21480
rect 1584 21403 1636 21412
rect 1584 21369 1593 21403
rect 1593 21369 1627 21403
rect 1627 21369 1636 21403
rect 1584 21360 1636 21369
rect 9956 21360 10008 21412
rect 1400 21292 1452 21344
rect 1768 21292 1820 21344
rect 6920 21292 6972 21344
rect 8760 21292 8812 21344
rect 9588 21292 9640 21344
rect 2582 21190 2634 21242
rect 2646 21190 2698 21242
rect 2710 21190 2762 21242
rect 2774 21190 2826 21242
rect 2838 21190 2890 21242
rect 5845 21190 5897 21242
rect 5909 21190 5961 21242
rect 5973 21190 6025 21242
rect 6037 21190 6089 21242
rect 6101 21190 6153 21242
rect 9109 21190 9161 21242
rect 9173 21190 9225 21242
rect 9237 21190 9289 21242
rect 9301 21190 9353 21242
rect 9365 21190 9417 21242
rect 8484 20884 8536 20936
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 11152 20859 11204 20868
rect 11152 20825 11161 20859
rect 11161 20825 11195 20859
rect 11195 20825 11204 20859
rect 11152 20816 11204 20825
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 4213 20646 4265 20698
rect 4277 20646 4329 20698
rect 4341 20646 4393 20698
rect 4405 20646 4457 20698
rect 4469 20646 4521 20698
rect 7477 20646 7529 20698
rect 7541 20646 7593 20698
rect 7605 20646 7657 20698
rect 7669 20646 7721 20698
rect 7733 20646 7785 20698
rect 8024 20544 8076 20596
rect 10600 20544 10652 20596
rect 8668 20476 8720 20528
rect 9588 20476 9640 20528
rect 6736 20408 6788 20460
rect 8116 20408 8168 20460
rect 9496 20408 9548 20460
rect 8300 20272 8352 20324
rect 8944 20272 8996 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 2582 20102 2634 20154
rect 2646 20102 2698 20154
rect 2710 20102 2762 20154
rect 2774 20102 2826 20154
rect 2838 20102 2890 20154
rect 5845 20102 5897 20154
rect 5909 20102 5961 20154
rect 5973 20102 6025 20154
rect 6037 20102 6089 20154
rect 6101 20102 6153 20154
rect 9109 20102 9161 20154
rect 9173 20102 9225 20154
rect 9237 20102 9289 20154
rect 9301 20102 9353 20154
rect 9365 20102 9417 20154
rect 7932 20000 7984 20052
rect 8760 19932 8812 19984
rect 9312 19932 9364 19984
rect 9588 19864 9640 19916
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 10324 19864 10376 19916
rect 7840 19796 7892 19848
rect 8116 19796 8168 19848
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 7012 19660 7064 19712
rect 10048 19660 10100 19712
rect 4213 19558 4265 19610
rect 4277 19558 4329 19610
rect 4341 19558 4393 19610
rect 4405 19558 4457 19610
rect 4469 19558 4521 19610
rect 7477 19558 7529 19610
rect 7541 19558 7593 19610
rect 7605 19558 7657 19610
rect 7669 19558 7721 19610
rect 7733 19558 7785 19610
rect 8300 19456 8352 19508
rect 7932 19388 7984 19440
rect 6920 19320 6972 19372
rect 8300 19363 8352 19372
rect 8300 19329 8309 19363
rect 8309 19329 8343 19363
rect 8343 19329 8352 19363
rect 8300 19320 8352 19329
rect 9680 19388 9732 19440
rect 9036 19320 9088 19372
rect 9956 19431 10008 19440
rect 9956 19397 9965 19431
rect 9965 19397 9999 19431
rect 9999 19397 10008 19431
rect 9956 19388 10008 19397
rect 10324 19388 10376 19440
rect 9864 19320 9916 19372
rect 10508 19320 10560 19372
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2582 19014 2634 19066
rect 2646 19014 2698 19066
rect 2710 19014 2762 19066
rect 2774 19014 2826 19066
rect 2838 19014 2890 19066
rect 5845 19014 5897 19066
rect 5909 19014 5961 19066
rect 5973 19014 6025 19066
rect 6037 19014 6089 19066
rect 6101 19014 6153 19066
rect 9109 19014 9161 19066
rect 9173 19014 9225 19066
rect 9237 19014 9289 19066
rect 9301 19014 9353 19066
rect 9365 19014 9417 19066
rect 7288 18912 7340 18964
rect 9772 18912 9824 18964
rect 10232 18955 10284 18964
rect 10232 18921 10241 18955
rect 10241 18921 10275 18955
rect 10275 18921 10284 18955
rect 10232 18912 10284 18921
rect 10324 18776 10376 18828
rect 7840 18708 7892 18760
rect 8668 18708 8720 18760
rect 1400 18572 1452 18624
rect 9680 18572 9732 18624
rect 4213 18470 4265 18522
rect 4277 18470 4329 18522
rect 4341 18470 4393 18522
rect 4405 18470 4457 18522
rect 4469 18470 4521 18522
rect 7477 18470 7529 18522
rect 7541 18470 7593 18522
rect 7605 18470 7657 18522
rect 7669 18470 7721 18522
rect 7733 18470 7785 18522
rect 7104 18411 7156 18420
rect 7104 18377 7113 18411
rect 7113 18377 7147 18411
rect 7147 18377 7156 18411
rect 7104 18368 7156 18377
rect 8852 18368 8904 18420
rect 9588 18368 9640 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 8392 18275 8444 18284
rect 8392 18241 8401 18275
rect 8401 18241 8435 18275
rect 8435 18241 8444 18275
rect 8392 18232 8444 18241
rect 1584 18139 1636 18148
rect 1584 18105 1593 18139
rect 1593 18105 1627 18139
rect 1627 18105 1636 18139
rect 1584 18096 1636 18105
rect 7840 18028 7892 18080
rect 2582 17926 2634 17978
rect 2646 17926 2698 17978
rect 2710 17926 2762 17978
rect 2774 17926 2826 17978
rect 2838 17926 2890 17978
rect 5845 17926 5897 17978
rect 5909 17926 5961 17978
rect 5973 17926 6025 17978
rect 6037 17926 6089 17978
rect 6101 17926 6153 17978
rect 9109 17926 9161 17978
rect 9173 17926 9225 17978
rect 9237 17926 9289 17978
rect 9301 17926 9353 17978
rect 9365 17926 9417 17978
rect 9036 17824 9088 17876
rect 5356 17756 5408 17808
rect 5632 17688 5684 17740
rect 2964 17620 3016 17672
rect 7012 17620 7064 17672
rect 7380 17620 7432 17672
rect 9128 17552 9180 17604
rect 9864 17731 9916 17740
rect 9864 17697 9873 17731
rect 9873 17697 9907 17731
rect 9907 17697 9916 17731
rect 9864 17688 9916 17697
rect 10324 17688 10376 17740
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 6460 17484 6512 17536
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 8116 17527 8168 17536
rect 8116 17493 8125 17527
rect 8125 17493 8159 17527
rect 8159 17493 8168 17527
rect 8116 17484 8168 17493
rect 8760 17484 8812 17536
rect 9772 17527 9824 17536
rect 9772 17493 9781 17527
rect 9781 17493 9815 17527
rect 9815 17493 9824 17527
rect 9772 17484 9824 17493
rect 9864 17484 9916 17536
rect 4213 17382 4265 17434
rect 4277 17382 4329 17434
rect 4341 17382 4393 17434
rect 4405 17382 4457 17434
rect 4469 17382 4521 17434
rect 7477 17382 7529 17434
rect 7541 17382 7593 17434
rect 7605 17382 7657 17434
rect 7669 17382 7721 17434
rect 7733 17382 7785 17434
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 9588 17280 9640 17332
rect 3976 17212 4028 17264
rect 7656 17212 7708 17264
rect 7748 17212 7800 17264
rect 6184 17144 6236 17196
rect 6460 17187 6512 17196
rect 6460 17153 6469 17187
rect 6469 17153 6503 17187
rect 6503 17153 6512 17187
rect 6460 17144 6512 17153
rect 7196 17144 7248 17196
rect 8300 17144 8352 17196
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 10324 17076 10376 17128
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 6276 16940 6328 16992
rect 2582 16838 2634 16890
rect 2646 16838 2698 16890
rect 2710 16838 2762 16890
rect 2774 16838 2826 16890
rect 2838 16838 2890 16890
rect 5845 16838 5897 16890
rect 5909 16838 5961 16890
rect 5973 16838 6025 16890
rect 6037 16838 6089 16890
rect 6101 16838 6153 16890
rect 9109 16838 9161 16890
rect 9173 16838 9225 16890
rect 9237 16838 9289 16890
rect 9301 16838 9353 16890
rect 9365 16838 9417 16890
rect 7196 16736 7248 16788
rect 7656 16736 7708 16788
rect 9956 16736 10008 16788
rect 7012 16600 7064 16652
rect 7380 16600 7432 16652
rect 7932 16600 7984 16652
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 8484 16600 8536 16652
rect 10324 16600 10376 16652
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 7748 16464 7800 16516
rect 8116 16464 8168 16516
rect 6920 16396 6972 16448
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7196 16396 7248 16405
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 9220 16532 9272 16584
rect 11612 16532 11664 16584
rect 4213 16294 4265 16346
rect 4277 16294 4329 16346
rect 4341 16294 4393 16346
rect 4405 16294 4457 16346
rect 4469 16294 4521 16346
rect 7477 16294 7529 16346
rect 7541 16294 7593 16346
rect 7605 16294 7657 16346
rect 7669 16294 7721 16346
rect 7733 16294 7785 16346
rect 11060 16260 11112 16312
rect 7840 16167 7892 16176
rect 7840 16133 7874 16167
rect 7874 16133 7892 16167
rect 7840 16124 7892 16133
rect 10232 16192 10284 16244
rect 9680 16124 9732 16176
rect 11888 16124 11940 16176
rect 6920 16056 6972 16108
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 7196 16056 7248 16108
rect 6736 15988 6788 16040
rect 9588 15988 9640 16040
rect 10324 15988 10376 16040
rect 10048 15920 10100 15972
rect 480 15852 532 15904
rect 5356 15852 5408 15904
rect 7288 15852 7340 15904
rect 7932 15852 7984 15904
rect 2582 15750 2634 15802
rect 2646 15750 2698 15802
rect 2710 15750 2762 15802
rect 2774 15750 2826 15802
rect 2838 15750 2890 15802
rect 5845 15750 5897 15802
rect 5909 15750 5961 15802
rect 5973 15750 6025 15802
rect 6037 15750 6089 15802
rect 6101 15750 6153 15802
rect 9109 15750 9161 15802
rect 9173 15750 9225 15802
rect 9237 15750 9289 15802
rect 9301 15750 9353 15802
rect 9365 15750 9417 15802
rect 5356 15648 5408 15700
rect 8300 15580 8352 15632
rect 7196 15512 7248 15564
rect 7288 15512 7340 15564
rect 10140 15580 10192 15632
rect 6828 15444 6880 15496
rect 8116 15444 8168 15496
rect 8300 15444 8352 15496
rect 9404 15444 9456 15496
rect 9772 15444 9824 15496
rect 10324 15512 10376 15564
rect 6644 15376 6696 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 6736 15308 6788 15360
rect 8668 15308 8720 15360
rect 8944 15308 8996 15360
rect 9404 15351 9456 15360
rect 9404 15317 9413 15351
rect 9413 15317 9447 15351
rect 9447 15317 9456 15351
rect 9404 15308 9456 15317
rect 9772 15351 9824 15360
rect 9772 15317 9781 15351
rect 9781 15317 9815 15351
rect 9815 15317 9824 15351
rect 9772 15308 9824 15317
rect 4213 15206 4265 15258
rect 4277 15206 4329 15258
rect 4341 15206 4393 15258
rect 4405 15206 4457 15258
rect 4469 15206 4521 15258
rect 7477 15206 7529 15258
rect 7541 15206 7593 15258
rect 7605 15206 7657 15258
rect 7669 15206 7721 15258
rect 7733 15206 7785 15258
rect 7932 15104 7984 15156
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 8668 15104 8720 15113
rect 8852 15104 8904 15156
rect 9772 15104 9824 15156
rect 8300 15036 8352 15088
rect 11520 15104 11572 15156
rect 7472 14968 7524 15020
rect 8484 14968 8536 15020
rect 5632 14900 5684 14952
rect 7840 14832 7892 14884
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 7104 14764 7156 14816
rect 7380 14764 7432 14816
rect 7656 14764 7708 14816
rect 8392 14900 8444 14952
rect 9036 14968 9088 15020
rect 10324 14900 10376 14952
rect 8944 14764 8996 14816
rect 2582 14662 2634 14714
rect 2646 14662 2698 14714
rect 2710 14662 2762 14714
rect 2774 14662 2826 14714
rect 2838 14662 2890 14714
rect 5845 14662 5897 14714
rect 5909 14662 5961 14714
rect 5973 14662 6025 14714
rect 6037 14662 6089 14714
rect 6101 14662 6153 14714
rect 9109 14662 9161 14714
rect 9173 14662 9225 14714
rect 9237 14662 9289 14714
rect 9301 14662 9353 14714
rect 9365 14662 9417 14714
rect 8944 14560 8996 14612
rect 5264 14535 5316 14544
rect 5264 14501 5273 14535
rect 5273 14501 5307 14535
rect 5307 14501 5316 14535
rect 5264 14492 5316 14501
rect 6920 14492 6972 14544
rect 7288 14467 7340 14476
rect 7288 14433 7297 14467
rect 7297 14433 7331 14467
rect 7331 14433 7340 14467
rect 7748 14492 7800 14544
rect 8116 14492 8168 14544
rect 7288 14424 7340 14433
rect 8944 14424 8996 14476
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 6920 14356 6972 14408
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 7932 14356 7984 14408
rect 9128 14356 9180 14408
rect 10324 14424 10376 14476
rect 7380 14288 7432 14340
rect 8300 14288 8352 14340
rect 1584 14263 1636 14272
rect 1584 14229 1593 14263
rect 1593 14229 1627 14263
rect 1627 14229 1636 14263
rect 1584 14220 1636 14229
rect 6276 14220 6328 14272
rect 7288 14220 7340 14272
rect 8852 14220 8904 14272
rect 9404 14263 9456 14272
rect 9404 14229 9413 14263
rect 9413 14229 9447 14263
rect 9447 14229 9456 14263
rect 9404 14220 9456 14229
rect 4213 14118 4265 14170
rect 4277 14118 4329 14170
rect 4341 14118 4393 14170
rect 4405 14118 4457 14170
rect 4469 14118 4521 14170
rect 7477 14118 7529 14170
rect 7541 14118 7593 14170
rect 7605 14118 7657 14170
rect 7669 14118 7721 14170
rect 7733 14118 7785 14170
rect 5632 14059 5684 14068
rect 5632 14025 5641 14059
rect 5641 14025 5675 14059
rect 5675 14025 5684 14059
rect 5632 14016 5684 14025
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7104 14016 7156 14068
rect 8024 14016 8076 14068
rect 8392 14016 8444 14068
rect 9956 14016 10008 14068
rect 7656 13948 7708 14000
rect 9404 13948 9456 14000
rect 6736 13880 6788 13932
rect 7196 13812 7248 13864
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 9036 13880 9088 13932
rect 9680 13880 9732 13932
rect 7564 13812 7616 13821
rect 7656 13744 7708 13796
rect 9128 13812 9180 13864
rect 9956 13855 10008 13864
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 5632 13676 5684 13728
rect 7288 13676 7340 13728
rect 8300 13676 8352 13728
rect 2582 13574 2634 13626
rect 2646 13574 2698 13626
rect 2710 13574 2762 13626
rect 2774 13574 2826 13626
rect 2838 13574 2890 13626
rect 5845 13574 5897 13626
rect 5909 13574 5961 13626
rect 5973 13574 6025 13626
rect 6037 13574 6089 13626
rect 6101 13574 6153 13626
rect 9109 13574 9161 13626
rect 9173 13574 9225 13626
rect 9237 13574 9289 13626
rect 9301 13574 9353 13626
rect 9365 13574 9417 13626
rect 6828 13472 6880 13524
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 8300 13404 8352 13456
rect 5356 13379 5408 13388
rect 5356 13345 5365 13379
rect 5365 13345 5399 13379
rect 5399 13345 5408 13379
rect 5356 13336 5408 13345
rect 5632 13379 5684 13388
rect 5632 13345 5641 13379
rect 5641 13345 5675 13379
rect 5675 13345 5684 13379
rect 5632 13336 5684 13345
rect 7564 13336 7616 13388
rect 6092 13268 6144 13320
rect 6184 13268 6236 13320
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 6552 13132 6604 13184
rect 6736 13200 6788 13252
rect 8024 13268 8076 13320
rect 8668 13200 8720 13252
rect 9588 13404 9640 13456
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 9496 13132 9548 13184
rect 9772 13175 9824 13184
rect 9772 13141 9781 13175
rect 9781 13141 9815 13175
rect 9815 13141 9824 13175
rect 9772 13132 9824 13141
rect 4213 13030 4265 13082
rect 4277 13030 4329 13082
rect 4341 13030 4393 13082
rect 4405 13030 4457 13082
rect 4469 13030 4521 13082
rect 7477 13030 7529 13082
rect 7541 13030 7593 13082
rect 7605 13030 7657 13082
rect 7669 13030 7721 13082
rect 7733 13030 7785 13082
rect 7012 12928 7064 12980
rect 7380 12928 7432 12980
rect 7840 12928 7892 12980
rect 8944 12928 8996 12980
rect 9588 12928 9640 12980
rect 8208 12860 8260 12912
rect 8852 12860 8904 12912
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 7104 12792 7156 12844
rect 7380 12792 7432 12844
rect 8944 12792 8996 12844
rect 9404 12792 9456 12844
rect 8852 12724 8904 12776
rect 7012 12656 7064 12708
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 2582 12486 2634 12538
rect 2646 12486 2698 12538
rect 2710 12486 2762 12538
rect 2774 12486 2826 12538
rect 2838 12486 2890 12538
rect 5845 12486 5897 12538
rect 5909 12486 5961 12538
rect 5973 12486 6025 12538
rect 6037 12486 6089 12538
rect 6101 12486 6153 12538
rect 9109 12486 9161 12538
rect 9173 12486 9225 12538
rect 9237 12486 9289 12538
rect 9301 12486 9353 12538
rect 9365 12486 9417 12538
rect 940 12384 992 12436
rect 6184 12384 6236 12436
rect 6460 12384 6512 12436
rect 8024 12384 8076 12436
rect 8852 12384 8904 12436
rect 5816 12180 5868 12232
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 6368 12223 6420 12232
rect 5908 12180 5960 12189
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 6552 12180 6604 12189
rect 9680 12180 9732 12232
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 8392 12112 8444 12164
rect 9496 12112 9548 12164
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 9680 12044 9732 12096
rect 4213 11942 4265 11994
rect 4277 11942 4329 11994
rect 4341 11942 4393 11994
rect 4405 11942 4457 11994
rect 4469 11942 4521 11994
rect 7477 11942 7529 11994
rect 7541 11942 7593 11994
rect 7605 11942 7657 11994
rect 7669 11942 7721 11994
rect 7733 11942 7785 11994
rect 5816 11840 5868 11892
rect 8392 11840 8444 11892
rect 8484 11840 8536 11892
rect 9404 11772 9456 11824
rect 6644 11704 6696 11756
rect 6828 11747 6880 11756
rect 6828 11713 6862 11747
rect 6862 11713 6880 11747
rect 6828 11704 6880 11713
rect 8208 11704 8260 11756
rect 1400 11568 1452 11620
rect 6552 11568 6604 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 8116 11500 8168 11552
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5845 11398 5897 11450
rect 5909 11398 5961 11450
rect 5973 11398 6025 11450
rect 6037 11398 6089 11450
rect 6101 11398 6153 11450
rect 9109 11398 9161 11450
rect 9173 11398 9225 11450
rect 9237 11398 9289 11450
rect 9301 11398 9353 11450
rect 9365 11398 9417 11450
rect 6828 11296 6880 11348
rect 6552 11228 6604 11280
rect 7932 11296 7984 11348
rect 8944 11296 8996 11348
rect 9864 11296 9916 11348
rect 9772 11228 9824 11280
rect 9404 11160 9456 11212
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 7380 11024 7432 11076
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 4213 10854 4265 10906
rect 4277 10854 4329 10906
rect 4341 10854 4393 10906
rect 4405 10854 4457 10906
rect 4469 10854 4521 10906
rect 7477 10854 7529 10906
rect 7541 10854 7593 10906
rect 7605 10854 7657 10906
rect 7669 10854 7721 10906
rect 7733 10854 7785 10906
rect 5632 10752 5684 10804
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 8760 10684 8812 10736
rect 9496 10684 9548 10736
rect 7196 10616 7248 10668
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 8760 10548 8812 10600
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 7104 10480 7156 10532
rect 9404 10523 9456 10532
rect 9404 10489 9413 10523
rect 9413 10489 9447 10523
rect 9447 10489 9456 10523
rect 9404 10480 9456 10489
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 9772 10412 9824 10464
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5845 10310 5897 10362
rect 5909 10310 5961 10362
rect 5973 10310 6025 10362
rect 6037 10310 6089 10362
rect 6101 10310 6153 10362
rect 9109 10310 9161 10362
rect 9173 10310 9225 10362
rect 9237 10310 9289 10362
rect 9301 10310 9353 10362
rect 9365 10310 9417 10362
rect 7196 10251 7248 10260
rect 7196 10217 7205 10251
rect 7205 10217 7239 10251
rect 7239 10217 7248 10251
rect 7196 10208 7248 10217
rect 8760 10208 8812 10260
rect 9680 10140 9732 10192
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 4712 9936 4764 9988
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 4213 9766 4265 9818
rect 4277 9766 4329 9818
rect 4341 9766 4393 9818
rect 4405 9766 4457 9818
rect 4469 9766 4521 9818
rect 7477 9766 7529 9818
rect 7541 9766 7593 9818
rect 7605 9766 7657 9818
rect 7669 9766 7721 9818
rect 7733 9766 7785 9818
rect 8484 9596 8536 9648
rect 8852 9639 8904 9648
rect 8852 9605 8861 9639
rect 8861 9605 8895 9639
rect 8895 9605 8904 9639
rect 8852 9596 8904 9605
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 1860 9392 1912 9444
rect 8852 9392 8904 9444
rect 9220 9392 9272 9444
rect 5540 9324 5592 9376
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5845 9222 5897 9274
rect 5909 9222 5961 9274
rect 5973 9222 6025 9274
rect 6037 9222 6089 9274
rect 6101 9222 6153 9274
rect 9109 9222 9161 9274
rect 9173 9222 9225 9274
rect 9237 9222 9289 9274
rect 9301 9222 9353 9274
rect 9365 9222 9417 9274
rect 5448 9120 5500 9172
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 4213 8678 4265 8730
rect 4277 8678 4329 8730
rect 4341 8678 4393 8730
rect 4405 8678 4457 8730
rect 4469 8678 4521 8730
rect 7477 8678 7529 8730
rect 7541 8678 7593 8730
rect 7605 8678 7657 8730
rect 7669 8678 7721 8730
rect 7733 8678 7785 8730
rect 8944 8576 8996 8628
rect 9588 8508 9640 8560
rect 756 8440 808 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 1584 8304 1636 8313
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5845 8134 5897 8186
rect 5909 8134 5961 8186
rect 5973 8134 6025 8186
rect 6037 8134 6089 8186
rect 6101 8134 6153 8186
rect 9109 8134 9161 8186
rect 9173 8134 9225 8186
rect 9237 8134 9289 8186
rect 9301 8134 9353 8186
rect 9365 8134 9417 8186
rect 1676 7828 1728 7880
rect 9772 7803 9824 7812
rect 9772 7769 9781 7803
rect 9781 7769 9815 7803
rect 9815 7769 9824 7803
rect 9772 7760 9824 7769
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 4213 7590 4265 7642
rect 4277 7590 4329 7642
rect 4341 7590 4393 7642
rect 4405 7590 4457 7642
rect 4469 7590 4521 7642
rect 7477 7590 7529 7642
rect 7541 7590 7593 7642
rect 7605 7590 7657 7642
rect 7669 7590 7721 7642
rect 7733 7590 7785 7642
rect 5172 7488 5224 7540
rect 1216 7352 1268 7404
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9680 7352 9732 7404
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 8392 7216 8444 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 8576 7148 8628 7200
rect 8760 7148 8812 7200
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5845 7046 5897 7098
rect 5909 7046 5961 7098
rect 5973 7046 6025 7098
rect 6037 7046 6089 7098
rect 6101 7046 6153 7098
rect 9109 7046 9161 7098
rect 9173 7046 9225 7098
rect 9237 7046 9289 7098
rect 9301 7046 9353 7098
rect 9365 7046 9417 7098
rect 8852 6808 8904 6860
rect 9956 6851 10008 6860
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 9036 6672 9088 6724
rect 8668 6604 8720 6656
rect 4213 6502 4265 6554
rect 4277 6502 4329 6554
rect 4341 6502 4393 6554
rect 4405 6502 4457 6554
rect 4469 6502 4521 6554
rect 7477 6502 7529 6554
rect 7541 6502 7593 6554
rect 7605 6502 7657 6554
rect 7669 6502 7721 6554
rect 7733 6502 7785 6554
rect 8852 6400 8904 6452
rect 1492 6264 1544 6316
rect 6184 6264 6236 6316
rect 1584 6171 1636 6180
rect 1584 6137 1593 6171
rect 1593 6137 1627 6171
rect 1627 6137 1636 6171
rect 1584 6128 1636 6137
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5845 5958 5897 6010
rect 5909 5958 5961 6010
rect 5973 5958 6025 6010
rect 6037 5958 6089 6010
rect 6101 5958 6153 6010
rect 9109 5958 9161 6010
rect 9173 5958 9225 6010
rect 9237 5958 9289 6010
rect 9301 5958 9353 6010
rect 9365 5958 9417 6010
rect 8852 5720 8904 5772
rect 9956 5720 10008 5772
rect 5724 5652 5776 5704
rect 6736 5652 6788 5704
rect 8024 5652 8076 5704
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 8576 5516 8628 5568
rect 4213 5414 4265 5466
rect 4277 5414 4329 5466
rect 4341 5414 4393 5466
rect 4405 5414 4457 5466
rect 4469 5414 4521 5466
rect 7477 5414 7529 5466
rect 7541 5414 7593 5466
rect 7605 5414 7657 5466
rect 7669 5414 7721 5466
rect 7733 5414 7785 5466
rect 9680 5312 9732 5364
rect 1768 5176 1820 5228
rect 8116 5176 8168 5228
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 8760 5108 8812 5160
rect 9588 5108 9640 5160
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 5540 5040 5592 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5845 4870 5897 4922
rect 5909 4870 5961 4922
rect 5973 4870 6025 4922
rect 6037 4870 6089 4922
rect 6101 4870 6153 4922
rect 9109 4870 9161 4922
rect 9173 4870 9225 4922
rect 9237 4870 9289 4922
rect 9301 4870 9353 4922
rect 9365 4870 9417 4922
rect 9588 4768 9640 4820
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 8392 4564 8444 4616
rect 8760 4564 8812 4616
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 9404 4471 9456 4480
rect 9404 4437 9413 4471
rect 9413 4437 9447 4471
rect 9447 4437 9456 4471
rect 9404 4428 9456 4437
rect 4213 4326 4265 4378
rect 4277 4326 4329 4378
rect 4341 4326 4393 4378
rect 4405 4326 4457 4378
rect 4469 4326 4521 4378
rect 7477 4326 7529 4378
rect 7541 4326 7593 4378
rect 7605 4326 7657 4378
rect 7669 4326 7721 4378
rect 7733 4326 7785 4378
rect 8024 4224 8076 4276
rect 9404 4156 9456 4208
rect 9128 4088 9180 4140
rect 9496 4088 9548 4140
rect 8944 4020 8996 4072
rect 9220 4020 9272 4072
rect 9036 3952 9088 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5845 3782 5897 3834
rect 5909 3782 5961 3834
rect 5973 3782 6025 3834
rect 6037 3782 6089 3834
rect 6101 3782 6153 3834
rect 9109 3782 9161 3834
rect 9173 3782 9225 3834
rect 9237 3782 9289 3834
rect 9301 3782 9353 3834
rect 9365 3782 9417 3834
rect 9772 3680 9824 3732
rect 8668 3544 8720 3596
rect 8852 3544 8904 3596
rect 8116 3476 8168 3528
rect 9496 3476 9548 3528
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 4213 3238 4265 3290
rect 4277 3238 4329 3290
rect 4341 3238 4393 3290
rect 4405 3238 4457 3290
rect 4469 3238 4521 3290
rect 7477 3238 7529 3290
rect 7541 3238 7593 3290
rect 7605 3238 7657 3290
rect 7669 3238 7721 3290
rect 7733 3238 7785 3290
rect 9956 3136 10008 3188
rect 8576 3068 8628 3120
rect 8116 3000 8168 3052
rect 8944 2932 8996 2984
rect 7840 2907 7892 2916
rect 7840 2873 7849 2907
rect 7849 2873 7883 2907
rect 7883 2873 7892 2907
rect 7840 2864 7892 2873
rect 8300 2864 8352 2916
rect 8576 2864 8628 2916
rect 1400 2796 1452 2848
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5845 2694 5897 2746
rect 5909 2694 5961 2746
rect 5973 2694 6025 2746
rect 6037 2694 6089 2746
rect 6101 2694 6153 2746
rect 9109 2694 9161 2746
rect 9173 2694 9225 2746
rect 9237 2694 9289 2746
rect 9301 2694 9353 2746
rect 9365 2694 9417 2746
rect 1492 2388 1544 2440
rect 5540 2456 5592 2508
rect 7932 2456 7984 2508
rect 8484 2456 8536 2508
rect 7104 2388 7156 2440
rect 8576 2388 8628 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2320 2295 2372 2304
rect 2320 2261 2329 2295
rect 2329 2261 2363 2295
rect 2363 2261 2372 2295
rect 2320 2252 2372 2261
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 4213 2150 4265 2202
rect 4277 2150 4329 2202
rect 4341 2150 4393 2202
rect 4405 2150 4457 2202
rect 4469 2150 4521 2202
rect 7477 2150 7529 2202
rect 7541 2150 7593 2202
rect 7605 2150 7657 2202
rect 7669 2150 7721 2202
rect 7733 2150 7785 2202
<< metal2 >>
rect 3238 79656 3294 79665
rect 3238 79591 3294 79600
rect 7562 79656 7618 79665
rect 7562 79591 7618 79600
rect 1398 78976 1454 78985
rect 1398 78911 1454 78920
rect 1412 77586 1440 78911
rect 2962 78296 3018 78305
rect 2962 78231 3018 78240
rect 2582 77820 2890 77840
rect 2582 77818 2588 77820
rect 2644 77818 2668 77820
rect 2724 77818 2748 77820
rect 2804 77818 2828 77820
rect 2884 77818 2890 77820
rect 2644 77766 2646 77818
rect 2826 77766 2828 77818
rect 2582 77764 2588 77766
rect 2644 77764 2668 77766
rect 2724 77764 2748 77766
rect 2804 77764 2828 77766
rect 2884 77764 2890 77766
rect 2582 77744 2890 77764
rect 2870 77616 2926 77625
rect 1400 77580 1452 77586
rect 2870 77551 2926 77560
rect 1400 77522 1452 77528
rect 2884 77518 2912 77551
rect 2872 77512 2924 77518
rect 2872 77454 2924 77460
rect 2976 77110 3004 78231
rect 3148 77444 3200 77450
rect 3148 77386 3200 77392
rect 3056 77376 3108 77382
rect 3056 77318 3108 77324
rect 2964 77104 3016 77110
rect 2964 77046 3016 77052
rect 1584 77036 1636 77042
rect 1584 76978 1636 76984
rect 1596 76945 1624 76978
rect 1582 76936 1638 76945
rect 1582 76871 1638 76880
rect 2964 76900 3016 76906
rect 2964 76842 3016 76848
rect 2582 76732 2890 76752
rect 2582 76730 2588 76732
rect 2644 76730 2668 76732
rect 2724 76730 2748 76732
rect 2804 76730 2828 76732
rect 2884 76730 2890 76732
rect 2644 76678 2646 76730
rect 2826 76678 2828 76730
rect 2582 76676 2588 76678
rect 2644 76676 2668 76678
rect 2724 76676 2748 76678
rect 2804 76676 2828 76678
rect 2884 76676 2890 76678
rect 2582 76656 2890 76676
rect 1584 76424 1636 76430
rect 1584 76366 1636 76372
rect 1596 76265 1624 76366
rect 2136 76288 2188 76294
rect 1582 76256 1638 76265
rect 2136 76230 2188 76236
rect 1582 76191 1638 76200
rect 1768 75948 1820 75954
rect 1768 75890 1820 75896
rect 1400 75880 1452 75886
rect 1400 75822 1452 75828
rect 1412 75585 1440 75822
rect 1398 75576 1454 75585
rect 1398 75511 1454 75520
rect 1584 74860 1636 74866
rect 1584 74802 1636 74808
rect 1596 73681 1624 74802
rect 1582 73672 1638 73681
rect 1582 73607 1638 73616
rect 1676 73160 1728 73166
rect 1676 73102 1728 73108
rect 940 72684 992 72690
rect 940 72626 992 72632
rect 952 68882 980 72626
rect 1584 72072 1636 72078
rect 1584 72014 1636 72020
rect 1596 71641 1624 72014
rect 1582 71632 1638 71641
rect 1492 71596 1544 71602
rect 1582 71567 1638 71576
rect 1492 71538 1544 71544
rect 1400 70984 1452 70990
rect 1398 70952 1400 70961
rect 1452 70952 1454 70961
rect 1398 70887 1454 70896
rect 1504 70553 1532 71538
rect 1490 70544 1546 70553
rect 1490 70479 1546 70488
rect 1124 69896 1176 69902
rect 1124 69838 1176 69844
rect 940 68876 992 68882
rect 940 68818 992 68824
rect 848 59968 900 59974
rect 848 59910 900 59916
rect 664 59424 716 59430
rect 664 59366 716 59372
rect 388 53984 440 53990
rect 388 53926 440 53932
rect 400 43994 428 53926
rect 480 50856 532 50862
rect 480 50798 532 50804
rect 388 43988 440 43994
rect 388 43930 440 43936
rect 492 15910 520 50798
rect 572 49088 624 49094
rect 572 49030 624 49036
rect 584 38554 612 49030
rect 572 38548 624 38554
rect 572 38490 624 38496
rect 676 34542 704 59366
rect 756 47592 808 47598
rect 756 47534 808 47540
rect 664 34536 716 34542
rect 664 34478 716 34484
rect 480 15904 532 15910
rect 480 15846 532 15852
rect 768 8498 796 47534
rect 860 43926 888 59910
rect 952 51066 980 68818
rect 1032 63980 1084 63986
rect 1032 63922 1084 63928
rect 1044 63073 1072 63922
rect 1030 63064 1086 63073
rect 1030 62999 1086 63008
rect 1032 57044 1084 57050
rect 1032 56986 1084 56992
rect 940 51060 992 51066
rect 940 51002 992 51008
rect 848 43920 900 43926
rect 848 43862 900 43868
rect 940 41744 992 41750
rect 940 41686 992 41692
rect 952 12442 980 41686
rect 1044 25226 1072 56986
rect 1136 47258 1164 69838
rect 1216 69420 1268 69426
rect 1216 69362 1268 69368
rect 1228 50522 1256 69362
rect 1584 68808 1636 68814
rect 1584 68750 1636 68756
rect 1596 68377 1624 68750
rect 1582 68368 1638 68377
rect 1492 68332 1544 68338
rect 1582 68303 1638 68312
rect 1492 68274 1544 68280
rect 1308 68264 1360 68270
rect 1308 68206 1360 68212
rect 1216 50516 1268 50522
rect 1216 50458 1268 50464
rect 1124 47252 1176 47258
rect 1124 47194 1176 47200
rect 1320 46170 1348 68206
rect 1400 67720 1452 67726
rect 1398 67688 1400 67697
rect 1452 67688 1454 67697
rect 1398 67623 1454 67632
rect 1504 67017 1532 68274
rect 1584 68196 1636 68202
rect 1584 68138 1636 68144
rect 1490 67008 1546 67017
rect 1490 66943 1546 66952
rect 1596 66858 1624 68138
rect 1504 66830 1624 66858
rect 1400 64456 1452 64462
rect 1400 64398 1452 64404
rect 1412 63753 1440 64398
rect 1398 63744 1454 63753
rect 1398 63679 1454 63688
rect 1400 63368 1452 63374
rect 1400 63310 1452 63316
rect 1412 62393 1440 63310
rect 1398 62384 1454 62393
rect 1398 62319 1454 62328
rect 1400 61804 1452 61810
rect 1400 61746 1452 61752
rect 1412 61169 1440 61746
rect 1398 61160 1454 61169
rect 1398 61095 1454 61104
rect 1504 54194 1532 66830
rect 1582 65784 1638 65793
rect 1582 65719 1638 65728
rect 1596 65550 1624 65719
rect 1584 65544 1636 65550
rect 1584 65486 1636 65492
rect 1688 60654 1716 73102
rect 1780 73030 1808 75890
rect 1860 75268 1912 75274
rect 1860 75210 1912 75216
rect 1872 75041 1900 75210
rect 1952 75200 2004 75206
rect 1952 75142 2004 75148
rect 1858 75032 1914 75041
rect 1858 74967 1914 74976
rect 1964 73778 1992 75142
rect 2044 74656 2096 74662
rect 2044 74598 2096 74604
rect 1952 73772 2004 73778
rect 1952 73714 2004 73720
rect 1952 73636 2004 73642
rect 1952 73578 2004 73584
rect 1768 73024 1820 73030
rect 1768 72966 1820 72972
rect 1768 72820 1820 72826
rect 1768 72762 1820 72768
rect 1780 69902 1808 72762
rect 1860 72616 1912 72622
rect 1860 72558 1912 72564
rect 1872 69970 1900 72558
rect 1860 69964 1912 69970
rect 1860 69906 1912 69912
rect 1768 69896 1820 69902
rect 1768 69838 1820 69844
rect 1964 68202 1992 73578
rect 2056 72826 2084 74598
rect 2148 74118 2176 76230
rect 2582 75644 2890 75664
rect 2582 75642 2588 75644
rect 2644 75642 2668 75644
rect 2724 75642 2748 75644
rect 2804 75642 2828 75644
rect 2884 75642 2890 75644
rect 2644 75590 2646 75642
rect 2826 75590 2828 75642
rect 2582 75588 2588 75590
rect 2644 75588 2668 75590
rect 2724 75588 2748 75590
rect 2804 75588 2828 75590
rect 2884 75588 2890 75590
rect 2582 75568 2890 75588
rect 2228 74860 2280 74866
rect 2228 74802 2280 74808
rect 2240 74361 2268 74802
rect 2504 74792 2556 74798
rect 2504 74734 2556 74740
rect 2226 74352 2282 74361
rect 2516 74322 2544 74734
rect 2582 74556 2890 74576
rect 2582 74554 2588 74556
rect 2644 74554 2668 74556
rect 2724 74554 2748 74556
rect 2804 74554 2828 74556
rect 2884 74554 2890 74556
rect 2644 74502 2646 74554
rect 2826 74502 2828 74554
rect 2582 74500 2588 74502
rect 2644 74500 2668 74502
rect 2724 74500 2748 74502
rect 2804 74500 2828 74502
rect 2884 74500 2890 74502
rect 2582 74480 2890 74500
rect 2226 74287 2282 74296
rect 2504 74316 2556 74322
rect 2504 74258 2556 74264
rect 2320 74248 2372 74254
rect 2320 74190 2372 74196
rect 2136 74112 2188 74118
rect 2136 74054 2188 74060
rect 2148 73370 2176 74054
rect 2136 73364 2188 73370
rect 2136 73306 2188 73312
rect 2136 73024 2188 73030
rect 2136 72966 2188 72972
rect 2044 72820 2096 72826
rect 2044 72762 2096 72768
rect 2044 71936 2096 71942
rect 2044 71878 2096 71884
rect 2056 69562 2084 71878
rect 2148 71534 2176 72966
rect 2228 72752 2280 72758
rect 2228 72694 2280 72700
rect 2240 72622 2268 72694
rect 2228 72616 2280 72622
rect 2228 72558 2280 72564
rect 2226 72312 2282 72321
rect 2226 72247 2282 72256
rect 2240 72078 2268 72247
rect 2228 72072 2280 72078
rect 2228 72014 2280 72020
rect 2332 71618 2360 74190
rect 2412 73772 2464 73778
rect 2412 73714 2464 73720
rect 2240 71590 2360 71618
rect 2136 71528 2188 71534
rect 2136 71470 2188 71476
rect 2136 71052 2188 71058
rect 2136 70994 2188 71000
rect 2148 69902 2176 70994
rect 2240 70514 2268 71590
rect 2320 71528 2372 71534
rect 2320 71470 2372 71476
rect 2228 70508 2280 70514
rect 2228 70450 2280 70456
rect 2332 70394 2360 71470
rect 2240 70366 2360 70394
rect 2136 69896 2188 69902
rect 2136 69838 2188 69844
rect 2044 69556 2096 69562
rect 2044 69498 2096 69504
rect 1952 68196 2004 68202
rect 1952 68138 2004 68144
rect 1768 68128 1820 68134
rect 1768 68070 1820 68076
rect 1780 67386 1808 68070
rect 1952 67720 2004 67726
rect 1952 67662 2004 67668
rect 1768 67380 1820 67386
rect 1768 67322 1820 67328
rect 1780 66162 1808 67322
rect 1860 67176 1912 67182
rect 1860 67118 1912 67124
rect 1768 66156 1820 66162
rect 1768 66098 1820 66104
rect 1872 66094 1900 67118
rect 1860 66088 1912 66094
rect 1860 66030 1912 66036
rect 1860 65068 1912 65074
rect 1860 65010 1912 65016
rect 1872 64433 1900 65010
rect 1858 64424 1914 64433
rect 1858 64359 1914 64368
rect 1768 63776 1820 63782
rect 1768 63718 1820 63724
rect 1676 60648 1728 60654
rect 1676 60590 1728 60596
rect 1584 60512 1636 60518
rect 1584 60454 1636 60460
rect 1596 59537 1624 60454
rect 1582 59528 1638 59537
rect 1582 59463 1638 59472
rect 1582 58440 1638 58449
rect 1582 58375 1584 58384
rect 1636 58375 1638 58384
rect 1584 58346 1636 58352
rect 1584 57792 1636 57798
rect 1582 57760 1584 57769
rect 1636 57760 1638 57769
rect 1582 57695 1638 57704
rect 1676 57520 1728 57526
rect 1676 57462 1728 57468
rect 1584 57248 1636 57254
rect 1584 57190 1636 57196
rect 1596 57089 1624 57190
rect 1582 57080 1638 57089
rect 1582 57015 1638 57024
rect 1584 56704 1636 56710
rect 1584 56646 1636 56652
rect 1596 56545 1624 56646
rect 1582 56536 1638 56545
rect 1582 56471 1638 56480
rect 1584 56160 1636 56166
rect 1584 56102 1636 56108
rect 1596 55865 1624 56102
rect 1582 55856 1638 55865
rect 1582 55791 1638 55800
rect 1584 55616 1636 55622
rect 1584 55558 1636 55564
rect 1596 55185 1624 55558
rect 1582 55176 1638 55185
rect 1582 55111 1638 55120
rect 1584 55072 1636 55078
rect 1584 55014 1636 55020
rect 1596 54505 1624 55014
rect 1688 54874 1716 57462
rect 1676 54868 1728 54874
rect 1676 54810 1728 54816
rect 1676 54528 1728 54534
rect 1582 54496 1638 54505
rect 1676 54470 1728 54476
rect 1582 54431 1638 54440
rect 1492 54188 1544 54194
rect 1492 54130 1544 54136
rect 1582 53816 1638 53825
rect 1582 53751 1584 53760
rect 1636 53751 1638 53760
rect 1584 53722 1636 53728
rect 1492 53576 1544 53582
rect 1492 53518 1544 53524
rect 1400 51400 1452 51406
rect 1400 51342 1452 51348
rect 1412 51241 1440 51342
rect 1398 51232 1454 51241
rect 1398 51167 1454 51176
rect 1308 46164 1360 46170
rect 1308 46106 1360 46112
rect 1400 45484 1452 45490
rect 1400 45426 1452 45432
rect 1412 45257 1440 45426
rect 1504 45354 1532 53518
rect 1584 53236 1636 53242
rect 1584 53178 1636 53184
rect 1596 53145 1624 53178
rect 1582 53136 1638 53145
rect 1582 53071 1638 53080
rect 1688 52494 1716 54470
rect 1676 52488 1728 52494
rect 1676 52430 1728 52436
rect 1584 48680 1636 48686
rect 1584 48622 1636 48628
rect 1492 45348 1544 45354
rect 1492 45290 1544 45296
rect 1398 45248 1454 45257
rect 1398 45183 1454 45192
rect 1596 45082 1624 48622
rect 1584 45076 1636 45082
rect 1584 45018 1636 45024
rect 1584 44328 1636 44334
rect 1584 44270 1636 44276
rect 1492 43988 1544 43994
rect 1492 43930 1544 43936
rect 1216 43716 1268 43722
rect 1216 43658 1268 43664
rect 1124 43172 1176 43178
rect 1124 43114 1176 43120
rect 1136 35894 1164 43114
rect 1228 37210 1256 43658
rect 1400 42696 1452 42702
rect 1398 42664 1400 42673
rect 1452 42664 1454 42673
rect 1398 42599 1454 42608
rect 1400 42220 1452 42226
rect 1400 42162 1452 42168
rect 1412 41993 1440 42162
rect 1398 41984 1454 41993
rect 1398 41919 1454 41928
rect 1400 41608 1452 41614
rect 1400 41550 1452 41556
rect 1412 41313 1440 41550
rect 1398 41304 1454 41313
rect 1398 41239 1454 41248
rect 1308 41064 1360 41070
rect 1308 41006 1360 41012
rect 1320 38434 1348 41006
rect 1400 39976 1452 39982
rect 1398 39944 1400 39953
rect 1452 39944 1454 39953
rect 1398 39879 1454 39888
rect 1504 38978 1532 43930
rect 1596 42362 1624 44270
rect 1584 42356 1636 42362
rect 1584 42298 1636 42304
rect 1584 40112 1636 40118
rect 1584 40054 1636 40060
rect 1596 39098 1624 40054
rect 1688 40050 1716 52430
rect 1780 45422 1808 63718
rect 1860 62212 1912 62218
rect 1860 62154 1912 62160
rect 1872 61713 1900 62154
rect 1858 61704 1914 61713
rect 1858 61639 1914 61648
rect 1860 60036 1912 60042
rect 1860 59978 1912 59984
rect 1872 59809 1900 59978
rect 1858 59800 1914 59809
rect 1858 59735 1914 59744
rect 1860 59628 1912 59634
rect 1860 59570 1912 59576
rect 1872 59129 1900 59570
rect 1858 59120 1914 59129
rect 1858 59055 1914 59064
rect 1860 57384 1912 57390
rect 1860 57326 1912 57332
rect 1872 52154 1900 57326
rect 1964 54738 1992 67662
rect 2056 66620 2084 69498
rect 2148 69358 2176 69838
rect 2136 69352 2188 69358
rect 2136 69294 2188 69300
rect 2136 66632 2188 66638
rect 2056 66592 2136 66620
rect 2136 66574 2188 66580
rect 2240 66484 2268 70366
rect 2320 68672 2372 68678
rect 2320 68614 2372 68620
rect 2056 66456 2268 66484
rect 2056 60858 2084 66456
rect 2228 65544 2280 65550
rect 2228 65486 2280 65492
rect 2240 65113 2268 65486
rect 2226 65104 2282 65113
rect 2226 65039 2282 65048
rect 2332 63034 2360 68614
rect 2320 63028 2372 63034
rect 2320 62970 2372 62976
rect 2228 62824 2280 62830
rect 2228 62766 2280 62772
rect 2240 61266 2268 62766
rect 2228 61260 2280 61266
rect 2228 61202 2280 61208
rect 2332 61198 2360 62970
rect 2320 61192 2372 61198
rect 2320 61134 2372 61140
rect 2044 60852 2096 60858
rect 2044 60794 2096 60800
rect 2044 60648 2096 60654
rect 2044 60590 2096 60596
rect 1952 54732 2004 54738
rect 1952 54674 2004 54680
rect 1952 54188 2004 54194
rect 1952 54130 2004 54136
rect 1860 52148 1912 52154
rect 1860 52090 1912 52096
rect 1860 52012 1912 52018
rect 1860 51954 1912 51960
rect 1872 51921 1900 51954
rect 1858 51912 1914 51921
rect 1858 51847 1914 51856
rect 1860 50924 1912 50930
rect 1860 50866 1912 50872
rect 1872 50561 1900 50866
rect 1858 50552 1914 50561
rect 1858 50487 1914 50496
rect 1860 50244 1912 50250
rect 1860 50186 1912 50192
rect 1872 49881 1900 50186
rect 1858 49872 1914 49881
rect 1858 49807 1914 49816
rect 1860 49224 1912 49230
rect 1858 49192 1860 49201
rect 1912 49192 1914 49201
rect 1858 49127 1914 49136
rect 1860 48748 1912 48754
rect 1860 48690 1912 48696
rect 1872 48521 1900 48690
rect 1858 48512 1914 48521
rect 1858 48447 1914 48456
rect 1860 48068 1912 48074
rect 1860 48010 1912 48016
rect 1872 47841 1900 48010
rect 1858 47832 1914 47841
rect 1964 47802 1992 54130
rect 2056 48278 2084 60590
rect 2228 55276 2280 55282
rect 2228 55218 2280 55224
rect 2136 54732 2188 54738
rect 2136 54674 2188 54680
rect 2148 52426 2176 54674
rect 2136 52420 2188 52426
rect 2136 52362 2188 52368
rect 2044 48272 2096 48278
rect 2044 48214 2096 48220
rect 2136 48272 2188 48278
rect 2136 48214 2188 48220
rect 1858 47767 1914 47776
rect 1952 47796 2004 47802
rect 1952 47738 2004 47744
rect 1860 47660 1912 47666
rect 1860 47602 1912 47608
rect 1872 47297 1900 47602
rect 1858 47288 1914 47297
rect 1858 47223 1914 47232
rect 1860 46980 1912 46986
rect 1860 46922 1912 46928
rect 1872 46617 1900 46922
rect 1858 46608 1914 46617
rect 1858 46543 1914 46552
rect 1860 45960 1912 45966
rect 1858 45928 1860 45937
rect 1912 45928 1914 45937
rect 1858 45863 1914 45872
rect 1952 45552 2004 45558
rect 1952 45494 2004 45500
rect 1768 45416 1820 45422
rect 1768 45358 1820 45364
rect 1768 45076 1820 45082
rect 1768 45018 1820 45024
rect 1676 40044 1728 40050
rect 1676 39986 1728 39992
rect 1676 39568 1728 39574
rect 1676 39510 1728 39516
rect 1584 39092 1636 39098
rect 1584 39034 1636 39040
rect 1400 38956 1452 38962
rect 1504 38950 1624 38978
rect 1400 38898 1452 38904
rect 1412 38593 1440 38898
rect 1398 38584 1454 38593
rect 1398 38519 1454 38528
rect 1320 38406 1532 38434
rect 1400 38344 1452 38350
rect 1400 38286 1452 38292
rect 1412 37913 1440 38286
rect 1398 37904 1454 37913
rect 1308 37868 1360 37874
rect 1398 37839 1454 37848
rect 1308 37810 1360 37816
rect 1320 37369 1348 37810
rect 1306 37360 1362 37369
rect 1306 37295 1362 37304
rect 1228 37182 1348 37210
rect 1136 35866 1256 35894
rect 1032 25220 1084 25226
rect 1032 25162 1084 25168
rect 940 12436 992 12442
rect 940 12378 992 12384
rect 756 8492 808 8498
rect 756 8434 808 8440
rect 1228 7410 1256 35866
rect 1320 31770 1348 37182
rect 1400 36712 1452 36718
rect 1398 36680 1400 36689
rect 1452 36680 1454 36689
rect 1398 36615 1454 36624
rect 1400 36032 1452 36038
rect 1400 35974 1452 35980
rect 1412 35290 1440 35974
rect 1400 35284 1452 35290
rect 1400 35226 1452 35232
rect 1400 33992 1452 33998
rect 1398 33960 1400 33969
rect 1452 33960 1454 33969
rect 1398 33895 1454 33904
rect 1400 33448 1452 33454
rect 1400 33390 1452 33396
rect 1412 33289 1440 33390
rect 1398 33280 1454 33289
rect 1398 33215 1454 33224
rect 1320 31742 1440 31770
rect 1412 21350 1440 31742
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1412 18290 1440 18566
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1400 11620 1452 11626
rect 1400 11562 1452 11568
rect 1216 7404 1268 7410
rect 1216 7346 1268 7352
rect 1412 4706 1440 11562
rect 1504 6322 1532 38406
rect 1596 36786 1624 38950
rect 1584 36780 1636 36786
rect 1584 36722 1636 36728
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1596 36009 1624 36110
rect 1582 36000 1638 36009
rect 1582 35935 1638 35944
rect 1584 35692 1636 35698
rect 1584 35634 1636 35640
rect 1596 35329 1624 35634
rect 1582 35320 1638 35329
rect 1582 35255 1638 35264
rect 1584 35080 1636 35086
rect 1584 35022 1636 35028
rect 1596 34649 1624 35022
rect 1582 34640 1638 34649
rect 1582 34575 1638 34584
rect 1584 32904 1636 32910
rect 1584 32846 1636 32852
rect 1596 32745 1624 32846
rect 1582 32736 1638 32745
rect 1582 32671 1638 32680
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1596 32065 1624 32370
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1596 31385 1624 31758
rect 1582 31376 1638 31385
rect 1582 31311 1638 31320
rect 1582 30696 1638 30705
rect 1582 30631 1638 30640
rect 1596 30598 1624 30631
rect 1584 30592 1636 30598
rect 1584 30534 1636 30540
rect 1584 30048 1636 30054
rect 1582 30016 1584 30025
rect 1636 30016 1638 30025
rect 1582 29951 1638 29960
rect 1584 29504 1636 29510
rect 1584 29446 1636 29452
rect 1596 29345 1624 29446
rect 1582 29336 1638 29345
rect 1582 29271 1638 29280
rect 1584 29028 1636 29034
rect 1584 28970 1636 28976
rect 1596 28665 1624 28970
rect 1582 28656 1638 28665
rect 1582 28591 1638 28600
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 1596 28121 1624 28358
rect 1582 28112 1638 28121
rect 1582 28047 1638 28056
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 1596 27334 1624 27367
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1584 26784 1636 26790
rect 1582 26752 1584 26761
rect 1636 26752 1638 26761
rect 1582 26687 1638 26696
rect 1584 26240 1636 26246
rect 1584 26182 1636 26188
rect 1596 26081 1624 26182
rect 1582 26072 1638 26081
rect 1582 26007 1638 26016
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1596 25401 1624 25638
rect 1582 25392 1638 25401
rect 1582 25327 1638 25336
rect 1582 24712 1638 24721
rect 1582 24647 1584 24656
rect 1636 24647 1638 24656
rect 1584 24618 1636 24624
rect 1584 24064 1636 24070
rect 1582 24032 1584 24041
rect 1636 24032 1638 24041
rect 1582 23967 1638 23976
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1596 22817 1624 22918
rect 1582 22808 1638 22817
rect 1582 22743 1638 22752
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22137 1624 22374
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 1582 21448 1638 21457
rect 1582 21383 1584 21392
rect 1636 21383 1638 21392
rect 1584 21354 1636 21360
rect 1584 20800 1636 20806
rect 1582 20768 1584 20777
rect 1636 20768 1638 20777
rect 1582 20703 1638 20712
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20097 1624 20198
rect 1582 20088 1638 20097
rect 1582 20023 1638 20032
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1596 19417 1624 19654
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1596 18873 1624 19110
rect 1582 18864 1638 18873
rect 1582 18799 1638 18808
rect 1582 18184 1638 18193
rect 1582 18119 1584 18128
rect 1636 18119 1638 18128
rect 1584 18090 1636 18096
rect 1584 17536 1636 17542
rect 1582 17504 1584 17513
rect 1636 17504 1638 17513
rect 1582 17439 1638 17448
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16833 1624 16934
rect 1582 16824 1638 16833
rect 1582 16759 1638 16768
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16153 1624 16390
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1582 15464 1638 15473
rect 1582 15399 1638 15408
rect 1596 15366 1624 15399
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1584 14816 1636 14822
rect 1582 14784 1584 14793
rect 1636 14784 1638 14793
rect 1582 14719 1638 14728
rect 1584 14272 1636 14278
rect 1582 14240 1584 14249
rect 1636 14240 1638 14249
rect 1582 14175 1638 14184
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 13569 1624 13670
rect 1582 13560 1638 13569
rect 1582 13495 1638 13504
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12889 1624 13126
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1582 12200 1638 12209
rect 1582 12135 1638 12144
rect 1596 12102 1624 12135
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1584 11552 1636 11558
rect 1582 11520 1584 11529
rect 1636 11520 1638 11529
rect 1582 11455 1638 11464
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10849 1624 10950
rect 1582 10840 1638 10849
rect 1582 10775 1638 10784
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10169 1624 10406
rect 1582 10160 1638 10169
rect 1582 10095 1638 10104
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9625 1624 9862
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8838 1624 8871
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 8265 1624 8298
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1688 7886 1716 39510
rect 1780 39114 1808 45018
rect 1860 44804 1912 44810
rect 1860 44746 1912 44752
rect 1872 44577 1900 44746
rect 1858 44568 1914 44577
rect 1858 44503 1914 44512
rect 1860 44396 1912 44402
rect 1860 44338 1912 44344
rect 1872 43897 1900 44338
rect 1858 43888 1914 43897
rect 1858 43823 1914 43832
rect 1860 43308 1912 43314
rect 1860 43250 1912 43256
rect 1872 43217 1900 43250
rect 1858 43208 1914 43217
rect 1858 43143 1914 43152
rect 1860 41132 1912 41138
rect 1860 41074 1912 41080
rect 1872 40633 1900 41074
rect 1858 40624 1914 40633
rect 1858 40559 1914 40568
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 39273 1900 40394
rect 1858 39264 1914 39273
rect 1858 39199 1914 39208
rect 1780 39086 1900 39114
rect 1768 37120 1820 37126
rect 1768 37062 1820 37068
rect 1780 36922 1808 37062
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7585 1624 7686
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1582 6216 1638 6225
rect 1582 6151 1584 6160
rect 1636 6151 1638 6160
rect 1584 6122 1636 6128
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1582 5471 1638 5480
rect 1780 5234 1808 21286
rect 1872 9450 1900 39086
rect 1964 38826 1992 45494
rect 2044 44260 2096 44266
rect 2044 44202 2096 44208
rect 2056 40662 2084 44202
rect 2148 41206 2176 48214
rect 2240 47802 2268 55218
rect 2320 54596 2372 54602
rect 2320 54538 2372 54544
rect 2332 54210 2360 54538
rect 2424 54330 2452 73714
rect 2516 73710 2544 74258
rect 2504 73704 2556 73710
rect 2504 73646 2556 73652
rect 2516 73234 2544 73646
rect 2582 73468 2890 73488
rect 2582 73466 2588 73468
rect 2644 73466 2668 73468
rect 2724 73466 2748 73468
rect 2804 73466 2828 73468
rect 2884 73466 2890 73468
rect 2644 73414 2646 73466
rect 2826 73414 2828 73466
rect 2582 73412 2588 73414
rect 2644 73412 2668 73414
rect 2724 73412 2748 73414
rect 2804 73412 2828 73414
rect 2884 73412 2890 73414
rect 2582 73392 2890 73412
rect 2596 73296 2648 73302
rect 2596 73238 2648 73244
rect 2504 73228 2556 73234
rect 2504 73170 2556 73176
rect 2516 72758 2544 73170
rect 2504 72752 2556 72758
rect 2504 72694 2556 72700
rect 2608 72570 2636 73238
rect 2872 73160 2924 73166
rect 2872 73102 2924 73108
rect 2884 73001 2912 73102
rect 2870 72992 2926 73001
rect 2870 72927 2926 72936
rect 2976 72690 3004 76842
rect 3068 75002 3096 77318
rect 3056 74996 3108 75002
rect 3056 74938 3108 74944
rect 2964 72684 3016 72690
rect 2964 72626 3016 72632
rect 2516 72542 2636 72570
rect 2516 70650 2544 72542
rect 2582 72380 2890 72400
rect 2582 72378 2588 72380
rect 2644 72378 2668 72380
rect 2724 72378 2748 72380
rect 2804 72378 2828 72380
rect 2884 72378 2890 72380
rect 2644 72326 2646 72378
rect 2826 72326 2828 72378
rect 2582 72324 2588 72326
rect 2644 72324 2668 72326
rect 2724 72324 2748 72326
rect 2804 72324 2828 72326
rect 2884 72324 2890 72326
rect 2582 72304 2890 72324
rect 2582 71292 2890 71312
rect 2582 71290 2588 71292
rect 2644 71290 2668 71292
rect 2724 71290 2748 71292
rect 2804 71290 2828 71292
rect 2884 71290 2890 71292
rect 2644 71238 2646 71290
rect 2826 71238 2828 71290
rect 2582 71236 2588 71238
rect 2644 71236 2668 71238
rect 2724 71236 2748 71238
rect 2804 71236 2828 71238
rect 2884 71236 2890 71238
rect 2582 71216 2890 71236
rect 2596 71052 2648 71058
rect 2596 70994 2648 71000
rect 2504 70644 2556 70650
rect 2504 70586 2556 70592
rect 2608 70514 2636 70994
rect 2596 70508 2648 70514
rect 2596 70450 2648 70456
rect 2582 70204 2890 70224
rect 2582 70202 2588 70204
rect 2644 70202 2668 70204
rect 2724 70202 2748 70204
rect 2804 70202 2828 70204
rect 2884 70202 2890 70204
rect 2644 70150 2646 70202
rect 2826 70150 2828 70202
rect 2582 70148 2588 70150
rect 2644 70148 2668 70150
rect 2724 70148 2748 70150
rect 2804 70148 2828 70150
rect 2884 70148 2890 70150
rect 2582 70128 2890 70148
rect 2872 69896 2924 69902
rect 2872 69838 2924 69844
rect 2884 69329 2912 69838
rect 2870 69320 2926 69329
rect 2504 69284 2556 69290
rect 2870 69255 2926 69264
rect 2504 69226 2556 69232
rect 2516 68746 2544 69226
rect 2582 69116 2890 69136
rect 2582 69114 2588 69116
rect 2644 69114 2668 69116
rect 2724 69114 2748 69116
rect 2804 69114 2828 69116
rect 2884 69114 2890 69116
rect 2644 69062 2646 69114
rect 2826 69062 2828 69114
rect 2582 69060 2588 69062
rect 2644 69060 2668 69062
rect 2724 69060 2748 69062
rect 2804 69060 2828 69062
rect 2884 69060 2890 69062
rect 2582 69040 2890 69060
rect 2976 68882 3004 72626
rect 3068 69426 3096 74938
rect 3160 74934 3188 77386
rect 3252 77042 3280 79591
rect 5845 77820 6153 77840
rect 5845 77818 5851 77820
rect 5907 77818 5931 77820
rect 5987 77818 6011 77820
rect 6067 77818 6091 77820
rect 6147 77818 6153 77820
rect 5907 77766 5909 77818
rect 6089 77766 6091 77818
rect 5845 77764 5851 77766
rect 5907 77764 5931 77766
rect 5987 77764 6011 77766
rect 6067 77764 6091 77766
rect 6147 77764 6153 77766
rect 5845 77744 6153 77764
rect 7576 77722 7604 79591
rect 8574 79248 8630 79257
rect 8574 79183 8630 79192
rect 8206 78296 8262 78305
rect 8206 78231 8262 78240
rect 8220 77722 8248 78231
rect 7564 77716 7616 77722
rect 7564 77658 7616 77664
rect 8208 77716 8260 77722
rect 8208 77658 8260 77664
rect 6184 77512 6236 77518
rect 6184 77454 6236 77460
rect 4213 77276 4521 77296
rect 4213 77274 4219 77276
rect 4275 77274 4299 77276
rect 4355 77274 4379 77276
rect 4435 77274 4459 77276
rect 4515 77274 4521 77276
rect 4275 77222 4277 77274
rect 4457 77222 4459 77274
rect 4213 77220 4219 77222
rect 4275 77220 4299 77222
rect 4355 77220 4379 77222
rect 4435 77220 4459 77222
rect 4515 77220 4521 77222
rect 4213 77200 4521 77220
rect 3700 77172 3752 77178
rect 3700 77114 3752 77120
rect 3240 77036 3292 77042
rect 3240 76978 3292 76984
rect 3332 76968 3384 76974
rect 3332 76910 3384 76916
rect 3148 74928 3200 74934
rect 3148 74870 3200 74876
rect 3148 74792 3200 74798
rect 3148 74734 3200 74740
rect 3160 74534 3188 74734
rect 3160 74506 3280 74534
rect 3148 72208 3200 72214
rect 3148 72150 3200 72156
rect 3056 69420 3108 69426
rect 3056 69362 3108 69368
rect 2964 68876 3016 68882
rect 2964 68818 3016 68824
rect 2504 68740 2556 68746
rect 2504 68682 2556 68688
rect 2516 68202 2544 68682
rect 2504 68196 2556 68202
rect 2504 68138 2556 68144
rect 2516 67182 2544 68138
rect 2582 68028 2890 68048
rect 2582 68026 2588 68028
rect 2644 68026 2668 68028
rect 2724 68026 2748 68028
rect 2804 68026 2828 68028
rect 2884 68026 2890 68028
rect 2644 67974 2646 68026
rect 2826 67974 2828 68026
rect 2582 67972 2588 67974
rect 2644 67972 2668 67974
rect 2724 67972 2748 67974
rect 2804 67972 2828 67974
rect 2884 67972 2890 67974
rect 2582 67952 2890 67972
rect 2964 67244 3016 67250
rect 2964 67186 3016 67192
rect 2504 67176 2556 67182
rect 2504 67118 2556 67124
rect 2516 66638 2544 67118
rect 2582 66940 2890 66960
rect 2582 66938 2588 66940
rect 2644 66938 2668 66940
rect 2724 66938 2748 66940
rect 2804 66938 2828 66940
rect 2884 66938 2890 66940
rect 2644 66886 2646 66938
rect 2826 66886 2828 66938
rect 2582 66884 2588 66886
rect 2644 66884 2668 66886
rect 2724 66884 2748 66886
rect 2804 66884 2828 66886
rect 2884 66884 2890 66886
rect 2582 66864 2890 66884
rect 2504 66632 2556 66638
rect 2504 66574 2556 66580
rect 2516 66162 2544 66574
rect 2976 66337 3004 67186
rect 2962 66328 3018 66337
rect 2962 66263 3018 66272
rect 3160 66230 3188 72150
rect 3252 70394 3280 74506
rect 3344 73914 3372 76910
rect 3332 73908 3384 73914
rect 3332 73850 3384 73856
rect 3712 73778 3740 77114
rect 5845 76732 6153 76752
rect 5845 76730 5851 76732
rect 5907 76730 5931 76732
rect 5987 76730 6011 76732
rect 6067 76730 6091 76732
rect 6147 76730 6153 76732
rect 5907 76678 5909 76730
rect 6089 76678 6091 76730
rect 5845 76676 5851 76678
rect 5907 76676 5931 76678
rect 5987 76676 6011 76678
rect 6067 76676 6091 76678
rect 6147 76676 6153 76678
rect 5845 76656 6153 76676
rect 4213 76188 4521 76208
rect 4213 76186 4219 76188
rect 4275 76186 4299 76188
rect 4355 76186 4379 76188
rect 4435 76186 4459 76188
rect 4515 76186 4521 76188
rect 4275 76134 4277 76186
rect 4457 76134 4459 76186
rect 4213 76132 4219 76134
rect 4275 76132 4299 76134
rect 4355 76132 4379 76134
rect 4435 76132 4459 76134
rect 4515 76132 4521 76134
rect 4213 76112 4521 76132
rect 5845 75644 6153 75664
rect 5845 75642 5851 75644
rect 5907 75642 5931 75644
rect 5987 75642 6011 75644
rect 6067 75642 6091 75644
rect 6147 75642 6153 75644
rect 5907 75590 5909 75642
rect 6089 75590 6091 75642
rect 5845 75588 5851 75590
rect 5907 75588 5931 75590
rect 5987 75588 6011 75590
rect 6067 75588 6091 75590
rect 6147 75588 6153 75590
rect 5845 75568 6153 75588
rect 4213 75100 4521 75120
rect 4213 75098 4219 75100
rect 4275 75098 4299 75100
rect 4355 75098 4379 75100
rect 4435 75098 4459 75100
rect 4515 75098 4521 75100
rect 4275 75046 4277 75098
rect 4457 75046 4459 75098
rect 4213 75044 4219 75046
rect 4275 75044 4299 75046
rect 4355 75044 4379 75046
rect 4435 75044 4459 75046
rect 4515 75044 4521 75046
rect 4213 75024 4521 75044
rect 4620 74656 4672 74662
rect 4620 74598 4672 74604
rect 4213 74012 4521 74032
rect 4213 74010 4219 74012
rect 4275 74010 4299 74012
rect 4355 74010 4379 74012
rect 4435 74010 4459 74012
rect 4515 74010 4521 74012
rect 4275 73958 4277 74010
rect 4457 73958 4459 74010
rect 4213 73956 4219 73958
rect 4275 73956 4299 73958
rect 4355 73956 4379 73958
rect 4435 73956 4459 73958
rect 4515 73956 4521 73958
rect 4213 73936 4521 73956
rect 3700 73772 3752 73778
rect 3700 73714 3752 73720
rect 4068 73772 4120 73778
rect 4068 73714 4120 73720
rect 3712 72146 3740 73714
rect 3700 72140 3752 72146
rect 3700 72082 3752 72088
rect 4080 72078 4108 73714
rect 4213 72924 4521 72944
rect 4213 72922 4219 72924
rect 4275 72922 4299 72924
rect 4355 72922 4379 72924
rect 4435 72922 4459 72924
rect 4515 72922 4521 72924
rect 4275 72870 4277 72922
rect 4457 72870 4459 72922
rect 4213 72868 4219 72870
rect 4275 72868 4299 72870
rect 4355 72868 4379 72870
rect 4435 72868 4459 72870
rect 4515 72868 4521 72870
rect 4213 72848 4521 72868
rect 4068 72072 4120 72078
rect 4068 72014 4120 72020
rect 3884 70848 3936 70854
rect 3884 70790 3936 70796
rect 3252 70366 3372 70394
rect 3344 69494 3372 70366
rect 3516 69828 3568 69834
rect 3516 69770 3568 69776
rect 3332 69488 3384 69494
rect 3332 69430 3384 69436
rect 3424 69216 3476 69222
rect 3424 69158 3476 69164
rect 3240 68740 3292 68746
rect 3240 68682 3292 68688
rect 3056 66224 3108 66230
rect 3056 66166 3108 66172
rect 3148 66224 3200 66230
rect 3148 66166 3200 66172
rect 2504 66156 2556 66162
rect 2504 66098 2556 66104
rect 2964 66088 3016 66094
rect 2964 66030 3016 66036
rect 2582 65852 2890 65872
rect 2582 65850 2588 65852
rect 2644 65850 2668 65852
rect 2724 65850 2748 65852
rect 2804 65850 2828 65852
rect 2884 65850 2890 65852
rect 2644 65798 2646 65850
rect 2826 65798 2828 65850
rect 2582 65796 2588 65798
rect 2644 65796 2668 65798
rect 2724 65796 2748 65798
rect 2804 65796 2828 65798
rect 2884 65796 2890 65798
rect 2582 65776 2890 65796
rect 2582 64764 2890 64784
rect 2582 64762 2588 64764
rect 2644 64762 2668 64764
rect 2724 64762 2748 64764
rect 2804 64762 2828 64764
rect 2884 64762 2890 64764
rect 2644 64710 2646 64762
rect 2826 64710 2828 64762
rect 2582 64708 2588 64710
rect 2644 64708 2668 64710
rect 2724 64708 2748 64710
rect 2804 64708 2828 64710
rect 2884 64708 2890 64710
rect 2582 64688 2890 64708
rect 2582 63676 2890 63696
rect 2582 63674 2588 63676
rect 2644 63674 2668 63676
rect 2724 63674 2748 63676
rect 2804 63674 2828 63676
rect 2884 63674 2890 63676
rect 2644 63622 2646 63674
rect 2826 63622 2828 63674
rect 2582 63620 2588 63622
rect 2644 63620 2668 63622
rect 2724 63620 2748 63622
rect 2804 63620 2828 63622
rect 2884 63620 2890 63622
rect 2582 63600 2890 63620
rect 2596 63504 2648 63510
rect 2596 63446 2648 63452
rect 2504 63368 2556 63374
rect 2504 63310 2556 63316
rect 2516 62830 2544 63310
rect 2504 62824 2556 62830
rect 2608 62801 2636 63446
rect 2976 63442 3004 66030
rect 3068 65754 3096 66166
rect 3056 65748 3108 65754
rect 3056 65690 3108 65696
rect 2964 63436 3016 63442
rect 2964 63378 3016 63384
rect 2504 62766 2556 62772
rect 2594 62792 2650 62801
rect 2516 61198 2544 62766
rect 2594 62727 2650 62736
rect 2582 62588 2890 62608
rect 2582 62586 2588 62588
rect 2644 62586 2668 62588
rect 2724 62586 2748 62588
rect 2804 62586 2828 62588
rect 2884 62586 2890 62588
rect 2644 62534 2646 62586
rect 2826 62534 2828 62586
rect 2582 62532 2588 62534
rect 2644 62532 2668 62534
rect 2724 62532 2748 62534
rect 2804 62532 2828 62534
rect 2884 62532 2890 62534
rect 2582 62512 2890 62532
rect 2582 61500 2890 61520
rect 2582 61498 2588 61500
rect 2644 61498 2668 61500
rect 2724 61498 2748 61500
rect 2804 61498 2828 61500
rect 2884 61498 2890 61500
rect 2644 61446 2646 61498
rect 2826 61446 2828 61498
rect 2582 61444 2588 61446
rect 2644 61444 2668 61446
rect 2724 61444 2748 61446
rect 2804 61444 2828 61446
rect 2884 61444 2890 61446
rect 2582 61424 2890 61444
rect 2504 61192 2556 61198
rect 2504 61134 2556 61140
rect 2516 60790 2544 61134
rect 2504 60784 2556 60790
rect 2504 60726 2556 60732
rect 2976 60734 3004 63378
rect 3160 63238 3188 66166
rect 3148 63232 3200 63238
rect 3148 63174 3200 63180
rect 2516 54602 2544 60726
rect 2780 60716 2832 60722
rect 2976 60706 3096 60734
rect 2780 60658 2832 60664
rect 2792 60625 2820 60658
rect 2778 60616 2834 60625
rect 2778 60551 2834 60560
rect 2582 60412 2890 60432
rect 2582 60410 2588 60412
rect 2644 60410 2668 60412
rect 2724 60410 2748 60412
rect 2804 60410 2828 60412
rect 2884 60410 2890 60412
rect 2644 60358 2646 60410
rect 2826 60358 2828 60410
rect 2582 60356 2588 60358
rect 2644 60356 2668 60358
rect 2724 60356 2748 60358
rect 2804 60356 2828 60358
rect 2884 60356 2890 60358
rect 2582 60336 2890 60356
rect 2582 59324 2890 59344
rect 2582 59322 2588 59324
rect 2644 59322 2668 59324
rect 2724 59322 2748 59324
rect 2804 59322 2828 59324
rect 2884 59322 2890 59324
rect 2644 59270 2646 59322
rect 2826 59270 2828 59322
rect 2582 59268 2588 59270
rect 2644 59268 2668 59270
rect 2724 59268 2748 59270
rect 2804 59268 2828 59270
rect 2884 59268 2890 59270
rect 2582 59248 2890 59268
rect 2582 58236 2890 58256
rect 2582 58234 2588 58236
rect 2644 58234 2668 58236
rect 2724 58234 2748 58236
rect 2804 58234 2828 58236
rect 2884 58234 2890 58236
rect 2644 58182 2646 58234
rect 2826 58182 2828 58234
rect 2582 58180 2588 58182
rect 2644 58180 2668 58182
rect 2724 58180 2748 58182
rect 2804 58180 2828 58182
rect 2884 58180 2890 58182
rect 2582 58160 2890 58180
rect 2582 57148 2890 57168
rect 2582 57146 2588 57148
rect 2644 57146 2668 57148
rect 2724 57146 2748 57148
rect 2804 57146 2828 57148
rect 2884 57146 2890 57148
rect 2644 57094 2646 57146
rect 2826 57094 2828 57146
rect 2582 57092 2588 57094
rect 2644 57092 2668 57094
rect 2724 57092 2748 57094
rect 2804 57092 2828 57094
rect 2884 57092 2890 57094
rect 2582 57072 2890 57092
rect 2964 56364 3016 56370
rect 2964 56306 3016 56312
rect 2582 56060 2890 56080
rect 2582 56058 2588 56060
rect 2644 56058 2668 56060
rect 2724 56058 2748 56060
rect 2804 56058 2828 56060
rect 2884 56058 2890 56060
rect 2644 56006 2646 56058
rect 2826 56006 2828 56058
rect 2582 56004 2588 56006
rect 2644 56004 2668 56006
rect 2724 56004 2748 56006
rect 2804 56004 2828 56006
rect 2884 56004 2890 56006
rect 2582 55984 2890 56004
rect 2976 55706 3004 56306
rect 3068 55842 3096 60706
rect 3252 56982 3280 68682
rect 3436 66706 3464 69158
rect 3424 66700 3476 66706
rect 3424 66642 3476 66648
rect 3436 63322 3464 66642
rect 3344 63294 3464 63322
rect 3240 56976 3292 56982
rect 3240 56918 3292 56924
rect 3068 55814 3280 55842
rect 2976 55678 3188 55706
rect 2582 54972 2890 54992
rect 2582 54970 2588 54972
rect 2644 54970 2668 54972
rect 2724 54970 2748 54972
rect 2804 54970 2828 54972
rect 2884 54970 2890 54972
rect 2644 54918 2646 54970
rect 2826 54918 2828 54970
rect 2582 54916 2588 54918
rect 2644 54916 2668 54918
rect 2724 54916 2748 54918
rect 2804 54916 2828 54918
rect 2884 54916 2890 54918
rect 2582 54896 2890 54916
rect 2504 54596 2556 54602
rect 2504 54538 2556 54544
rect 2412 54324 2464 54330
rect 2412 54266 2464 54272
rect 2332 54182 2452 54210
rect 2424 54126 2452 54182
rect 2412 54120 2464 54126
rect 2412 54062 2464 54068
rect 2424 52494 2452 54062
rect 3056 53984 3108 53990
rect 3056 53926 3108 53932
rect 2582 53884 2890 53904
rect 2582 53882 2588 53884
rect 2644 53882 2668 53884
rect 2724 53882 2748 53884
rect 2804 53882 2828 53884
rect 2884 53882 2890 53884
rect 2644 53830 2646 53882
rect 2826 53830 2828 53882
rect 2582 53828 2588 53830
rect 2644 53828 2668 53830
rect 2724 53828 2748 53830
rect 2804 53828 2828 53830
rect 2884 53828 2890 53830
rect 2582 53808 2890 53828
rect 2504 53100 2556 53106
rect 2504 53042 2556 53048
rect 2412 52488 2464 52494
rect 2412 52430 2464 52436
rect 2424 51474 2452 52430
rect 2412 51468 2464 51474
rect 2412 51410 2464 51416
rect 2516 51066 2544 53042
rect 2582 52796 2890 52816
rect 2582 52794 2588 52796
rect 2644 52794 2668 52796
rect 2724 52794 2748 52796
rect 2804 52794 2828 52796
rect 2884 52794 2890 52796
rect 2644 52742 2646 52794
rect 2826 52742 2828 52794
rect 2582 52740 2588 52742
rect 2644 52740 2668 52742
rect 2724 52740 2748 52742
rect 2804 52740 2828 52742
rect 2884 52740 2890 52742
rect 2582 52720 2890 52740
rect 2780 52624 2832 52630
rect 2780 52566 2832 52572
rect 2792 52465 2820 52566
rect 2964 52488 3016 52494
rect 2778 52456 2834 52465
rect 2964 52430 3016 52436
rect 2778 52391 2834 52400
rect 2582 51708 2890 51728
rect 2582 51706 2588 51708
rect 2644 51706 2668 51708
rect 2724 51706 2748 51708
rect 2804 51706 2828 51708
rect 2884 51706 2890 51708
rect 2644 51654 2646 51706
rect 2826 51654 2828 51706
rect 2582 51652 2588 51654
rect 2644 51652 2668 51654
rect 2724 51652 2748 51654
rect 2804 51652 2828 51654
rect 2884 51652 2890 51654
rect 2582 51632 2890 51652
rect 2596 51536 2648 51542
rect 2596 51478 2648 51484
rect 2504 51060 2556 51066
rect 2504 51002 2556 51008
rect 2608 50708 2636 51478
rect 2976 51218 3004 52430
rect 3068 51241 3096 53926
rect 2516 50680 2636 50708
rect 2884 51190 3004 51218
rect 3054 51232 3110 51241
rect 2884 50708 2912 51190
rect 3054 51167 3110 51176
rect 3160 51066 3188 55678
rect 3148 51060 3200 51066
rect 3148 51002 3200 51008
rect 3146 50960 3202 50969
rect 3146 50895 3202 50904
rect 2884 50680 3004 50708
rect 2412 49700 2464 49706
rect 2412 49642 2464 49648
rect 2320 49632 2372 49638
rect 2320 49574 2372 49580
rect 2228 47796 2280 47802
rect 2228 47738 2280 47744
rect 2332 45558 2360 49574
rect 2320 45552 2372 45558
rect 2320 45494 2372 45500
rect 2228 45416 2280 45422
rect 2228 45358 2280 45364
rect 2136 41200 2188 41206
rect 2136 41142 2188 41148
rect 2044 40656 2096 40662
rect 2044 40598 2096 40604
rect 2044 40044 2096 40050
rect 2044 39986 2096 39992
rect 1952 38820 2004 38826
rect 1952 38762 2004 38768
rect 2056 35894 2084 39986
rect 2240 39545 2268 45358
rect 2320 44192 2372 44198
rect 2320 44134 2372 44140
rect 2226 39536 2282 39545
rect 2332 39506 2360 44134
rect 2424 41818 2452 49642
rect 2516 48314 2544 50680
rect 2582 50620 2890 50640
rect 2582 50618 2588 50620
rect 2644 50618 2668 50620
rect 2724 50618 2748 50620
rect 2804 50618 2828 50620
rect 2884 50618 2890 50620
rect 2644 50566 2646 50618
rect 2826 50566 2828 50618
rect 2582 50564 2588 50566
rect 2644 50564 2668 50566
rect 2724 50564 2748 50566
rect 2804 50564 2828 50566
rect 2884 50564 2890 50566
rect 2582 50544 2890 50564
rect 2582 49532 2890 49552
rect 2582 49530 2588 49532
rect 2644 49530 2668 49532
rect 2724 49530 2748 49532
rect 2804 49530 2828 49532
rect 2884 49530 2890 49532
rect 2644 49478 2646 49530
rect 2826 49478 2828 49530
rect 2582 49476 2588 49478
rect 2644 49476 2668 49478
rect 2724 49476 2748 49478
rect 2804 49476 2828 49478
rect 2884 49476 2890 49478
rect 2582 49456 2890 49476
rect 2582 48444 2890 48464
rect 2582 48442 2588 48444
rect 2644 48442 2668 48444
rect 2724 48442 2748 48444
rect 2804 48442 2828 48444
rect 2884 48442 2890 48444
rect 2644 48390 2646 48442
rect 2826 48390 2828 48442
rect 2582 48388 2588 48390
rect 2644 48388 2668 48390
rect 2724 48388 2748 48390
rect 2804 48388 2828 48390
rect 2884 48388 2890 48390
rect 2582 48368 2890 48388
rect 2516 48286 2912 48314
rect 2502 47560 2558 47569
rect 2884 47530 2912 48286
rect 2502 47495 2558 47504
rect 2872 47524 2924 47530
rect 2516 44334 2544 47495
rect 2872 47466 2924 47472
rect 2582 47356 2890 47376
rect 2582 47354 2588 47356
rect 2644 47354 2668 47356
rect 2724 47354 2748 47356
rect 2804 47354 2828 47356
rect 2884 47354 2890 47356
rect 2644 47302 2646 47354
rect 2826 47302 2828 47354
rect 2582 47300 2588 47302
rect 2644 47300 2668 47302
rect 2724 47300 2748 47302
rect 2804 47300 2828 47302
rect 2884 47300 2890 47302
rect 2582 47280 2890 47300
rect 2582 46268 2890 46288
rect 2582 46266 2588 46268
rect 2644 46266 2668 46268
rect 2724 46266 2748 46268
rect 2804 46266 2828 46268
rect 2884 46266 2890 46268
rect 2644 46214 2646 46266
rect 2826 46214 2828 46266
rect 2582 46212 2588 46214
rect 2644 46212 2668 46214
rect 2724 46212 2748 46214
rect 2804 46212 2828 46214
rect 2884 46212 2890 46214
rect 2582 46192 2890 46212
rect 2582 45180 2890 45200
rect 2582 45178 2588 45180
rect 2644 45178 2668 45180
rect 2724 45178 2748 45180
rect 2804 45178 2828 45180
rect 2884 45178 2890 45180
rect 2644 45126 2646 45178
rect 2826 45126 2828 45178
rect 2582 45124 2588 45126
rect 2644 45124 2668 45126
rect 2724 45124 2748 45126
rect 2804 45124 2828 45126
rect 2884 45124 2890 45126
rect 2582 45104 2890 45124
rect 2504 44328 2556 44334
rect 2504 44270 2556 44276
rect 2582 44092 2890 44112
rect 2582 44090 2588 44092
rect 2644 44090 2668 44092
rect 2724 44090 2748 44092
rect 2804 44090 2828 44092
rect 2884 44090 2890 44092
rect 2644 44038 2646 44090
rect 2826 44038 2828 44090
rect 2582 44036 2588 44038
rect 2644 44036 2668 44038
rect 2724 44036 2748 44038
rect 2804 44036 2828 44038
rect 2884 44036 2890 44038
rect 2582 44016 2890 44036
rect 2504 43920 2556 43926
rect 2504 43862 2556 43868
rect 2412 41812 2464 41818
rect 2412 41754 2464 41760
rect 2516 41414 2544 43862
rect 2582 43004 2890 43024
rect 2582 43002 2588 43004
rect 2644 43002 2668 43004
rect 2724 43002 2748 43004
rect 2804 43002 2828 43004
rect 2884 43002 2890 43004
rect 2644 42950 2646 43002
rect 2826 42950 2828 43002
rect 2582 42948 2588 42950
rect 2644 42948 2668 42950
rect 2724 42948 2748 42950
rect 2804 42948 2828 42950
rect 2884 42948 2890 42950
rect 2582 42928 2890 42948
rect 2582 41916 2890 41936
rect 2582 41914 2588 41916
rect 2644 41914 2668 41916
rect 2724 41914 2748 41916
rect 2804 41914 2828 41916
rect 2884 41914 2890 41916
rect 2644 41862 2646 41914
rect 2826 41862 2828 41914
rect 2582 41860 2588 41862
rect 2644 41860 2668 41862
rect 2724 41860 2748 41862
rect 2804 41860 2828 41862
rect 2884 41860 2890 41862
rect 2582 41840 2890 41860
rect 2424 41386 2544 41414
rect 2226 39471 2282 39480
rect 2320 39500 2372 39506
rect 2320 39442 2372 39448
rect 2228 39296 2280 39302
rect 2228 39238 2280 39244
rect 2240 37262 2268 39238
rect 2228 37256 2280 37262
rect 2228 37198 2280 37204
rect 1964 35866 2084 35894
rect 1964 29170 1992 35866
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 2056 32570 2084 35022
rect 2240 33114 2268 37198
rect 2332 37126 2360 39442
rect 2320 37120 2372 37126
rect 2320 37062 2372 37068
rect 2424 36938 2452 41386
rect 2504 41268 2556 41274
rect 2504 41210 2556 41216
rect 2516 39642 2544 41210
rect 2582 40828 2890 40848
rect 2582 40826 2588 40828
rect 2644 40826 2668 40828
rect 2724 40826 2748 40828
rect 2804 40826 2828 40828
rect 2884 40826 2890 40828
rect 2644 40774 2646 40826
rect 2826 40774 2828 40826
rect 2582 40772 2588 40774
rect 2644 40772 2668 40774
rect 2724 40772 2748 40774
rect 2804 40772 2828 40774
rect 2884 40772 2890 40774
rect 2582 40752 2890 40772
rect 2582 39740 2890 39760
rect 2582 39738 2588 39740
rect 2644 39738 2668 39740
rect 2724 39738 2748 39740
rect 2804 39738 2828 39740
rect 2884 39738 2890 39740
rect 2644 39686 2646 39738
rect 2826 39686 2828 39738
rect 2582 39684 2588 39686
rect 2644 39684 2668 39686
rect 2724 39684 2748 39686
rect 2804 39684 2828 39686
rect 2884 39684 2890 39686
rect 2582 39664 2890 39684
rect 2504 39636 2556 39642
rect 2504 39578 2556 39584
rect 2504 39364 2556 39370
rect 2504 39306 2556 39312
rect 2516 37330 2544 39306
rect 2582 38652 2890 38672
rect 2582 38650 2588 38652
rect 2644 38650 2668 38652
rect 2724 38650 2748 38652
rect 2804 38650 2828 38652
rect 2884 38650 2890 38652
rect 2644 38598 2646 38650
rect 2826 38598 2828 38650
rect 2582 38596 2588 38598
rect 2644 38596 2668 38598
rect 2724 38596 2748 38598
rect 2804 38596 2828 38598
rect 2884 38596 2890 38598
rect 2582 38576 2890 38596
rect 2686 37768 2742 37777
rect 2686 37703 2688 37712
rect 2740 37703 2742 37712
rect 2688 37674 2740 37680
rect 2582 37564 2890 37584
rect 2582 37562 2588 37564
rect 2644 37562 2668 37564
rect 2724 37562 2748 37564
rect 2804 37562 2828 37564
rect 2884 37562 2890 37564
rect 2644 37510 2646 37562
rect 2826 37510 2828 37562
rect 2582 37508 2588 37510
rect 2644 37508 2668 37510
rect 2724 37508 2748 37510
rect 2804 37508 2828 37510
rect 2884 37508 2890 37510
rect 2582 37488 2890 37508
rect 2504 37324 2556 37330
rect 2504 37266 2556 37272
rect 2332 36910 2452 36938
rect 2332 36242 2360 36910
rect 2516 36242 2544 37266
rect 2582 36476 2890 36496
rect 2582 36474 2588 36476
rect 2644 36474 2668 36476
rect 2724 36474 2748 36476
rect 2804 36474 2828 36476
rect 2884 36474 2890 36476
rect 2644 36422 2646 36474
rect 2826 36422 2828 36474
rect 2582 36420 2588 36422
rect 2644 36420 2668 36422
rect 2724 36420 2748 36422
rect 2804 36420 2828 36422
rect 2884 36420 2890 36422
rect 2582 36400 2890 36420
rect 2320 36236 2372 36242
rect 2320 36178 2372 36184
rect 2504 36236 2556 36242
rect 2504 36178 2556 36184
rect 2332 35154 2360 36178
rect 2412 36168 2464 36174
rect 2412 36110 2464 36116
rect 2320 35148 2372 35154
rect 2320 35090 2372 35096
rect 2424 35086 2452 36110
rect 2516 35136 2544 36178
rect 2582 35388 2890 35408
rect 2582 35386 2588 35388
rect 2644 35386 2668 35388
rect 2724 35386 2748 35388
rect 2804 35386 2828 35388
rect 2884 35386 2890 35388
rect 2644 35334 2646 35386
rect 2826 35334 2828 35386
rect 2582 35332 2588 35334
rect 2644 35332 2668 35334
rect 2724 35332 2748 35334
rect 2804 35332 2828 35334
rect 2884 35332 2890 35334
rect 2582 35312 2890 35332
rect 2596 35148 2648 35154
rect 2516 35108 2596 35136
rect 2596 35090 2648 35096
rect 2412 35080 2464 35086
rect 2412 35022 2464 35028
rect 2424 34610 2544 34626
rect 2608 34610 2636 35090
rect 2424 34604 2556 34610
rect 2424 34598 2504 34604
rect 2320 34536 2372 34542
rect 2320 34478 2372 34484
rect 2228 33108 2280 33114
rect 2228 33050 2280 33056
rect 2332 32910 2360 34478
rect 2320 32904 2372 32910
rect 2320 32846 2372 32852
rect 2424 32858 2452 34598
rect 2504 34546 2556 34552
rect 2596 34604 2648 34610
rect 2596 34546 2648 34552
rect 2608 34456 2636 34546
rect 2516 34428 2636 34456
rect 2516 32978 2544 34428
rect 2582 34300 2890 34320
rect 2582 34298 2588 34300
rect 2644 34298 2668 34300
rect 2724 34298 2748 34300
rect 2804 34298 2828 34300
rect 2884 34298 2890 34300
rect 2644 34246 2646 34298
rect 2826 34246 2828 34298
rect 2582 34244 2588 34246
rect 2644 34244 2668 34246
rect 2724 34244 2748 34246
rect 2804 34244 2828 34246
rect 2884 34244 2890 34246
rect 2582 34224 2890 34244
rect 2582 33212 2890 33232
rect 2582 33210 2588 33212
rect 2644 33210 2668 33212
rect 2724 33210 2748 33212
rect 2804 33210 2828 33212
rect 2884 33210 2890 33212
rect 2644 33158 2646 33210
rect 2826 33158 2828 33210
rect 2582 33156 2588 33158
rect 2644 33156 2668 33158
rect 2724 33156 2748 33158
rect 2804 33156 2828 33158
rect 2884 33156 2890 33158
rect 2582 33136 2890 33156
rect 2504 32972 2556 32978
rect 2504 32914 2556 32920
rect 2424 32830 2544 32858
rect 2516 32774 2544 32830
rect 2136 32768 2188 32774
rect 2136 32710 2188 32716
rect 2504 32768 2556 32774
rect 2504 32710 2556 32716
rect 2148 32570 2176 32710
rect 2044 32564 2096 32570
rect 2044 32506 2096 32512
rect 2136 32564 2188 32570
rect 2136 32506 2188 32512
rect 2516 32026 2544 32710
rect 2582 32124 2890 32144
rect 2582 32122 2588 32124
rect 2644 32122 2668 32124
rect 2724 32122 2748 32124
rect 2804 32122 2828 32124
rect 2884 32122 2890 32124
rect 2644 32070 2646 32122
rect 2826 32070 2828 32122
rect 2582 32068 2588 32070
rect 2644 32068 2668 32070
rect 2724 32068 2748 32070
rect 2804 32068 2828 32070
rect 2884 32068 2890 32070
rect 2582 32048 2890 32068
rect 2504 32020 2556 32026
rect 2504 31962 2556 31968
rect 2582 31036 2890 31056
rect 2582 31034 2588 31036
rect 2644 31034 2668 31036
rect 2724 31034 2748 31036
rect 2804 31034 2828 31036
rect 2884 31034 2890 31036
rect 2644 30982 2646 31034
rect 2826 30982 2828 31034
rect 2582 30980 2588 30982
rect 2644 30980 2668 30982
rect 2724 30980 2748 30982
rect 2804 30980 2828 30982
rect 2884 30980 2890 30982
rect 2582 30960 2890 30980
rect 2582 29948 2890 29968
rect 2582 29946 2588 29948
rect 2644 29946 2668 29948
rect 2724 29946 2748 29948
rect 2804 29946 2828 29948
rect 2884 29946 2890 29948
rect 2644 29894 2646 29946
rect 2826 29894 2828 29946
rect 2582 29892 2588 29894
rect 2644 29892 2668 29894
rect 2724 29892 2748 29894
rect 2804 29892 2828 29894
rect 2884 29892 2890 29894
rect 2582 29872 2890 29892
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 2582 28860 2890 28880
rect 2582 28858 2588 28860
rect 2644 28858 2668 28860
rect 2724 28858 2748 28860
rect 2804 28858 2828 28860
rect 2884 28858 2890 28860
rect 2644 28806 2646 28858
rect 2826 28806 2828 28858
rect 2582 28804 2588 28806
rect 2644 28804 2668 28806
rect 2724 28804 2748 28806
rect 2804 28804 2828 28806
rect 2884 28804 2890 28806
rect 2582 28784 2890 28804
rect 2582 27772 2890 27792
rect 2582 27770 2588 27772
rect 2644 27770 2668 27772
rect 2724 27770 2748 27772
rect 2804 27770 2828 27772
rect 2884 27770 2890 27772
rect 2644 27718 2646 27770
rect 2826 27718 2828 27770
rect 2582 27716 2588 27718
rect 2644 27716 2668 27718
rect 2724 27716 2748 27718
rect 2804 27716 2828 27718
rect 2884 27716 2890 27718
rect 2582 27696 2890 27716
rect 2582 26684 2890 26704
rect 2582 26682 2588 26684
rect 2644 26682 2668 26684
rect 2724 26682 2748 26684
rect 2804 26682 2828 26684
rect 2884 26682 2890 26684
rect 2644 26630 2646 26682
rect 2826 26630 2828 26682
rect 2582 26628 2588 26630
rect 2644 26628 2668 26630
rect 2724 26628 2748 26630
rect 2804 26628 2828 26630
rect 2884 26628 2890 26630
rect 2582 26608 2890 26628
rect 2582 25596 2890 25616
rect 2582 25594 2588 25596
rect 2644 25594 2668 25596
rect 2724 25594 2748 25596
rect 2804 25594 2828 25596
rect 2884 25594 2890 25596
rect 2644 25542 2646 25594
rect 2826 25542 2828 25594
rect 2582 25540 2588 25542
rect 2644 25540 2668 25542
rect 2724 25540 2748 25542
rect 2804 25540 2828 25542
rect 2884 25540 2890 25542
rect 2582 25520 2890 25540
rect 2582 24508 2890 24528
rect 2582 24506 2588 24508
rect 2644 24506 2668 24508
rect 2724 24506 2748 24508
rect 2804 24506 2828 24508
rect 2884 24506 2890 24508
rect 2644 24454 2646 24506
rect 2826 24454 2828 24506
rect 2582 24452 2588 24454
rect 2644 24452 2668 24454
rect 2724 24452 2748 24454
rect 2804 24452 2828 24454
rect 2884 24452 2890 24454
rect 2582 24432 2890 24452
rect 2582 23420 2890 23440
rect 2582 23418 2588 23420
rect 2644 23418 2668 23420
rect 2724 23418 2748 23420
rect 2804 23418 2828 23420
rect 2884 23418 2890 23420
rect 2644 23366 2646 23418
rect 2826 23366 2828 23418
rect 2582 23364 2588 23366
rect 2644 23364 2668 23366
rect 2724 23364 2748 23366
rect 2804 23364 2828 23366
rect 2884 23364 2890 23366
rect 2582 23344 2890 23364
rect 2582 22332 2890 22352
rect 2582 22330 2588 22332
rect 2644 22330 2668 22332
rect 2724 22330 2748 22332
rect 2804 22330 2828 22332
rect 2884 22330 2890 22332
rect 2644 22278 2646 22330
rect 2826 22278 2828 22330
rect 2582 22276 2588 22278
rect 2644 22276 2668 22278
rect 2724 22276 2748 22278
rect 2804 22276 2828 22278
rect 2884 22276 2890 22278
rect 2582 22256 2890 22276
rect 2582 21244 2890 21264
rect 2582 21242 2588 21244
rect 2644 21242 2668 21244
rect 2724 21242 2748 21244
rect 2804 21242 2828 21244
rect 2884 21242 2890 21244
rect 2644 21190 2646 21242
rect 2826 21190 2828 21242
rect 2582 21188 2588 21190
rect 2644 21188 2668 21190
rect 2724 21188 2748 21190
rect 2804 21188 2828 21190
rect 2884 21188 2890 21190
rect 2582 21168 2890 21188
rect 2582 20156 2890 20176
rect 2582 20154 2588 20156
rect 2644 20154 2668 20156
rect 2724 20154 2748 20156
rect 2804 20154 2828 20156
rect 2884 20154 2890 20156
rect 2644 20102 2646 20154
rect 2826 20102 2828 20154
rect 2582 20100 2588 20102
rect 2644 20100 2668 20102
rect 2724 20100 2748 20102
rect 2804 20100 2828 20102
rect 2884 20100 2890 20102
rect 2582 20080 2890 20100
rect 2582 19068 2890 19088
rect 2582 19066 2588 19068
rect 2644 19066 2668 19068
rect 2724 19066 2748 19068
rect 2804 19066 2828 19068
rect 2884 19066 2890 19068
rect 2644 19014 2646 19066
rect 2826 19014 2828 19066
rect 2582 19012 2588 19014
rect 2644 19012 2668 19014
rect 2724 19012 2748 19014
rect 2804 19012 2828 19014
rect 2884 19012 2890 19014
rect 2582 18992 2890 19012
rect 2582 17980 2890 18000
rect 2582 17978 2588 17980
rect 2644 17978 2668 17980
rect 2724 17978 2748 17980
rect 2804 17978 2828 17980
rect 2884 17978 2890 17980
rect 2644 17926 2646 17978
rect 2826 17926 2828 17978
rect 2582 17924 2588 17926
rect 2644 17924 2668 17926
rect 2724 17924 2748 17926
rect 2804 17924 2828 17926
rect 2884 17924 2890 17926
rect 2582 17904 2890 17924
rect 2976 17678 3004 50680
rect 3056 50244 3108 50250
rect 3056 50186 3108 50192
rect 3068 36242 3096 50186
rect 3056 36236 3108 36242
rect 3056 36178 3108 36184
rect 3160 34678 3188 50895
rect 3252 44470 3280 55814
rect 3344 45014 3372 63294
rect 3528 63186 3556 69770
rect 3792 69352 3844 69358
rect 3792 69294 3844 69300
rect 3608 66700 3660 66706
rect 3608 66642 3660 66648
rect 3620 66094 3648 66642
rect 3608 66088 3660 66094
rect 3608 66030 3660 66036
rect 3620 63442 3648 66030
rect 3608 63436 3660 63442
rect 3608 63378 3660 63384
rect 3436 63158 3556 63186
rect 3332 45008 3384 45014
rect 3332 44950 3384 44956
rect 3332 44872 3384 44878
rect 3332 44814 3384 44820
rect 3240 44464 3292 44470
rect 3240 44406 3292 44412
rect 3240 42220 3292 42226
rect 3344 42208 3372 44814
rect 3292 42180 3372 42208
rect 3240 42162 3292 42168
rect 3252 39506 3280 42162
rect 3332 41540 3384 41546
rect 3332 41482 3384 41488
rect 3344 40050 3372 41482
rect 3332 40044 3384 40050
rect 3332 39986 3384 39992
rect 3240 39500 3292 39506
rect 3240 39442 3292 39448
rect 3436 36854 3464 63158
rect 3516 62212 3568 62218
rect 3516 62154 3568 62160
rect 3528 42566 3556 62154
rect 3608 61668 3660 61674
rect 3608 61610 3660 61616
rect 3620 58682 3648 61610
rect 3608 58676 3660 58682
rect 3608 58618 3660 58624
rect 3804 57974 3832 69294
rect 3896 68474 3924 70790
rect 3976 69896 4028 69902
rect 3976 69838 4028 69844
rect 3988 69737 4016 69838
rect 3974 69728 4030 69737
rect 3974 69663 4030 69672
rect 3884 68468 3936 68474
rect 3884 68410 3936 68416
rect 3976 60580 4028 60586
rect 3976 60522 4028 60528
rect 3884 58676 3936 58682
rect 3884 58618 3936 58624
rect 3712 57946 3832 57974
rect 3608 56976 3660 56982
rect 3608 56918 3660 56924
rect 3620 50969 3648 56918
rect 3606 50960 3662 50969
rect 3606 50895 3662 50904
rect 3608 50856 3660 50862
rect 3608 50798 3660 50804
rect 3620 49774 3648 50798
rect 3608 49768 3660 49774
rect 3712 49745 3740 57946
rect 3792 56840 3844 56846
rect 3792 56782 3844 56788
rect 3608 49710 3660 49716
rect 3698 49736 3754 49745
rect 3698 49671 3754 49680
rect 3804 49609 3832 56782
rect 3606 49600 3662 49609
rect 3606 49535 3662 49544
rect 3790 49600 3846 49609
rect 3790 49535 3846 49544
rect 3620 47734 3648 49535
rect 3698 49464 3754 49473
rect 3698 49399 3754 49408
rect 3792 49428 3844 49434
rect 3608 47728 3660 47734
rect 3608 47670 3660 47676
rect 3608 47524 3660 47530
rect 3608 47466 3660 47472
rect 3620 43382 3648 47466
rect 3608 43376 3660 43382
rect 3608 43318 3660 43324
rect 3608 42696 3660 42702
rect 3608 42638 3660 42644
rect 3516 42560 3568 42566
rect 3516 42502 3568 42508
rect 3516 41676 3568 41682
rect 3516 41618 3568 41624
rect 3424 36848 3476 36854
rect 3424 36790 3476 36796
rect 3148 34672 3200 34678
rect 3148 34614 3200 34620
rect 3424 33652 3476 33658
rect 3424 33594 3476 33600
rect 3436 23730 3464 33594
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3528 21690 3556 41618
rect 3620 26382 3648 42638
rect 3712 38962 3740 49399
rect 3792 49370 3844 49376
rect 3804 45506 3832 49370
rect 3896 45626 3924 58618
rect 3884 45620 3936 45626
rect 3884 45562 3936 45568
rect 3804 45478 3924 45506
rect 3790 45384 3846 45393
rect 3790 45319 3846 45328
rect 3804 41614 3832 45319
rect 3792 41608 3844 41614
rect 3792 41550 3844 41556
rect 3792 41472 3844 41478
rect 3792 41414 3844 41420
rect 3700 38956 3752 38962
rect 3700 38898 3752 38904
rect 3608 26376 3660 26382
rect 3608 26318 3660 26324
rect 3804 22778 3832 41414
rect 3896 40118 3924 45478
rect 3988 44198 4016 60522
rect 4080 49366 4108 72014
rect 4213 71836 4521 71856
rect 4213 71834 4219 71836
rect 4275 71834 4299 71836
rect 4355 71834 4379 71836
rect 4435 71834 4459 71836
rect 4515 71834 4521 71836
rect 4275 71782 4277 71834
rect 4457 71782 4459 71834
rect 4213 71780 4219 71782
rect 4275 71780 4299 71782
rect 4355 71780 4379 71782
rect 4435 71780 4459 71782
rect 4515 71780 4521 71782
rect 4213 71760 4521 71780
rect 4632 70990 4660 74598
rect 5845 74556 6153 74576
rect 5845 74554 5851 74556
rect 5907 74554 5931 74556
rect 5987 74554 6011 74556
rect 6067 74554 6091 74556
rect 6147 74554 6153 74556
rect 5907 74502 5909 74554
rect 6089 74502 6091 74554
rect 5845 74500 5851 74502
rect 5907 74500 5931 74502
rect 5987 74500 6011 74502
rect 6067 74500 6091 74502
rect 6147 74500 6153 74502
rect 5845 74480 6153 74500
rect 6196 74458 6224 77454
rect 7477 77276 7785 77296
rect 7477 77274 7483 77276
rect 7539 77274 7563 77276
rect 7619 77274 7643 77276
rect 7699 77274 7723 77276
rect 7779 77274 7785 77276
rect 7539 77222 7541 77274
rect 7721 77222 7723 77274
rect 7477 77220 7483 77222
rect 7539 77220 7563 77222
rect 7619 77220 7643 77222
rect 7699 77220 7723 77222
rect 7779 77220 7785 77222
rect 7477 77200 7785 77220
rect 8588 77178 8616 79183
rect 9494 78704 9550 78713
rect 9494 78639 9550 78648
rect 9109 77820 9417 77840
rect 9109 77818 9115 77820
rect 9171 77818 9195 77820
rect 9251 77818 9275 77820
rect 9331 77818 9355 77820
rect 9411 77818 9417 77820
rect 9171 77766 9173 77818
rect 9353 77766 9355 77818
rect 9109 77764 9115 77766
rect 9171 77764 9195 77766
rect 9251 77764 9275 77766
rect 9331 77764 9355 77766
rect 9411 77764 9417 77766
rect 9109 77744 9417 77764
rect 8944 77512 8996 77518
rect 8944 77454 8996 77460
rect 8576 77172 8628 77178
rect 8576 77114 8628 77120
rect 8392 77036 8444 77042
rect 8392 76978 8444 76984
rect 6460 76832 6512 76838
rect 6460 76774 6512 76780
rect 6184 74452 6236 74458
rect 6184 74394 6236 74400
rect 6472 74186 6500 76774
rect 8300 76424 8352 76430
rect 8300 76366 8352 76372
rect 7477 76188 7785 76208
rect 7477 76186 7483 76188
rect 7539 76186 7563 76188
rect 7619 76186 7643 76188
rect 7699 76186 7723 76188
rect 7779 76186 7785 76188
rect 7539 76134 7541 76186
rect 7721 76134 7723 76186
rect 7477 76132 7483 76134
rect 7539 76132 7563 76134
rect 7619 76132 7643 76134
rect 7699 76132 7723 76134
rect 7779 76132 7785 76134
rect 7477 76112 7785 76132
rect 7477 75100 7785 75120
rect 7477 75098 7483 75100
rect 7539 75098 7563 75100
rect 7619 75098 7643 75100
rect 7699 75098 7723 75100
rect 7779 75098 7785 75100
rect 7539 75046 7541 75098
rect 7721 75046 7723 75098
rect 7477 75044 7483 75046
rect 7539 75044 7563 75046
rect 7619 75044 7643 75046
rect 7699 75044 7723 75046
rect 7779 75044 7785 75046
rect 7477 75024 7785 75044
rect 6828 74316 6880 74322
rect 6828 74258 6880 74264
rect 6460 74180 6512 74186
rect 6460 74122 6512 74128
rect 6644 74180 6696 74186
rect 6644 74122 6696 74128
rect 6368 74112 6420 74118
rect 6368 74054 6420 74060
rect 5845 73468 6153 73488
rect 5845 73466 5851 73468
rect 5907 73466 5931 73468
rect 5987 73466 6011 73468
rect 6067 73466 6091 73468
rect 6147 73466 6153 73468
rect 5907 73414 5909 73466
rect 6089 73414 6091 73466
rect 5845 73412 5851 73414
rect 5907 73412 5931 73414
rect 5987 73412 6011 73414
rect 6067 73412 6091 73414
rect 6147 73412 6153 73414
rect 5845 73392 6153 73412
rect 5845 72380 6153 72400
rect 5845 72378 5851 72380
rect 5907 72378 5931 72380
rect 5987 72378 6011 72380
rect 6067 72378 6091 72380
rect 6147 72378 6153 72380
rect 5907 72326 5909 72378
rect 6089 72326 6091 72378
rect 5845 72324 5851 72326
rect 5907 72324 5931 72326
rect 5987 72324 6011 72326
rect 6067 72324 6091 72326
rect 6147 72324 6153 72326
rect 5845 72304 6153 72324
rect 6184 72208 6236 72214
rect 6184 72150 6236 72156
rect 4804 72004 4856 72010
rect 4804 71946 4856 71952
rect 5724 72004 5776 72010
rect 5724 71946 5776 71952
rect 4620 70984 4672 70990
rect 4620 70926 4672 70932
rect 4213 70748 4521 70768
rect 4213 70746 4219 70748
rect 4275 70746 4299 70748
rect 4355 70746 4379 70748
rect 4435 70746 4459 70748
rect 4515 70746 4521 70748
rect 4275 70694 4277 70746
rect 4457 70694 4459 70746
rect 4213 70692 4219 70694
rect 4275 70692 4299 70694
rect 4355 70692 4379 70694
rect 4435 70692 4459 70694
rect 4515 70692 4521 70694
rect 4213 70672 4521 70692
rect 4213 69660 4521 69680
rect 4213 69658 4219 69660
rect 4275 69658 4299 69660
rect 4355 69658 4379 69660
rect 4435 69658 4459 69660
rect 4515 69658 4521 69660
rect 4275 69606 4277 69658
rect 4457 69606 4459 69658
rect 4213 69604 4219 69606
rect 4275 69604 4299 69606
rect 4355 69604 4379 69606
rect 4435 69604 4459 69606
rect 4515 69604 4521 69606
rect 4213 69584 4521 69604
rect 4213 68572 4521 68592
rect 4213 68570 4219 68572
rect 4275 68570 4299 68572
rect 4355 68570 4379 68572
rect 4435 68570 4459 68572
rect 4515 68570 4521 68572
rect 4275 68518 4277 68570
rect 4457 68518 4459 68570
rect 4213 68516 4219 68518
rect 4275 68516 4299 68518
rect 4355 68516 4379 68518
rect 4435 68516 4459 68518
rect 4515 68516 4521 68518
rect 4213 68496 4521 68516
rect 4632 68406 4660 70926
rect 4620 68400 4672 68406
rect 4620 68342 4672 68348
rect 4620 68264 4672 68270
rect 4620 68206 4672 68212
rect 4213 67484 4521 67504
rect 4213 67482 4219 67484
rect 4275 67482 4299 67484
rect 4355 67482 4379 67484
rect 4435 67482 4459 67484
rect 4515 67482 4521 67484
rect 4275 67430 4277 67482
rect 4457 67430 4459 67482
rect 4213 67428 4219 67430
rect 4275 67428 4299 67430
rect 4355 67428 4379 67430
rect 4435 67428 4459 67430
rect 4515 67428 4521 67430
rect 4213 67408 4521 67428
rect 4213 66396 4521 66416
rect 4213 66394 4219 66396
rect 4275 66394 4299 66396
rect 4355 66394 4379 66396
rect 4435 66394 4459 66396
rect 4515 66394 4521 66396
rect 4275 66342 4277 66394
rect 4457 66342 4459 66394
rect 4213 66340 4219 66342
rect 4275 66340 4299 66342
rect 4355 66340 4379 66342
rect 4435 66340 4459 66342
rect 4515 66340 4521 66342
rect 4213 66320 4521 66340
rect 4213 65308 4521 65328
rect 4213 65306 4219 65308
rect 4275 65306 4299 65308
rect 4355 65306 4379 65308
rect 4435 65306 4459 65308
rect 4515 65306 4521 65308
rect 4275 65254 4277 65306
rect 4457 65254 4459 65306
rect 4213 65252 4219 65254
rect 4275 65252 4299 65254
rect 4355 65252 4379 65254
rect 4435 65252 4459 65254
rect 4515 65252 4521 65254
rect 4213 65232 4521 65252
rect 4213 64220 4521 64240
rect 4213 64218 4219 64220
rect 4275 64218 4299 64220
rect 4355 64218 4379 64220
rect 4435 64218 4459 64220
rect 4515 64218 4521 64220
rect 4275 64166 4277 64218
rect 4457 64166 4459 64218
rect 4213 64164 4219 64166
rect 4275 64164 4299 64166
rect 4355 64164 4379 64166
rect 4435 64164 4459 64166
rect 4515 64164 4521 64166
rect 4213 64144 4521 64164
rect 4213 63132 4521 63152
rect 4213 63130 4219 63132
rect 4275 63130 4299 63132
rect 4355 63130 4379 63132
rect 4435 63130 4459 63132
rect 4515 63130 4521 63132
rect 4275 63078 4277 63130
rect 4457 63078 4459 63130
rect 4213 63076 4219 63078
rect 4275 63076 4299 63078
rect 4355 63076 4379 63078
rect 4435 63076 4459 63078
rect 4515 63076 4521 63078
rect 4213 63056 4521 63076
rect 4213 62044 4521 62064
rect 4213 62042 4219 62044
rect 4275 62042 4299 62044
rect 4355 62042 4379 62044
rect 4435 62042 4459 62044
rect 4515 62042 4521 62044
rect 4275 61990 4277 62042
rect 4457 61990 4459 62042
rect 4213 61988 4219 61990
rect 4275 61988 4299 61990
rect 4355 61988 4379 61990
rect 4435 61988 4459 61990
rect 4515 61988 4521 61990
rect 4213 61968 4521 61988
rect 4213 60956 4521 60976
rect 4213 60954 4219 60956
rect 4275 60954 4299 60956
rect 4355 60954 4379 60956
rect 4435 60954 4459 60956
rect 4515 60954 4521 60956
rect 4275 60902 4277 60954
rect 4457 60902 4459 60954
rect 4213 60900 4219 60902
rect 4275 60900 4299 60902
rect 4355 60900 4379 60902
rect 4435 60900 4459 60902
rect 4515 60900 4521 60902
rect 4213 60880 4521 60900
rect 4213 59868 4521 59888
rect 4213 59866 4219 59868
rect 4275 59866 4299 59868
rect 4355 59866 4379 59868
rect 4435 59866 4459 59868
rect 4515 59866 4521 59868
rect 4275 59814 4277 59866
rect 4457 59814 4459 59866
rect 4213 59812 4219 59814
rect 4275 59812 4299 59814
rect 4355 59812 4379 59814
rect 4435 59812 4459 59814
rect 4515 59812 4521 59814
rect 4213 59792 4521 59812
rect 4213 58780 4521 58800
rect 4213 58778 4219 58780
rect 4275 58778 4299 58780
rect 4355 58778 4379 58780
rect 4435 58778 4459 58780
rect 4515 58778 4521 58780
rect 4275 58726 4277 58778
rect 4457 58726 4459 58778
rect 4213 58724 4219 58726
rect 4275 58724 4299 58726
rect 4355 58724 4379 58726
rect 4435 58724 4459 58726
rect 4515 58724 4521 58726
rect 4213 58704 4521 58724
rect 4213 57692 4521 57712
rect 4213 57690 4219 57692
rect 4275 57690 4299 57692
rect 4355 57690 4379 57692
rect 4435 57690 4459 57692
rect 4515 57690 4521 57692
rect 4275 57638 4277 57690
rect 4457 57638 4459 57690
rect 4213 57636 4219 57638
rect 4275 57636 4299 57638
rect 4355 57636 4379 57638
rect 4435 57636 4459 57638
rect 4515 57636 4521 57638
rect 4213 57616 4521 57636
rect 4213 56604 4521 56624
rect 4213 56602 4219 56604
rect 4275 56602 4299 56604
rect 4355 56602 4379 56604
rect 4435 56602 4459 56604
rect 4515 56602 4521 56604
rect 4275 56550 4277 56602
rect 4457 56550 4459 56602
rect 4213 56548 4219 56550
rect 4275 56548 4299 56550
rect 4355 56548 4379 56550
rect 4435 56548 4459 56550
rect 4515 56548 4521 56550
rect 4213 56528 4521 56548
rect 4213 55516 4521 55536
rect 4213 55514 4219 55516
rect 4275 55514 4299 55516
rect 4355 55514 4379 55516
rect 4435 55514 4459 55516
rect 4515 55514 4521 55516
rect 4275 55462 4277 55514
rect 4457 55462 4459 55514
rect 4213 55460 4219 55462
rect 4275 55460 4299 55462
rect 4355 55460 4379 55462
rect 4435 55460 4459 55462
rect 4515 55460 4521 55462
rect 4213 55440 4521 55460
rect 4213 54428 4521 54448
rect 4213 54426 4219 54428
rect 4275 54426 4299 54428
rect 4355 54426 4379 54428
rect 4435 54426 4459 54428
rect 4515 54426 4521 54428
rect 4275 54374 4277 54426
rect 4457 54374 4459 54426
rect 4213 54372 4219 54374
rect 4275 54372 4299 54374
rect 4355 54372 4379 54374
rect 4435 54372 4459 54374
rect 4515 54372 4521 54374
rect 4213 54352 4521 54372
rect 4213 53340 4521 53360
rect 4213 53338 4219 53340
rect 4275 53338 4299 53340
rect 4355 53338 4379 53340
rect 4435 53338 4459 53340
rect 4515 53338 4521 53340
rect 4275 53286 4277 53338
rect 4457 53286 4459 53338
rect 4213 53284 4219 53286
rect 4275 53284 4299 53286
rect 4355 53284 4379 53286
rect 4435 53284 4459 53286
rect 4515 53284 4521 53286
rect 4213 53264 4521 53284
rect 4213 52252 4521 52272
rect 4213 52250 4219 52252
rect 4275 52250 4299 52252
rect 4355 52250 4379 52252
rect 4435 52250 4459 52252
rect 4515 52250 4521 52252
rect 4275 52198 4277 52250
rect 4457 52198 4459 52250
rect 4213 52196 4219 52198
rect 4275 52196 4299 52198
rect 4355 52196 4379 52198
rect 4435 52196 4459 52198
rect 4515 52196 4521 52198
rect 4213 52176 4521 52196
rect 4213 51164 4521 51184
rect 4213 51162 4219 51164
rect 4275 51162 4299 51164
rect 4355 51162 4379 51164
rect 4435 51162 4459 51164
rect 4515 51162 4521 51164
rect 4275 51110 4277 51162
rect 4457 51110 4459 51162
rect 4213 51108 4219 51110
rect 4275 51108 4299 51110
rect 4355 51108 4379 51110
rect 4435 51108 4459 51110
rect 4515 51108 4521 51110
rect 4213 51088 4521 51108
rect 4213 50076 4521 50096
rect 4213 50074 4219 50076
rect 4275 50074 4299 50076
rect 4355 50074 4379 50076
rect 4435 50074 4459 50076
rect 4515 50074 4521 50076
rect 4275 50022 4277 50074
rect 4457 50022 4459 50074
rect 4213 50020 4219 50022
rect 4275 50020 4299 50022
rect 4355 50020 4379 50022
rect 4435 50020 4459 50022
rect 4515 50020 4521 50022
rect 4213 50000 4521 50020
rect 4160 49768 4212 49774
rect 4160 49710 4212 49716
rect 4068 49360 4120 49366
rect 4068 49302 4120 49308
rect 4172 49178 4200 49710
rect 4080 49150 4200 49178
rect 4080 47258 4108 49150
rect 4213 48988 4521 49008
rect 4213 48986 4219 48988
rect 4275 48986 4299 48988
rect 4355 48986 4379 48988
rect 4435 48986 4459 48988
rect 4515 48986 4521 48988
rect 4275 48934 4277 48986
rect 4457 48934 4459 48986
rect 4213 48932 4219 48934
rect 4275 48932 4299 48934
rect 4355 48932 4379 48934
rect 4435 48932 4459 48934
rect 4515 48932 4521 48934
rect 4213 48912 4521 48932
rect 4213 47900 4521 47920
rect 4213 47898 4219 47900
rect 4275 47898 4299 47900
rect 4355 47898 4379 47900
rect 4435 47898 4459 47900
rect 4515 47898 4521 47900
rect 4275 47846 4277 47898
rect 4457 47846 4459 47898
rect 4213 47844 4219 47846
rect 4275 47844 4299 47846
rect 4355 47844 4379 47846
rect 4435 47844 4459 47846
rect 4515 47844 4521 47846
rect 4213 47824 4521 47844
rect 4068 47252 4120 47258
rect 4068 47194 4120 47200
rect 4213 46812 4521 46832
rect 4213 46810 4219 46812
rect 4275 46810 4299 46812
rect 4355 46810 4379 46812
rect 4435 46810 4459 46812
rect 4515 46810 4521 46812
rect 4275 46758 4277 46810
rect 4457 46758 4459 46810
rect 4213 46756 4219 46758
rect 4275 46756 4299 46758
rect 4355 46756 4379 46758
rect 4435 46756 4459 46758
rect 4515 46756 4521 46758
rect 4213 46736 4521 46756
rect 4068 46640 4120 46646
rect 4068 46582 4120 46588
rect 4080 45608 4108 46582
rect 4213 45724 4521 45744
rect 4213 45722 4219 45724
rect 4275 45722 4299 45724
rect 4355 45722 4379 45724
rect 4435 45722 4459 45724
rect 4515 45722 4521 45724
rect 4275 45670 4277 45722
rect 4457 45670 4459 45722
rect 4213 45668 4219 45670
rect 4275 45668 4299 45670
rect 4355 45668 4379 45670
rect 4435 45668 4459 45670
rect 4515 45668 4521 45670
rect 4213 45648 4521 45668
rect 4080 45580 4200 45608
rect 4068 45484 4120 45490
rect 4068 45426 4120 45432
rect 3976 44192 4028 44198
rect 3976 44134 4028 44140
rect 4080 43790 4108 45426
rect 4172 45422 4200 45580
rect 4160 45416 4212 45422
rect 4160 45358 4212 45364
rect 4172 44878 4200 45358
rect 4160 44872 4212 44878
rect 4160 44814 4212 44820
rect 4213 44636 4521 44656
rect 4213 44634 4219 44636
rect 4275 44634 4299 44636
rect 4355 44634 4379 44636
rect 4435 44634 4459 44636
rect 4515 44634 4521 44636
rect 4275 44582 4277 44634
rect 4457 44582 4459 44634
rect 4213 44580 4219 44582
rect 4275 44580 4299 44582
rect 4355 44580 4379 44582
rect 4435 44580 4459 44582
rect 4515 44580 4521 44582
rect 4213 44560 4521 44580
rect 4068 43784 4120 43790
rect 4068 43726 4120 43732
rect 3976 43376 4028 43382
rect 3976 43318 4028 43324
rect 3988 42786 4016 43318
rect 4080 42906 4108 43726
rect 4213 43548 4521 43568
rect 4213 43546 4219 43548
rect 4275 43546 4299 43548
rect 4355 43546 4379 43548
rect 4435 43546 4459 43548
rect 4515 43546 4521 43548
rect 4275 43494 4277 43546
rect 4457 43494 4459 43546
rect 4213 43492 4219 43494
rect 4275 43492 4299 43494
rect 4355 43492 4379 43494
rect 4435 43492 4459 43494
rect 4515 43492 4521 43494
rect 4213 43472 4521 43492
rect 4068 42900 4120 42906
rect 4068 42842 4120 42848
rect 3988 42758 4108 42786
rect 3976 42628 4028 42634
rect 3976 42570 4028 42576
rect 3884 40112 3936 40118
rect 3884 40054 3936 40060
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 3988 17270 4016 42570
rect 4080 24410 4108 42758
rect 4213 42460 4521 42480
rect 4213 42458 4219 42460
rect 4275 42458 4299 42460
rect 4355 42458 4379 42460
rect 4435 42458 4459 42460
rect 4515 42458 4521 42460
rect 4275 42406 4277 42458
rect 4457 42406 4459 42458
rect 4213 42404 4219 42406
rect 4275 42404 4299 42406
rect 4355 42404 4379 42406
rect 4435 42404 4459 42406
rect 4515 42404 4521 42406
rect 4213 42384 4521 42404
rect 4213 41372 4521 41392
rect 4213 41370 4219 41372
rect 4275 41370 4299 41372
rect 4355 41370 4379 41372
rect 4435 41370 4459 41372
rect 4515 41370 4521 41372
rect 4275 41318 4277 41370
rect 4457 41318 4459 41370
rect 4213 41316 4219 41318
rect 4275 41316 4299 41318
rect 4355 41316 4379 41318
rect 4435 41316 4459 41318
rect 4515 41316 4521 41318
rect 4213 41296 4521 41316
rect 4213 40284 4521 40304
rect 4213 40282 4219 40284
rect 4275 40282 4299 40284
rect 4355 40282 4379 40284
rect 4435 40282 4459 40284
rect 4515 40282 4521 40284
rect 4275 40230 4277 40282
rect 4457 40230 4459 40282
rect 4213 40228 4219 40230
rect 4275 40228 4299 40230
rect 4355 40228 4379 40230
rect 4435 40228 4459 40230
rect 4515 40228 4521 40230
rect 4213 40208 4521 40228
rect 4213 39196 4521 39216
rect 4213 39194 4219 39196
rect 4275 39194 4299 39196
rect 4355 39194 4379 39196
rect 4435 39194 4459 39196
rect 4515 39194 4521 39196
rect 4275 39142 4277 39194
rect 4457 39142 4459 39194
rect 4213 39140 4219 39142
rect 4275 39140 4299 39142
rect 4355 39140 4379 39142
rect 4435 39140 4459 39142
rect 4515 39140 4521 39142
rect 4213 39120 4521 39140
rect 4213 38108 4521 38128
rect 4213 38106 4219 38108
rect 4275 38106 4299 38108
rect 4355 38106 4379 38108
rect 4435 38106 4459 38108
rect 4515 38106 4521 38108
rect 4275 38054 4277 38106
rect 4457 38054 4459 38106
rect 4213 38052 4219 38054
rect 4275 38052 4299 38054
rect 4355 38052 4379 38054
rect 4435 38052 4459 38054
rect 4515 38052 4521 38054
rect 4213 38032 4521 38052
rect 4213 37020 4521 37040
rect 4213 37018 4219 37020
rect 4275 37018 4299 37020
rect 4355 37018 4379 37020
rect 4435 37018 4459 37020
rect 4515 37018 4521 37020
rect 4275 36966 4277 37018
rect 4457 36966 4459 37018
rect 4213 36964 4219 36966
rect 4275 36964 4299 36966
rect 4355 36964 4379 36966
rect 4435 36964 4459 36966
rect 4515 36964 4521 36966
rect 4213 36944 4521 36964
rect 4213 35932 4521 35952
rect 4213 35930 4219 35932
rect 4275 35930 4299 35932
rect 4355 35930 4379 35932
rect 4435 35930 4459 35932
rect 4515 35930 4521 35932
rect 4275 35878 4277 35930
rect 4457 35878 4459 35930
rect 4213 35876 4219 35878
rect 4275 35876 4299 35878
rect 4355 35876 4379 35878
rect 4435 35876 4459 35878
rect 4515 35876 4521 35878
rect 4213 35856 4521 35876
rect 4632 35086 4660 68206
rect 4712 52624 4764 52630
rect 4712 52566 4764 52572
rect 4724 48210 4752 52566
rect 4712 48204 4764 48210
rect 4712 48146 4764 48152
rect 4712 48068 4764 48074
rect 4712 48010 4764 48016
rect 4724 47598 4752 48010
rect 4712 47592 4764 47598
rect 4712 47534 4764 47540
rect 4712 47456 4764 47462
rect 4712 47398 4764 47404
rect 4724 46510 4752 47398
rect 4712 46504 4764 46510
rect 4712 46446 4764 46452
rect 4712 45552 4764 45558
rect 4712 45494 4764 45500
rect 4724 43858 4752 45494
rect 4712 43852 4764 43858
rect 4712 43794 4764 43800
rect 4712 43648 4764 43654
rect 4712 43590 4764 43596
rect 4620 35080 4672 35086
rect 4620 35022 4672 35028
rect 4213 34844 4521 34864
rect 4213 34842 4219 34844
rect 4275 34842 4299 34844
rect 4355 34842 4379 34844
rect 4435 34842 4459 34844
rect 4515 34842 4521 34844
rect 4275 34790 4277 34842
rect 4457 34790 4459 34842
rect 4213 34788 4219 34790
rect 4275 34788 4299 34790
rect 4355 34788 4379 34790
rect 4435 34788 4459 34790
rect 4515 34788 4521 34790
rect 4213 34768 4521 34788
rect 4213 33756 4521 33776
rect 4213 33754 4219 33756
rect 4275 33754 4299 33756
rect 4355 33754 4379 33756
rect 4435 33754 4459 33756
rect 4515 33754 4521 33756
rect 4275 33702 4277 33754
rect 4457 33702 4459 33754
rect 4213 33700 4219 33702
rect 4275 33700 4299 33702
rect 4355 33700 4379 33702
rect 4435 33700 4459 33702
rect 4515 33700 4521 33702
rect 4213 33680 4521 33700
rect 4213 32668 4521 32688
rect 4213 32666 4219 32668
rect 4275 32666 4299 32668
rect 4355 32666 4379 32668
rect 4435 32666 4459 32668
rect 4515 32666 4521 32668
rect 4275 32614 4277 32666
rect 4457 32614 4459 32666
rect 4213 32612 4219 32614
rect 4275 32612 4299 32614
rect 4355 32612 4379 32614
rect 4435 32612 4459 32614
rect 4515 32612 4521 32614
rect 4213 32592 4521 32612
rect 4213 31580 4521 31600
rect 4213 31578 4219 31580
rect 4275 31578 4299 31580
rect 4355 31578 4379 31580
rect 4435 31578 4459 31580
rect 4515 31578 4521 31580
rect 4275 31526 4277 31578
rect 4457 31526 4459 31578
rect 4213 31524 4219 31526
rect 4275 31524 4299 31526
rect 4355 31524 4379 31526
rect 4435 31524 4459 31526
rect 4515 31524 4521 31526
rect 4213 31504 4521 31524
rect 4213 30492 4521 30512
rect 4213 30490 4219 30492
rect 4275 30490 4299 30492
rect 4355 30490 4379 30492
rect 4435 30490 4459 30492
rect 4515 30490 4521 30492
rect 4275 30438 4277 30490
rect 4457 30438 4459 30490
rect 4213 30436 4219 30438
rect 4275 30436 4299 30438
rect 4355 30436 4379 30438
rect 4435 30436 4459 30438
rect 4515 30436 4521 30438
rect 4213 30416 4521 30436
rect 4213 29404 4521 29424
rect 4213 29402 4219 29404
rect 4275 29402 4299 29404
rect 4355 29402 4379 29404
rect 4435 29402 4459 29404
rect 4515 29402 4521 29404
rect 4275 29350 4277 29402
rect 4457 29350 4459 29402
rect 4213 29348 4219 29350
rect 4275 29348 4299 29350
rect 4355 29348 4379 29350
rect 4435 29348 4459 29350
rect 4515 29348 4521 29350
rect 4213 29328 4521 29348
rect 4213 28316 4521 28336
rect 4213 28314 4219 28316
rect 4275 28314 4299 28316
rect 4355 28314 4379 28316
rect 4435 28314 4459 28316
rect 4515 28314 4521 28316
rect 4275 28262 4277 28314
rect 4457 28262 4459 28314
rect 4213 28260 4219 28262
rect 4275 28260 4299 28262
rect 4355 28260 4379 28262
rect 4435 28260 4459 28262
rect 4515 28260 4521 28262
rect 4213 28240 4521 28260
rect 4213 27228 4521 27248
rect 4213 27226 4219 27228
rect 4275 27226 4299 27228
rect 4355 27226 4379 27228
rect 4435 27226 4459 27228
rect 4515 27226 4521 27228
rect 4275 27174 4277 27226
rect 4457 27174 4459 27226
rect 4213 27172 4219 27174
rect 4275 27172 4299 27174
rect 4355 27172 4379 27174
rect 4435 27172 4459 27174
rect 4515 27172 4521 27174
rect 4213 27152 4521 27172
rect 4213 26140 4521 26160
rect 4213 26138 4219 26140
rect 4275 26138 4299 26140
rect 4355 26138 4379 26140
rect 4435 26138 4459 26140
rect 4515 26138 4521 26140
rect 4275 26086 4277 26138
rect 4457 26086 4459 26138
rect 4213 26084 4219 26086
rect 4275 26084 4299 26086
rect 4355 26084 4379 26086
rect 4435 26084 4459 26086
rect 4515 26084 4521 26086
rect 4213 26064 4521 26084
rect 4213 25052 4521 25072
rect 4213 25050 4219 25052
rect 4275 25050 4299 25052
rect 4355 25050 4379 25052
rect 4435 25050 4459 25052
rect 4515 25050 4521 25052
rect 4275 24998 4277 25050
rect 4457 24998 4459 25050
rect 4213 24996 4219 24998
rect 4275 24996 4299 24998
rect 4355 24996 4379 24998
rect 4435 24996 4459 24998
rect 4515 24996 4521 24998
rect 4213 24976 4521 24996
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 4213 23964 4521 23984
rect 4213 23962 4219 23964
rect 4275 23962 4299 23964
rect 4355 23962 4379 23964
rect 4435 23962 4459 23964
rect 4515 23962 4521 23964
rect 4275 23910 4277 23962
rect 4457 23910 4459 23962
rect 4213 23908 4219 23910
rect 4275 23908 4299 23910
rect 4355 23908 4379 23910
rect 4435 23908 4459 23910
rect 4515 23908 4521 23910
rect 4213 23888 4521 23908
rect 4213 22876 4521 22896
rect 4213 22874 4219 22876
rect 4275 22874 4299 22876
rect 4355 22874 4379 22876
rect 4435 22874 4459 22876
rect 4515 22874 4521 22876
rect 4275 22822 4277 22874
rect 4457 22822 4459 22874
rect 4213 22820 4219 22822
rect 4275 22820 4299 22822
rect 4355 22820 4379 22822
rect 4435 22820 4459 22822
rect 4515 22820 4521 22822
rect 4213 22800 4521 22820
rect 4213 21788 4521 21808
rect 4213 21786 4219 21788
rect 4275 21786 4299 21788
rect 4355 21786 4379 21788
rect 4435 21786 4459 21788
rect 4515 21786 4521 21788
rect 4275 21734 4277 21786
rect 4457 21734 4459 21786
rect 4213 21732 4219 21734
rect 4275 21732 4299 21734
rect 4355 21732 4379 21734
rect 4435 21732 4459 21734
rect 4515 21732 4521 21734
rect 4213 21712 4521 21732
rect 4213 20700 4521 20720
rect 4213 20698 4219 20700
rect 4275 20698 4299 20700
rect 4355 20698 4379 20700
rect 4435 20698 4459 20700
rect 4515 20698 4521 20700
rect 4275 20646 4277 20698
rect 4457 20646 4459 20698
rect 4213 20644 4219 20646
rect 4275 20644 4299 20646
rect 4355 20644 4379 20646
rect 4435 20644 4459 20646
rect 4515 20644 4521 20646
rect 4213 20624 4521 20644
rect 4213 19612 4521 19632
rect 4213 19610 4219 19612
rect 4275 19610 4299 19612
rect 4355 19610 4379 19612
rect 4435 19610 4459 19612
rect 4515 19610 4521 19612
rect 4275 19558 4277 19610
rect 4457 19558 4459 19610
rect 4213 19556 4219 19558
rect 4275 19556 4299 19558
rect 4355 19556 4379 19558
rect 4435 19556 4459 19558
rect 4515 19556 4521 19558
rect 4213 19536 4521 19556
rect 4213 18524 4521 18544
rect 4213 18522 4219 18524
rect 4275 18522 4299 18524
rect 4355 18522 4379 18524
rect 4435 18522 4459 18524
rect 4515 18522 4521 18524
rect 4275 18470 4277 18522
rect 4457 18470 4459 18522
rect 4213 18468 4219 18470
rect 4275 18468 4299 18470
rect 4355 18468 4379 18470
rect 4435 18468 4459 18470
rect 4515 18468 4521 18470
rect 4213 18448 4521 18468
rect 4213 17436 4521 17456
rect 4213 17434 4219 17436
rect 4275 17434 4299 17436
rect 4355 17434 4379 17436
rect 4435 17434 4459 17436
rect 4515 17434 4521 17436
rect 4275 17382 4277 17434
rect 4457 17382 4459 17434
rect 4213 17380 4219 17382
rect 4275 17380 4299 17382
rect 4355 17380 4379 17382
rect 4435 17380 4459 17382
rect 4515 17380 4521 17382
rect 4213 17360 4521 17380
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 2582 16892 2890 16912
rect 2582 16890 2588 16892
rect 2644 16890 2668 16892
rect 2724 16890 2748 16892
rect 2804 16890 2828 16892
rect 2884 16890 2890 16892
rect 2644 16838 2646 16890
rect 2826 16838 2828 16890
rect 2582 16836 2588 16838
rect 2644 16836 2668 16838
rect 2724 16836 2748 16838
rect 2804 16836 2828 16838
rect 2884 16836 2890 16838
rect 2582 16816 2890 16836
rect 4213 16348 4521 16368
rect 4213 16346 4219 16348
rect 4275 16346 4299 16348
rect 4355 16346 4379 16348
rect 4435 16346 4459 16348
rect 4515 16346 4521 16348
rect 4275 16294 4277 16346
rect 4457 16294 4459 16346
rect 4213 16292 4219 16294
rect 4275 16292 4299 16294
rect 4355 16292 4379 16294
rect 4435 16292 4459 16294
rect 4515 16292 4521 16294
rect 4213 16272 4521 16292
rect 2582 15804 2890 15824
rect 2582 15802 2588 15804
rect 2644 15802 2668 15804
rect 2724 15802 2748 15804
rect 2804 15802 2828 15804
rect 2884 15802 2890 15804
rect 2644 15750 2646 15802
rect 2826 15750 2828 15802
rect 2582 15748 2588 15750
rect 2644 15748 2668 15750
rect 2724 15748 2748 15750
rect 2804 15748 2828 15750
rect 2884 15748 2890 15750
rect 2582 15728 2890 15748
rect 4213 15260 4521 15280
rect 4213 15258 4219 15260
rect 4275 15258 4299 15260
rect 4355 15258 4379 15260
rect 4435 15258 4459 15260
rect 4515 15258 4521 15260
rect 4275 15206 4277 15258
rect 4457 15206 4459 15258
rect 4213 15204 4219 15206
rect 4275 15204 4299 15206
rect 4355 15204 4379 15206
rect 4435 15204 4459 15206
rect 4515 15204 4521 15206
rect 4213 15184 4521 15204
rect 2582 14716 2890 14736
rect 2582 14714 2588 14716
rect 2644 14714 2668 14716
rect 2724 14714 2748 14716
rect 2804 14714 2828 14716
rect 2884 14714 2890 14716
rect 2644 14662 2646 14714
rect 2826 14662 2828 14714
rect 2582 14660 2588 14662
rect 2644 14660 2668 14662
rect 2724 14660 2748 14662
rect 2804 14660 2828 14662
rect 2884 14660 2890 14662
rect 2582 14640 2890 14660
rect 4213 14172 4521 14192
rect 4213 14170 4219 14172
rect 4275 14170 4299 14172
rect 4355 14170 4379 14172
rect 4435 14170 4459 14172
rect 4515 14170 4521 14172
rect 4275 14118 4277 14170
rect 4457 14118 4459 14170
rect 4213 14116 4219 14118
rect 4275 14116 4299 14118
rect 4355 14116 4379 14118
rect 4435 14116 4459 14118
rect 4515 14116 4521 14118
rect 4213 14096 4521 14116
rect 2582 13628 2890 13648
rect 2582 13626 2588 13628
rect 2644 13626 2668 13628
rect 2724 13626 2748 13628
rect 2804 13626 2828 13628
rect 2884 13626 2890 13628
rect 2644 13574 2646 13626
rect 2826 13574 2828 13626
rect 2582 13572 2588 13574
rect 2644 13572 2668 13574
rect 2724 13572 2748 13574
rect 2804 13572 2828 13574
rect 2884 13572 2890 13574
rect 2582 13552 2890 13572
rect 4213 13084 4521 13104
rect 4213 13082 4219 13084
rect 4275 13082 4299 13084
rect 4355 13082 4379 13084
rect 4435 13082 4459 13084
rect 4515 13082 4521 13084
rect 4275 13030 4277 13082
rect 4457 13030 4459 13082
rect 4213 13028 4219 13030
rect 4275 13028 4299 13030
rect 4355 13028 4379 13030
rect 4435 13028 4459 13030
rect 4515 13028 4521 13030
rect 4213 13008 4521 13028
rect 2582 12540 2890 12560
rect 2582 12538 2588 12540
rect 2644 12538 2668 12540
rect 2724 12538 2748 12540
rect 2804 12538 2828 12540
rect 2884 12538 2890 12540
rect 2644 12486 2646 12538
rect 2826 12486 2828 12538
rect 2582 12484 2588 12486
rect 2644 12484 2668 12486
rect 2724 12484 2748 12486
rect 2804 12484 2828 12486
rect 2884 12484 2890 12486
rect 2582 12464 2890 12484
rect 4213 11996 4521 12016
rect 4213 11994 4219 11996
rect 4275 11994 4299 11996
rect 4355 11994 4379 11996
rect 4435 11994 4459 11996
rect 4515 11994 4521 11996
rect 4275 11942 4277 11994
rect 4457 11942 4459 11994
rect 4213 11940 4219 11942
rect 4275 11940 4299 11942
rect 4355 11940 4379 11942
rect 4435 11940 4459 11942
rect 4515 11940 4521 11942
rect 4213 11920 4521 11940
rect 2582 11452 2890 11472
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 4213 10908 4521 10928
rect 4213 10906 4219 10908
rect 4275 10906 4299 10908
rect 4355 10906 4379 10908
rect 4435 10906 4459 10908
rect 4515 10906 4521 10908
rect 4275 10854 4277 10906
rect 4457 10854 4459 10906
rect 4213 10852 4219 10854
rect 4275 10852 4299 10854
rect 4355 10852 4379 10854
rect 4435 10852 4459 10854
rect 4515 10852 4521 10854
rect 4213 10832 4521 10852
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 4724 9994 4752 43590
rect 4816 38350 4844 71946
rect 5080 70508 5132 70514
rect 5080 70450 5132 70456
rect 4896 70440 4948 70446
rect 4896 70382 4948 70388
rect 4804 38344 4856 38350
rect 4804 38286 4856 38292
rect 4908 37874 4936 70382
rect 4988 61124 5040 61130
rect 4988 61066 5040 61072
rect 5000 40730 5028 61066
rect 5092 48822 5120 70450
rect 5632 66156 5684 66162
rect 5632 66098 5684 66104
rect 5172 66020 5224 66026
rect 5172 65962 5224 65968
rect 5080 48816 5132 48822
rect 5080 48758 5132 48764
rect 5080 47796 5132 47802
rect 5080 47738 5132 47744
rect 5092 46578 5120 47738
rect 5080 46572 5132 46578
rect 5080 46514 5132 46520
rect 5184 45778 5212 65962
rect 5356 61260 5408 61266
rect 5356 61202 5408 61208
rect 5264 57860 5316 57866
rect 5264 57802 5316 57808
rect 5276 50250 5304 57802
rect 5264 50244 5316 50250
rect 5264 50186 5316 50192
rect 5264 49972 5316 49978
rect 5264 49914 5316 49920
rect 5276 48226 5304 49914
rect 5368 48346 5396 61202
rect 5448 56976 5500 56982
rect 5448 56918 5500 56924
rect 5356 48340 5408 48346
rect 5356 48282 5408 48288
rect 5276 48198 5396 48226
rect 5264 48136 5316 48142
rect 5264 48078 5316 48084
rect 5092 45750 5212 45778
rect 5092 44266 5120 45750
rect 5172 45620 5224 45626
rect 5172 45562 5224 45568
rect 5080 44260 5132 44266
rect 5080 44202 5132 44208
rect 5080 43784 5132 43790
rect 5080 43726 5132 43732
rect 5092 42673 5120 43726
rect 5078 42664 5134 42673
rect 5078 42599 5134 42608
rect 5080 42288 5132 42294
rect 5080 42230 5132 42236
rect 4988 40724 5040 40730
rect 4988 40666 5040 40672
rect 5092 40610 5120 42230
rect 5184 42158 5212 45562
rect 5172 42152 5224 42158
rect 5172 42094 5224 42100
rect 5000 40582 5120 40610
rect 5000 39302 5028 40582
rect 5078 40488 5134 40497
rect 5078 40423 5134 40432
rect 4988 39296 5040 39302
rect 4988 39238 5040 39244
rect 4896 37868 4948 37874
rect 4896 37810 4948 37816
rect 4804 34740 4856 34746
rect 4804 34682 4856 34688
rect 4816 24206 4844 34682
rect 5000 33522 5028 39238
rect 4988 33516 5040 33522
rect 4988 33458 5040 33464
rect 4896 33040 4948 33046
rect 4896 32982 4948 32988
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4908 22642 4936 32982
rect 5092 31754 5120 40423
rect 5184 39438 5212 42094
rect 5172 39432 5224 39438
rect 5172 39374 5224 39380
rect 5172 39296 5224 39302
rect 5172 39238 5224 39244
rect 5184 32298 5212 39238
rect 5172 32292 5224 32298
rect 5172 32234 5224 32240
rect 5092 31726 5212 31754
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4213 9820 4521 9840
rect 4213 9818 4219 9820
rect 4275 9818 4299 9820
rect 4355 9818 4379 9820
rect 4435 9818 4459 9820
rect 4515 9818 4521 9820
rect 4275 9766 4277 9818
rect 4457 9766 4459 9818
rect 4213 9764 4219 9766
rect 4275 9764 4299 9766
rect 4355 9764 4379 9766
rect 4435 9764 4459 9766
rect 4515 9764 4521 9766
rect 4213 9744 4521 9764
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2582 9200 2890 9220
rect 4213 8732 4521 8752
rect 4213 8730 4219 8732
rect 4275 8730 4299 8732
rect 4355 8730 4379 8732
rect 4435 8730 4459 8732
rect 4515 8730 4521 8732
rect 4275 8678 4277 8730
rect 4457 8678 4459 8730
rect 4213 8676 4219 8678
rect 4275 8676 4299 8678
rect 4355 8676 4379 8678
rect 4435 8676 4459 8678
rect 4515 8676 4521 8678
rect 4213 8656 4521 8676
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 4213 7644 4521 7664
rect 4213 7642 4219 7644
rect 4275 7642 4299 7644
rect 4355 7642 4379 7644
rect 4435 7642 4459 7644
rect 4515 7642 4521 7644
rect 4275 7590 4277 7642
rect 4457 7590 4459 7642
rect 4213 7588 4219 7590
rect 4275 7588 4299 7590
rect 4355 7588 4379 7590
rect 4435 7588 4459 7590
rect 4515 7588 4521 7590
rect 4213 7568 4521 7588
rect 5184 7546 5212 31726
rect 5276 21978 5304 48078
rect 5368 43654 5396 48198
rect 5356 43648 5408 43654
rect 5356 43590 5408 43596
rect 5356 43376 5408 43382
rect 5356 43318 5408 43324
rect 5368 22094 5396 43318
rect 5460 41546 5488 56918
rect 5540 55752 5592 55758
rect 5540 55694 5592 55700
rect 5552 46714 5580 55694
rect 5540 46708 5592 46714
rect 5540 46650 5592 46656
rect 5644 44826 5672 66098
rect 5736 57390 5764 71946
rect 5845 71292 6153 71312
rect 5845 71290 5851 71292
rect 5907 71290 5931 71292
rect 5987 71290 6011 71292
rect 6067 71290 6091 71292
rect 6147 71290 6153 71292
rect 5907 71238 5909 71290
rect 6089 71238 6091 71290
rect 5845 71236 5851 71238
rect 5907 71236 5931 71238
rect 5987 71236 6011 71238
rect 6067 71236 6091 71238
rect 6147 71236 6153 71238
rect 5845 71216 6153 71236
rect 6196 70394 6224 72150
rect 6380 72010 6408 74054
rect 6656 72010 6684 74122
rect 6840 73710 6868 74258
rect 7477 74012 7785 74032
rect 7477 74010 7483 74012
rect 7539 74010 7563 74012
rect 7619 74010 7643 74012
rect 7699 74010 7723 74012
rect 7779 74010 7785 74012
rect 7539 73958 7541 74010
rect 7721 73958 7723 74010
rect 7477 73956 7483 73958
rect 7539 73956 7563 73958
rect 7619 73956 7643 73958
rect 7699 73956 7723 73958
rect 7779 73956 7785 73958
rect 7477 73936 7785 73956
rect 6828 73704 6880 73710
rect 6828 73646 6880 73652
rect 6840 73234 6868 73646
rect 6828 73228 6880 73234
rect 6828 73170 6880 73176
rect 6840 72162 6868 73170
rect 6920 73092 6972 73098
rect 6920 73034 6972 73040
rect 7380 73092 7432 73098
rect 7380 73034 7432 73040
rect 6932 72758 6960 73034
rect 7012 73024 7064 73030
rect 7288 73024 7340 73030
rect 7064 72972 7288 72978
rect 7012 72966 7340 72972
rect 7024 72950 7328 72966
rect 6920 72752 6972 72758
rect 6920 72694 6972 72700
rect 6840 72134 6960 72162
rect 6828 72072 6880 72078
rect 6828 72014 6880 72020
rect 6368 72004 6420 72010
rect 6368 71946 6420 71952
rect 6644 72004 6696 72010
rect 6644 71946 6696 71952
rect 6196 70366 6408 70394
rect 5845 70204 6153 70224
rect 5845 70202 5851 70204
rect 5907 70202 5931 70204
rect 5987 70202 6011 70204
rect 6067 70202 6091 70204
rect 6147 70202 6153 70204
rect 5907 70150 5909 70202
rect 6089 70150 6091 70202
rect 5845 70148 5851 70150
rect 5907 70148 5931 70150
rect 5987 70148 6011 70150
rect 6067 70148 6091 70150
rect 6147 70148 6153 70150
rect 5845 70128 6153 70148
rect 5845 69116 6153 69136
rect 5845 69114 5851 69116
rect 5907 69114 5931 69116
rect 5987 69114 6011 69116
rect 6067 69114 6091 69116
rect 6147 69114 6153 69116
rect 5907 69062 5909 69114
rect 6089 69062 6091 69114
rect 5845 69060 5851 69062
rect 5907 69060 5931 69062
rect 5987 69060 6011 69062
rect 6067 69060 6091 69062
rect 6147 69060 6153 69062
rect 5845 69040 6153 69060
rect 5845 68028 6153 68048
rect 5845 68026 5851 68028
rect 5907 68026 5931 68028
rect 5987 68026 6011 68028
rect 6067 68026 6091 68028
rect 6147 68026 6153 68028
rect 5907 67974 5909 68026
rect 6089 67974 6091 68026
rect 5845 67972 5851 67974
rect 5907 67972 5931 67974
rect 5987 67972 6011 67974
rect 6067 67972 6091 67974
rect 6147 67972 6153 67974
rect 5845 67952 6153 67972
rect 5845 66940 6153 66960
rect 5845 66938 5851 66940
rect 5907 66938 5931 66940
rect 5987 66938 6011 66940
rect 6067 66938 6091 66940
rect 6147 66938 6153 66940
rect 5907 66886 5909 66938
rect 6089 66886 6091 66938
rect 5845 66884 5851 66886
rect 5907 66884 5931 66886
rect 5987 66884 6011 66886
rect 6067 66884 6091 66886
rect 6147 66884 6153 66886
rect 5845 66864 6153 66884
rect 6276 66564 6328 66570
rect 6276 66506 6328 66512
rect 5845 65852 6153 65872
rect 5845 65850 5851 65852
rect 5907 65850 5931 65852
rect 5987 65850 6011 65852
rect 6067 65850 6091 65852
rect 6147 65850 6153 65852
rect 5907 65798 5909 65850
rect 6089 65798 6091 65850
rect 5845 65796 5851 65798
rect 5907 65796 5931 65798
rect 5987 65796 6011 65798
rect 6067 65796 6091 65798
rect 6147 65796 6153 65798
rect 5845 65776 6153 65796
rect 5845 64764 6153 64784
rect 5845 64762 5851 64764
rect 5907 64762 5931 64764
rect 5987 64762 6011 64764
rect 6067 64762 6091 64764
rect 6147 64762 6153 64764
rect 5907 64710 5909 64762
rect 6089 64710 6091 64762
rect 5845 64708 5851 64710
rect 5907 64708 5931 64710
rect 5987 64708 6011 64710
rect 6067 64708 6091 64710
rect 6147 64708 6153 64710
rect 5845 64688 6153 64708
rect 5845 63676 6153 63696
rect 5845 63674 5851 63676
rect 5907 63674 5931 63676
rect 5987 63674 6011 63676
rect 6067 63674 6091 63676
rect 6147 63674 6153 63676
rect 5907 63622 5909 63674
rect 6089 63622 6091 63674
rect 5845 63620 5851 63622
rect 5907 63620 5931 63622
rect 5987 63620 6011 63622
rect 6067 63620 6091 63622
rect 6147 63620 6153 63622
rect 5845 63600 6153 63620
rect 6184 62756 6236 62762
rect 6184 62698 6236 62704
rect 5845 62588 6153 62608
rect 5845 62586 5851 62588
rect 5907 62586 5931 62588
rect 5987 62586 6011 62588
rect 6067 62586 6091 62588
rect 6147 62586 6153 62588
rect 5907 62534 5909 62586
rect 6089 62534 6091 62586
rect 5845 62532 5851 62534
rect 5907 62532 5931 62534
rect 5987 62532 6011 62534
rect 6067 62532 6091 62534
rect 6147 62532 6153 62534
rect 5845 62512 6153 62532
rect 5845 61500 6153 61520
rect 5845 61498 5851 61500
rect 5907 61498 5931 61500
rect 5987 61498 6011 61500
rect 6067 61498 6091 61500
rect 6147 61498 6153 61500
rect 5907 61446 5909 61498
rect 6089 61446 6091 61498
rect 5845 61444 5851 61446
rect 5907 61444 5931 61446
rect 5987 61444 6011 61446
rect 6067 61444 6091 61446
rect 6147 61444 6153 61446
rect 5845 61424 6153 61444
rect 5845 60412 6153 60432
rect 5845 60410 5851 60412
rect 5907 60410 5931 60412
rect 5987 60410 6011 60412
rect 6067 60410 6091 60412
rect 6147 60410 6153 60412
rect 5907 60358 5909 60410
rect 6089 60358 6091 60410
rect 5845 60356 5851 60358
rect 5907 60356 5931 60358
rect 5987 60356 6011 60358
rect 6067 60356 6091 60358
rect 6147 60356 6153 60358
rect 5845 60336 6153 60356
rect 5845 59324 6153 59344
rect 5845 59322 5851 59324
rect 5907 59322 5931 59324
rect 5987 59322 6011 59324
rect 6067 59322 6091 59324
rect 6147 59322 6153 59324
rect 5907 59270 5909 59322
rect 6089 59270 6091 59322
rect 5845 59268 5851 59270
rect 5907 59268 5931 59270
rect 5987 59268 6011 59270
rect 6067 59268 6091 59270
rect 6147 59268 6153 59270
rect 5845 59248 6153 59268
rect 5845 58236 6153 58256
rect 5845 58234 5851 58236
rect 5907 58234 5931 58236
rect 5987 58234 6011 58236
rect 6067 58234 6091 58236
rect 6147 58234 6153 58236
rect 5907 58182 5909 58234
rect 6089 58182 6091 58234
rect 5845 58180 5851 58182
rect 5907 58180 5931 58182
rect 5987 58180 6011 58182
rect 6067 58180 6091 58182
rect 6147 58180 6153 58182
rect 5845 58160 6153 58180
rect 5724 57384 5776 57390
rect 5724 57326 5776 57332
rect 5724 57248 5776 57254
rect 5724 57190 5776 57196
rect 5736 57050 5764 57190
rect 5845 57148 6153 57168
rect 5845 57146 5851 57148
rect 5907 57146 5931 57148
rect 5987 57146 6011 57148
rect 6067 57146 6091 57148
rect 6147 57146 6153 57148
rect 5907 57094 5909 57146
rect 6089 57094 6091 57146
rect 5845 57092 5851 57094
rect 5907 57092 5931 57094
rect 5987 57092 6011 57094
rect 6067 57092 6091 57094
rect 6147 57092 6153 57094
rect 5845 57072 6153 57092
rect 5724 57044 5776 57050
rect 5724 56986 5776 56992
rect 5845 56060 6153 56080
rect 5845 56058 5851 56060
rect 5907 56058 5931 56060
rect 5987 56058 6011 56060
rect 6067 56058 6091 56060
rect 6147 56058 6153 56060
rect 5907 56006 5909 56058
rect 6089 56006 6091 56058
rect 5845 56004 5851 56006
rect 5907 56004 5931 56006
rect 5987 56004 6011 56006
rect 6067 56004 6091 56006
rect 6147 56004 6153 56006
rect 5845 55984 6153 56004
rect 5845 54972 6153 54992
rect 5845 54970 5851 54972
rect 5907 54970 5931 54972
rect 5987 54970 6011 54972
rect 6067 54970 6091 54972
rect 6147 54970 6153 54972
rect 5907 54918 5909 54970
rect 6089 54918 6091 54970
rect 5845 54916 5851 54918
rect 5907 54916 5931 54918
rect 5987 54916 6011 54918
rect 6067 54916 6091 54918
rect 6147 54916 6153 54918
rect 5845 54896 6153 54916
rect 5845 53884 6153 53904
rect 5845 53882 5851 53884
rect 5907 53882 5931 53884
rect 5987 53882 6011 53884
rect 6067 53882 6091 53884
rect 6147 53882 6153 53884
rect 5907 53830 5909 53882
rect 6089 53830 6091 53882
rect 5845 53828 5851 53830
rect 5907 53828 5931 53830
rect 5987 53828 6011 53830
rect 6067 53828 6091 53830
rect 6147 53828 6153 53830
rect 5845 53808 6153 53828
rect 5845 52796 6153 52816
rect 5845 52794 5851 52796
rect 5907 52794 5931 52796
rect 5987 52794 6011 52796
rect 6067 52794 6091 52796
rect 6147 52794 6153 52796
rect 5907 52742 5909 52794
rect 6089 52742 6091 52794
rect 5845 52740 5851 52742
rect 5907 52740 5931 52742
rect 5987 52740 6011 52742
rect 6067 52740 6091 52742
rect 6147 52740 6153 52742
rect 5845 52720 6153 52740
rect 5845 51708 6153 51728
rect 5845 51706 5851 51708
rect 5907 51706 5931 51708
rect 5987 51706 6011 51708
rect 6067 51706 6091 51708
rect 6147 51706 6153 51708
rect 5907 51654 5909 51706
rect 6089 51654 6091 51706
rect 5845 51652 5851 51654
rect 5907 51652 5931 51654
rect 5987 51652 6011 51654
rect 6067 51652 6091 51654
rect 6147 51652 6153 51654
rect 5845 51632 6153 51652
rect 5845 50620 6153 50640
rect 5845 50618 5851 50620
rect 5907 50618 5931 50620
rect 5987 50618 6011 50620
rect 6067 50618 6091 50620
rect 6147 50618 6153 50620
rect 5907 50566 5909 50618
rect 6089 50566 6091 50618
rect 5845 50564 5851 50566
rect 5907 50564 5931 50566
rect 5987 50564 6011 50566
rect 6067 50564 6091 50566
rect 6147 50564 6153 50566
rect 5845 50544 6153 50564
rect 5845 49532 6153 49552
rect 5845 49530 5851 49532
rect 5907 49530 5931 49532
rect 5987 49530 6011 49532
rect 6067 49530 6091 49532
rect 6147 49530 6153 49532
rect 5907 49478 5909 49530
rect 6089 49478 6091 49530
rect 5845 49476 5851 49478
rect 5907 49476 5931 49478
rect 5987 49476 6011 49478
rect 6067 49476 6091 49478
rect 6147 49476 6153 49478
rect 5845 49456 6153 49476
rect 5845 48444 6153 48464
rect 5845 48442 5851 48444
rect 5907 48442 5931 48444
rect 5987 48442 6011 48444
rect 6067 48442 6091 48444
rect 6147 48442 6153 48444
rect 5907 48390 5909 48442
rect 6089 48390 6091 48442
rect 5845 48388 5851 48390
rect 5907 48388 5931 48390
rect 5987 48388 6011 48390
rect 6067 48388 6091 48390
rect 6147 48388 6153 48390
rect 5845 48368 6153 48388
rect 5724 47456 5776 47462
rect 5724 47398 5776 47404
rect 5736 46646 5764 47398
rect 5845 47356 6153 47376
rect 5845 47354 5851 47356
rect 5907 47354 5931 47356
rect 5987 47354 6011 47356
rect 6067 47354 6091 47356
rect 6147 47354 6153 47356
rect 5907 47302 5909 47354
rect 6089 47302 6091 47354
rect 5845 47300 5851 47302
rect 5907 47300 5931 47302
rect 5987 47300 6011 47302
rect 6067 47300 6091 47302
rect 6147 47300 6153 47302
rect 5845 47280 6153 47300
rect 5724 46640 5776 46646
rect 5724 46582 5776 46588
rect 5724 46504 5776 46510
rect 5724 46446 5776 46452
rect 5552 44798 5672 44826
rect 5448 41540 5500 41546
rect 5448 41482 5500 41488
rect 5552 41274 5580 44798
rect 5632 44736 5684 44742
rect 5632 44678 5684 44684
rect 5540 41268 5592 41274
rect 5540 41210 5592 41216
rect 5448 40724 5500 40730
rect 5448 40666 5500 40672
rect 5460 32434 5488 40666
rect 5644 40526 5672 44678
rect 5632 40520 5684 40526
rect 5632 40462 5684 40468
rect 5632 40384 5684 40390
rect 5632 40326 5684 40332
rect 5644 39302 5672 40326
rect 5632 39296 5684 39302
rect 5632 39238 5684 39244
rect 5632 37188 5684 37194
rect 5632 37130 5684 37136
rect 5540 36304 5592 36310
rect 5540 36246 5592 36252
rect 5448 32428 5500 32434
rect 5448 32370 5500 32376
rect 5448 32292 5500 32298
rect 5448 32234 5500 32240
rect 5460 23186 5488 32234
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5368 22066 5488 22094
rect 5276 21950 5396 21978
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5276 14550 5304 21830
rect 5368 17814 5396 21950
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5368 15706 5396 15846
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5354 13424 5410 13433
rect 5354 13359 5356 13368
rect 5408 13359 5410 13368
rect 5356 13330 5408 13336
rect 5460 9178 5488 22066
rect 5552 9382 5580 36246
rect 5644 35834 5672 37130
rect 5632 35828 5684 35834
rect 5632 35770 5684 35776
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5644 17746 5672 22918
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5644 14074 5672 14894
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 13394 5672 13670
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 10810 5672 12786
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 4213 6556 4521 6576
rect 4213 6554 4219 6556
rect 4275 6554 4299 6556
rect 4355 6554 4379 6556
rect 4435 6554 4459 6556
rect 4515 6554 4521 6556
rect 4275 6502 4277 6554
rect 4457 6502 4459 6554
rect 4213 6500 4219 6502
rect 4275 6500 4299 6502
rect 4355 6500 4379 6502
rect 4435 6500 4459 6502
rect 4515 6500 4521 6502
rect 4213 6480 4521 6500
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 5736 5710 5764 46446
rect 5845 46268 6153 46288
rect 5845 46266 5851 46268
rect 5907 46266 5931 46268
rect 5987 46266 6011 46268
rect 6067 46266 6091 46268
rect 6147 46266 6153 46268
rect 5907 46214 5909 46266
rect 6089 46214 6091 46266
rect 5845 46212 5851 46214
rect 5907 46212 5931 46214
rect 5987 46212 6011 46214
rect 6067 46212 6091 46214
rect 6147 46212 6153 46214
rect 5845 46192 6153 46212
rect 5845 45180 6153 45200
rect 5845 45178 5851 45180
rect 5907 45178 5931 45180
rect 5987 45178 6011 45180
rect 6067 45178 6091 45180
rect 6147 45178 6153 45180
rect 5907 45126 5909 45178
rect 6089 45126 6091 45178
rect 5845 45124 5851 45126
rect 5907 45124 5931 45126
rect 5987 45124 6011 45126
rect 6067 45124 6091 45126
rect 6147 45124 6153 45126
rect 5845 45104 6153 45124
rect 5845 44092 6153 44112
rect 5845 44090 5851 44092
rect 5907 44090 5931 44092
rect 5987 44090 6011 44092
rect 6067 44090 6091 44092
rect 6147 44090 6153 44092
rect 5907 44038 5909 44090
rect 6089 44038 6091 44090
rect 5845 44036 5851 44038
rect 5907 44036 5931 44038
rect 5987 44036 6011 44038
rect 6067 44036 6091 44038
rect 6147 44036 6153 44038
rect 5845 44016 6153 44036
rect 5845 43004 6153 43024
rect 5845 43002 5851 43004
rect 5907 43002 5931 43004
rect 5987 43002 6011 43004
rect 6067 43002 6091 43004
rect 6147 43002 6153 43004
rect 5907 42950 5909 43002
rect 6089 42950 6091 43002
rect 5845 42948 5851 42950
rect 5907 42948 5931 42950
rect 5987 42948 6011 42950
rect 6067 42948 6091 42950
rect 6147 42948 6153 42950
rect 5845 42928 6153 42948
rect 6090 42664 6146 42673
rect 6090 42599 6146 42608
rect 6104 42226 6132 42599
rect 6092 42220 6144 42226
rect 6092 42162 6144 42168
rect 5845 41916 6153 41936
rect 5845 41914 5851 41916
rect 5907 41914 5931 41916
rect 5987 41914 6011 41916
rect 6067 41914 6091 41916
rect 6147 41914 6153 41916
rect 5907 41862 5909 41914
rect 6089 41862 6091 41914
rect 5845 41860 5851 41862
rect 5907 41860 5931 41862
rect 5987 41860 6011 41862
rect 6067 41860 6091 41862
rect 6147 41860 6153 41862
rect 5845 41840 6153 41860
rect 5845 40828 6153 40848
rect 5845 40826 5851 40828
rect 5907 40826 5931 40828
rect 5987 40826 6011 40828
rect 6067 40826 6091 40828
rect 6147 40826 6153 40828
rect 5907 40774 5909 40826
rect 6089 40774 6091 40826
rect 5845 40772 5851 40774
rect 5907 40772 5931 40774
rect 5987 40772 6011 40774
rect 6067 40772 6091 40774
rect 6147 40772 6153 40774
rect 5845 40752 6153 40772
rect 5845 39740 6153 39760
rect 5845 39738 5851 39740
rect 5907 39738 5931 39740
rect 5987 39738 6011 39740
rect 6067 39738 6091 39740
rect 6147 39738 6153 39740
rect 5907 39686 5909 39738
rect 6089 39686 6091 39738
rect 5845 39684 5851 39686
rect 5907 39684 5931 39686
rect 5987 39684 6011 39686
rect 6067 39684 6091 39686
rect 6147 39684 6153 39686
rect 5845 39664 6153 39684
rect 5845 38652 6153 38672
rect 5845 38650 5851 38652
rect 5907 38650 5931 38652
rect 5987 38650 6011 38652
rect 6067 38650 6091 38652
rect 6147 38650 6153 38652
rect 5907 38598 5909 38650
rect 6089 38598 6091 38650
rect 5845 38596 5851 38598
rect 5907 38596 5931 38598
rect 5987 38596 6011 38598
rect 6067 38596 6091 38598
rect 6147 38596 6153 38598
rect 5845 38576 6153 38596
rect 5845 37564 6153 37584
rect 5845 37562 5851 37564
rect 5907 37562 5931 37564
rect 5987 37562 6011 37564
rect 6067 37562 6091 37564
rect 6147 37562 6153 37564
rect 5907 37510 5909 37562
rect 6089 37510 6091 37562
rect 5845 37508 5851 37510
rect 5907 37508 5931 37510
rect 5987 37508 6011 37510
rect 6067 37508 6091 37510
rect 6147 37508 6153 37510
rect 5845 37488 6153 37508
rect 5845 36476 6153 36496
rect 5845 36474 5851 36476
rect 5907 36474 5931 36476
rect 5987 36474 6011 36476
rect 6067 36474 6091 36476
rect 6147 36474 6153 36476
rect 5907 36422 5909 36474
rect 6089 36422 6091 36474
rect 5845 36420 5851 36422
rect 5907 36420 5931 36422
rect 5987 36420 6011 36422
rect 6067 36420 6091 36422
rect 6147 36420 6153 36422
rect 5845 36400 6153 36420
rect 5845 35388 6153 35408
rect 5845 35386 5851 35388
rect 5907 35386 5931 35388
rect 5987 35386 6011 35388
rect 6067 35386 6091 35388
rect 6147 35386 6153 35388
rect 5907 35334 5909 35386
rect 6089 35334 6091 35386
rect 5845 35332 5851 35334
rect 5907 35332 5931 35334
rect 5987 35332 6011 35334
rect 6067 35332 6091 35334
rect 6147 35332 6153 35334
rect 5845 35312 6153 35332
rect 5845 34300 6153 34320
rect 5845 34298 5851 34300
rect 5907 34298 5931 34300
rect 5987 34298 6011 34300
rect 6067 34298 6091 34300
rect 6147 34298 6153 34300
rect 5907 34246 5909 34298
rect 6089 34246 6091 34298
rect 5845 34244 5851 34246
rect 5907 34244 5931 34246
rect 5987 34244 6011 34246
rect 6067 34244 6091 34246
rect 6147 34244 6153 34246
rect 5845 34224 6153 34244
rect 5845 33212 6153 33232
rect 5845 33210 5851 33212
rect 5907 33210 5931 33212
rect 5987 33210 6011 33212
rect 6067 33210 6091 33212
rect 6147 33210 6153 33212
rect 5907 33158 5909 33210
rect 6089 33158 6091 33210
rect 5845 33156 5851 33158
rect 5907 33156 5931 33158
rect 5987 33156 6011 33158
rect 6067 33156 6091 33158
rect 6147 33156 6153 33158
rect 5845 33136 6153 33156
rect 5845 32124 6153 32144
rect 5845 32122 5851 32124
rect 5907 32122 5931 32124
rect 5987 32122 6011 32124
rect 6067 32122 6091 32124
rect 6147 32122 6153 32124
rect 5907 32070 5909 32122
rect 6089 32070 6091 32122
rect 5845 32068 5851 32070
rect 5907 32068 5931 32070
rect 5987 32068 6011 32070
rect 6067 32068 6091 32070
rect 6147 32068 6153 32070
rect 5845 32048 6153 32068
rect 6196 31890 6224 62698
rect 6288 38298 6316 66506
rect 6380 44742 6408 70366
rect 6840 69018 6868 72014
rect 6932 72010 6960 72134
rect 6920 72004 6972 72010
rect 6920 71946 6972 71952
rect 6932 71058 6960 71946
rect 7104 71120 7156 71126
rect 7104 71062 7156 71068
rect 6920 71052 6972 71058
rect 6920 70994 6972 71000
rect 6828 69012 6880 69018
rect 6828 68954 6880 68960
rect 7012 68740 7064 68746
rect 7012 68682 7064 68688
rect 6920 67720 6972 67726
rect 6920 67662 6972 67668
rect 6736 65544 6788 65550
rect 6736 65486 6788 65492
rect 6552 65476 6604 65482
rect 6552 65418 6604 65424
rect 6460 63300 6512 63306
rect 6460 63242 6512 63248
rect 6368 44736 6420 44742
rect 6368 44678 6420 44684
rect 6368 43308 6420 43314
rect 6368 43250 6420 43256
rect 6380 42770 6408 43250
rect 6368 42764 6420 42770
rect 6368 42706 6420 42712
rect 6368 42560 6420 42566
rect 6368 42502 6420 42508
rect 6380 42294 6408 42502
rect 6368 42288 6420 42294
rect 6368 42230 6420 42236
rect 6368 42016 6420 42022
rect 6368 41958 6420 41964
rect 6380 41750 6408 41958
rect 6368 41744 6420 41750
rect 6368 41686 6420 41692
rect 6472 41414 6500 63242
rect 6564 53990 6592 65418
rect 6644 56840 6696 56846
rect 6644 56782 6696 56788
rect 6552 53984 6604 53990
rect 6552 53926 6604 53932
rect 6656 51610 6684 56782
rect 6644 51604 6696 51610
rect 6644 51546 6696 51552
rect 6644 51264 6696 51270
rect 6644 51206 6696 51212
rect 6552 49904 6604 49910
rect 6552 49846 6604 49852
rect 6564 42634 6592 49846
rect 6656 49434 6684 51206
rect 6644 49428 6696 49434
rect 6644 49370 6696 49376
rect 6644 47116 6696 47122
rect 6644 47058 6696 47064
rect 6656 43382 6684 47058
rect 6644 43376 6696 43382
rect 6644 43318 6696 43324
rect 6642 43072 6698 43081
rect 6642 43007 6698 43016
rect 6552 42628 6604 42634
rect 6552 42570 6604 42576
rect 6552 42288 6604 42294
rect 6552 42230 6604 42236
rect 6380 41386 6500 41414
rect 6380 38418 6408 41386
rect 6460 41132 6512 41138
rect 6460 41074 6512 41080
rect 6472 40118 6500 41074
rect 6460 40112 6512 40118
rect 6460 40054 6512 40060
rect 6368 38412 6420 38418
rect 6368 38354 6420 38360
rect 6288 38270 6408 38298
rect 6276 36916 6328 36922
rect 6276 36858 6328 36864
rect 6288 36242 6316 36858
rect 6276 36236 6328 36242
rect 6276 36178 6328 36184
rect 6380 35766 6408 38270
rect 6368 35760 6420 35766
rect 6368 35702 6420 35708
rect 6472 34066 6500 40054
rect 6564 39982 6592 42230
rect 6552 39976 6604 39982
rect 6552 39918 6604 39924
rect 6552 39840 6604 39846
rect 6552 39782 6604 39788
rect 6564 39506 6592 39782
rect 6552 39500 6604 39506
rect 6552 39442 6604 39448
rect 6564 39302 6592 39442
rect 6552 39296 6604 39302
rect 6552 39238 6604 39244
rect 6550 39128 6606 39137
rect 6550 39063 6606 39072
rect 6460 34060 6512 34066
rect 6460 34002 6512 34008
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 5845 31036 6153 31056
rect 5845 31034 5851 31036
rect 5907 31034 5931 31036
rect 5987 31034 6011 31036
rect 6067 31034 6091 31036
rect 6147 31034 6153 31036
rect 5907 30982 5909 31034
rect 6089 30982 6091 31034
rect 5845 30980 5851 30982
rect 5907 30980 5931 30982
rect 5987 30980 6011 30982
rect 6067 30980 6091 30982
rect 6147 30980 6153 30982
rect 5845 30960 6153 30980
rect 5845 29948 6153 29968
rect 5845 29946 5851 29948
rect 5907 29946 5931 29948
rect 5987 29946 6011 29948
rect 6067 29946 6091 29948
rect 6147 29946 6153 29948
rect 5907 29894 5909 29946
rect 6089 29894 6091 29946
rect 5845 29892 5851 29894
rect 5907 29892 5931 29894
rect 5987 29892 6011 29894
rect 6067 29892 6091 29894
rect 6147 29892 6153 29894
rect 5845 29872 6153 29892
rect 5845 28860 6153 28880
rect 5845 28858 5851 28860
rect 5907 28858 5931 28860
rect 5987 28858 6011 28860
rect 6067 28858 6091 28860
rect 6147 28858 6153 28860
rect 5907 28806 5909 28858
rect 6089 28806 6091 28858
rect 5845 28804 5851 28806
rect 5907 28804 5931 28806
rect 5987 28804 6011 28806
rect 6067 28804 6091 28806
rect 6147 28804 6153 28806
rect 5845 28784 6153 28804
rect 5845 27772 6153 27792
rect 5845 27770 5851 27772
rect 5907 27770 5931 27772
rect 5987 27770 6011 27772
rect 6067 27770 6091 27772
rect 6147 27770 6153 27772
rect 5907 27718 5909 27770
rect 6089 27718 6091 27770
rect 5845 27716 5851 27718
rect 5907 27716 5931 27718
rect 5987 27716 6011 27718
rect 6067 27716 6091 27718
rect 6147 27716 6153 27718
rect 5845 27696 6153 27716
rect 5845 26684 6153 26704
rect 5845 26682 5851 26684
rect 5907 26682 5931 26684
rect 5987 26682 6011 26684
rect 6067 26682 6091 26684
rect 6147 26682 6153 26684
rect 5907 26630 5909 26682
rect 6089 26630 6091 26682
rect 5845 26628 5851 26630
rect 5907 26628 5931 26630
rect 5987 26628 6011 26630
rect 6067 26628 6091 26630
rect 6147 26628 6153 26630
rect 5845 26608 6153 26628
rect 5845 25596 6153 25616
rect 5845 25594 5851 25596
rect 5907 25594 5931 25596
rect 5987 25594 6011 25596
rect 6067 25594 6091 25596
rect 6147 25594 6153 25596
rect 5907 25542 5909 25594
rect 6089 25542 6091 25594
rect 5845 25540 5851 25542
rect 5907 25540 5931 25542
rect 5987 25540 6011 25542
rect 6067 25540 6091 25542
rect 6147 25540 6153 25542
rect 5845 25520 6153 25540
rect 5845 24508 6153 24528
rect 5845 24506 5851 24508
rect 5907 24506 5931 24508
rect 5987 24506 6011 24508
rect 6067 24506 6091 24508
rect 6147 24506 6153 24508
rect 5907 24454 5909 24506
rect 6089 24454 6091 24506
rect 5845 24452 5851 24454
rect 5907 24452 5931 24454
rect 5987 24452 6011 24454
rect 6067 24452 6091 24454
rect 6147 24452 6153 24454
rect 5845 24432 6153 24452
rect 5845 23420 6153 23440
rect 5845 23418 5851 23420
rect 5907 23418 5931 23420
rect 5987 23418 6011 23420
rect 6067 23418 6091 23420
rect 6147 23418 6153 23420
rect 5907 23366 5909 23418
rect 6089 23366 6091 23418
rect 5845 23364 5851 23366
rect 5907 23364 5931 23366
rect 5987 23364 6011 23366
rect 6067 23364 6091 23366
rect 6147 23364 6153 23366
rect 5845 23344 6153 23364
rect 6564 22710 6592 39063
rect 6552 22704 6604 22710
rect 6552 22646 6604 22652
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 5845 22332 6153 22352
rect 5845 22330 5851 22332
rect 5907 22330 5931 22332
rect 5987 22330 6011 22332
rect 6067 22330 6091 22332
rect 6147 22330 6153 22332
rect 5907 22278 5909 22330
rect 6089 22278 6091 22330
rect 5845 22276 5851 22278
rect 5907 22276 5931 22278
rect 5987 22276 6011 22278
rect 6067 22276 6091 22278
rect 6147 22276 6153 22278
rect 5845 22256 6153 22276
rect 5845 21244 6153 21264
rect 5845 21242 5851 21244
rect 5907 21242 5931 21244
rect 5987 21242 6011 21244
rect 6067 21242 6091 21244
rect 6147 21242 6153 21244
rect 5907 21190 5909 21242
rect 6089 21190 6091 21242
rect 5845 21188 5851 21190
rect 5907 21188 5931 21190
rect 5987 21188 6011 21190
rect 6067 21188 6091 21190
rect 6147 21188 6153 21190
rect 5845 21168 6153 21188
rect 5845 20156 6153 20176
rect 5845 20154 5851 20156
rect 5907 20154 5931 20156
rect 5987 20154 6011 20156
rect 6067 20154 6091 20156
rect 6147 20154 6153 20156
rect 5907 20102 5909 20154
rect 6089 20102 6091 20154
rect 5845 20100 5851 20102
rect 5907 20100 5931 20102
rect 5987 20100 6011 20102
rect 6067 20100 6091 20102
rect 6147 20100 6153 20102
rect 5845 20080 6153 20100
rect 5845 19068 6153 19088
rect 5845 19066 5851 19068
rect 5907 19066 5931 19068
rect 5987 19066 6011 19068
rect 6067 19066 6091 19068
rect 6147 19066 6153 19068
rect 5907 19014 5909 19066
rect 6089 19014 6091 19066
rect 5845 19012 5851 19014
rect 5907 19012 5931 19014
rect 5987 19012 6011 19014
rect 6067 19012 6091 19014
rect 6147 19012 6153 19014
rect 5845 18992 6153 19012
rect 5845 17980 6153 18000
rect 5845 17978 5851 17980
rect 5907 17978 5931 17980
rect 5987 17978 6011 17980
rect 6067 17978 6091 17980
rect 6147 17978 6153 17980
rect 5907 17926 5909 17978
rect 6089 17926 6091 17978
rect 5845 17924 5851 17926
rect 5907 17924 5931 17926
rect 5987 17924 6011 17926
rect 6067 17924 6091 17926
rect 6147 17924 6153 17926
rect 5845 17904 6153 17924
rect 6196 17202 6224 22442
rect 6656 22094 6684 43007
rect 6748 26042 6776 65486
rect 6828 51808 6880 51814
rect 6828 51750 6880 51756
rect 6840 49910 6868 51750
rect 6828 49904 6880 49910
rect 6828 49846 6880 49852
rect 6828 49768 6880 49774
rect 6828 49710 6880 49716
rect 6840 42906 6868 49710
rect 6932 46050 6960 67662
rect 7024 66638 7052 68682
rect 7012 66632 7064 66638
rect 7012 66574 7064 66580
rect 7024 51241 7052 66574
rect 7116 62286 7144 71062
rect 7300 70514 7328 72950
rect 7288 70508 7340 70514
rect 7288 70450 7340 70456
rect 7392 70446 7420 73034
rect 7477 72924 7785 72944
rect 7477 72922 7483 72924
rect 7539 72922 7563 72924
rect 7619 72922 7643 72924
rect 7699 72922 7723 72924
rect 7779 72922 7785 72924
rect 7539 72870 7541 72922
rect 7721 72870 7723 72922
rect 7477 72868 7483 72870
rect 7539 72868 7563 72870
rect 7619 72868 7643 72870
rect 7699 72868 7723 72870
rect 7779 72868 7785 72870
rect 7477 72848 7785 72868
rect 8312 72826 8340 76366
rect 8404 74458 8432 76978
rect 8484 75948 8536 75954
rect 8484 75890 8536 75896
rect 8392 74452 8444 74458
rect 8392 74394 8444 74400
rect 8300 72820 8352 72826
rect 8300 72762 8352 72768
rect 8496 72486 8524 75890
rect 8956 74390 8984 77454
rect 9312 77376 9364 77382
rect 9310 77344 9312 77353
rect 9364 77344 9366 77353
rect 9310 77279 9366 77288
rect 9109 76732 9417 76752
rect 9109 76730 9115 76732
rect 9171 76730 9195 76732
rect 9251 76730 9275 76732
rect 9331 76730 9355 76732
rect 9411 76730 9417 76732
rect 9171 76678 9173 76730
rect 9353 76678 9355 76730
rect 9109 76676 9115 76678
rect 9171 76676 9195 76678
rect 9251 76676 9275 76678
rect 9331 76676 9355 76678
rect 9411 76676 9417 76678
rect 9109 76656 9417 76676
rect 9508 76634 9536 78639
rect 9586 77752 9642 77761
rect 9586 77687 9642 77696
rect 9600 77178 9628 77687
rect 10140 77376 10192 77382
rect 10140 77318 10192 77324
rect 9588 77172 9640 77178
rect 9588 77114 9640 77120
rect 10048 76832 10100 76838
rect 10152 76809 10180 77318
rect 10048 76774 10100 76780
rect 10138 76800 10194 76809
rect 9496 76628 9548 76634
rect 9496 76570 9548 76576
rect 10060 76401 10088 76774
rect 10138 76735 10194 76744
rect 10046 76392 10102 76401
rect 10046 76327 10102 76336
rect 10048 76288 10100 76294
rect 10048 76230 10100 76236
rect 9312 76084 9364 76090
rect 9312 76026 9364 76032
rect 9324 75857 9352 76026
rect 9864 75948 9916 75954
rect 9864 75890 9916 75896
rect 9310 75848 9366 75857
rect 9310 75783 9366 75792
rect 9109 75644 9417 75664
rect 9109 75642 9115 75644
rect 9171 75642 9195 75644
rect 9251 75642 9275 75644
rect 9331 75642 9355 75644
rect 9411 75642 9417 75644
rect 9171 75590 9173 75642
rect 9353 75590 9355 75642
rect 9109 75588 9115 75590
rect 9171 75588 9195 75590
rect 9251 75588 9275 75590
rect 9331 75588 9355 75590
rect 9411 75588 9417 75590
rect 9109 75568 9417 75588
rect 9109 74556 9417 74576
rect 9109 74554 9115 74556
rect 9171 74554 9195 74556
rect 9251 74554 9275 74556
rect 9331 74554 9355 74556
rect 9411 74554 9417 74556
rect 9171 74502 9173 74554
rect 9353 74502 9355 74554
rect 9109 74500 9115 74502
rect 9171 74500 9195 74502
rect 9251 74500 9275 74502
rect 9331 74500 9355 74502
rect 9411 74500 9417 74502
rect 9109 74480 9417 74500
rect 8944 74384 8996 74390
rect 8944 74326 8996 74332
rect 8668 73772 8720 73778
rect 8668 73714 8720 73720
rect 8576 73024 8628 73030
rect 8576 72966 8628 72972
rect 8484 72480 8536 72486
rect 8484 72422 8536 72428
rect 8588 71913 8616 72966
rect 8574 71904 8630 71913
rect 7477 71836 7785 71856
rect 8574 71839 8630 71848
rect 7477 71834 7483 71836
rect 7539 71834 7563 71836
rect 7619 71834 7643 71836
rect 7699 71834 7723 71836
rect 7779 71834 7785 71836
rect 7539 71782 7541 71834
rect 7721 71782 7723 71834
rect 7477 71780 7483 71782
rect 7539 71780 7563 71782
rect 7619 71780 7643 71782
rect 7699 71780 7723 71782
rect 7779 71780 7785 71782
rect 7477 71760 7785 71780
rect 7932 71052 7984 71058
rect 7932 70994 7984 71000
rect 7477 70748 7785 70768
rect 7477 70746 7483 70748
rect 7539 70746 7563 70748
rect 7619 70746 7643 70748
rect 7699 70746 7723 70748
rect 7779 70746 7785 70748
rect 7539 70694 7541 70746
rect 7721 70694 7723 70746
rect 7477 70692 7483 70694
rect 7539 70692 7563 70694
rect 7619 70692 7643 70694
rect 7699 70692 7723 70694
rect 7779 70692 7785 70694
rect 7477 70672 7785 70692
rect 7944 70514 7972 70994
rect 7932 70508 7984 70514
rect 7932 70450 7984 70456
rect 7380 70440 7432 70446
rect 7300 70388 7380 70394
rect 7300 70382 7432 70388
rect 7840 70440 7892 70446
rect 7840 70382 7892 70388
rect 7300 70366 7420 70382
rect 7196 70032 7248 70038
rect 7196 69974 7248 69980
rect 7208 68814 7236 69974
rect 7196 68808 7248 68814
rect 7196 68750 7248 68756
rect 7208 66638 7236 68750
rect 7196 66632 7248 66638
rect 7196 66574 7248 66580
rect 7104 62280 7156 62286
rect 7104 62222 7156 62228
rect 7116 60734 7144 62222
rect 7116 60706 7236 60734
rect 7104 60240 7156 60246
rect 7104 60182 7156 60188
rect 7010 51232 7066 51241
rect 7010 51167 7066 51176
rect 7010 51096 7066 51105
rect 7010 51031 7012 51040
rect 7064 51031 7066 51040
rect 7012 51002 7064 51008
rect 7010 50960 7066 50969
rect 7010 50895 7066 50904
rect 7024 49706 7052 50895
rect 7012 49700 7064 49706
rect 7012 49642 7064 49648
rect 7010 49600 7066 49609
rect 7010 49535 7066 49544
rect 7024 46170 7052 49535
rect 7116 46186 7144 60182
rect 7208 59974 7236 60706
rect 7196 59968 7248 59974
rect 7196 59910 7248 59916
rect 7196 59764 7248 59770
rect 7196 59706 7248 59712
rect 7208 51513 7236 59706
rect 7194 51504 7250 51513
rect 7194 51439 7250 51448
rect 7300 51066 7328 70366
rect 7477 69660 7785 69680
rect 7477 69658 7483 69660
rect 7539 69658 7563 69660
rect 7619 69658 7643 69660
rect 7699 69658 7723 69660
rect 7779 69658 7785 69660
rect 7539 69606 7541 69658
rect 7721 69606 7723 69658
rect 7477 69604 7483 69606
rect 7539 69604 7563 69606
rect 7619 69604 7643 69606
rect 7699 69604 7723 69606
rect 7779 69604 7785 69606
rect 7477 69584 7785 69604
rect 7477 68572 7785 68592
rect 7477 68570 7483 68572
rect 7539 68570 7563 68572
rect 7619 68570 7643 68572
rect 7699 68570 7723 68572
rect 7779 68570 7785 68572
rect 7539 68518 7541 68570
rect 7721 68518 7723 68570
rect 7477 68516 7483 68518
rect 7539 68516 7563 68518
rect 7619 68516 7643 68518
rect 7699 68516 7723 68518
rect 7779 68516 7785 68518
rect 7477 68496 7785 68516
rect 7477 67484 7785 67504
rect 7477 67482 7483 67484
rect 7539 67482 7563 67484
rect 7619 67482 7643 67484
rect 7699 67482 7723 67484
rect 7779 67482 7785 67484
rect 7539 67430 7541 67482
rect 7721 67430 7723 67482
rect 7477 67428 7483 67430
rect 7539 67428 7563 67430
rect 7619 67428 7643 67430
rect 7699 67428 7723 67430
rect 7779 67428 7785 67430
rect 7477 67408 7785 67428
rect 7380 67040 7432 67046
rect 7380 66982 7432 66988
rect 7392 65210 7420 66982
rect 7477 66396 7785 66416
rect 7477 66394 7483 66396
rect 7539 66394 7563 66396
rect 7619 66394 7643 66396
rect 7699 66394 7723 66396
rect 7779 66394 7785 66396
rect 7539 66342 7541 66394
rect 7721 66342 7723 66394
rect 7477 66340 7483 66342
rect 7539 66340 7563 66342
rect 7619 66340 7643 66342
rect 7699 66340 7723 66342
rect 7779 66340 7785 66342
rect 7477 66320 7785 66340
rect 7477 65308 7785 65328
rect 7477 65306 7483 65308
rect 7539 65306 7563 65308
rect 7619 65306 7643 65308
rect 7699 65306 7723 65308
rect 7779 65306 7785 65308
rect 7539 65254 7541 65306
rect 7721 65254 7723 65306
rect 7477 65252 7483 65254
rect 7539 65252 7563 65254
rect 7619 65252 7643 65254
rect 7699 65252 7723 65254
rect 7779 65252 7785 65254
rect 7477 65232 7785 65252
rect 7380 65204 7432 65210
rect 7380 65146 7432 65152
rect 7392 63034 7420 65146
rect 7477 64220 7785 64240
rect 7477 64218 7483 64220
rect 7539 64218 7563 64220
rect 7619 64218 7643 64220
rect 7699 64218 7723 64220
rect 7779 64218 7785 64220
rect 7539 64166 7541 64218
rect 7721 64166 7723 64218
rect 7477 64164 7483 64166
rect 7539 64164 7563 64166
rect 7619 64164 7643 64166
rect 7699 64164 7723 64166
rect 7779 64164 7785 64166
rect 7477 64144 7785 64164
rect 7477 63132 7785 63152
rect 7477 63130 7483 63132
rect 7539 63130 7563 63132
rect 7619 63130 7643 63132
rect 7699 63130 7723 63132
rect 7779 63130 7785 63132
rect 7539 63078 7541 63130
rect 7721 63078 7723 63130
rect 7477 63076 7483 63078
rect 7539 63076 7563 63078
rect 7619 63076 7643 63078
rect 7699 63076 7723 63078
rect 7779 63076 7785 63078
rect 7477 63056 7785 63076
rect 7380 63028 7432 63034
rect 7380 62970 7432 62976
rect 7380 62688 7432 62694
rect 7380 62630 7432 62636
rect 7392 51066 7420 62630
rect 7477 62044 7785 62064
rect 7477 62042 7483 62044
rect 7539 62042 7563 62044
rect 7619 62042 7643 62044
rect 7699 62042 7723 62044
rect 7779 62042 7785 62044
rect 7539 61990 7541 62042
rect 7721 61990 7723 62042
rect 7477 61988 7483 61990
rect 7539 61988 7563 61990
rect 7619 61988 7643 61990
rect 7699 61988 7723 61990
rect 7779 61988 7785 61990
rect 7477 61968 7785 61988
rect 7477 60956 7785 60976
rect 7477 60954 7483 60956
rect 7539 60954 7563 60956
rect 7619 60954 7643 60956
rect 7699 60954 7723 60956
rect 7779 60954 7785 60956
rect 7539 60902 7541 60954
rect 7721 60902 7723 60954
rect 7477 60900 7483 60902
rect 7539 60900 7563 60902
rect 7619 60900 7643 60902
rect 7699 60900 7723 60902
rect 7779 60900 7785 60902
rect 7477 60880 7785 60900
rect 7477 59868 7785 59888
rect 7477 59866 7483 59868
rect 7539 59866 7563 59868
rect 7619 59866 7643 59868
rect 7699 59866 7723 59868
rect 7779 59866 7785 59868
rect 7539 59814 7541 59866
rect 7721 59814 7723 59866
rect 7477 59812 7483 59814
rect 7539 59812 7563 59814
rect 7619 59812 7643 59814
rect 7699 59812 7723 59814
rect 7779 59812 7785 59814
rect 7477 59792 7785 59812
rect 7477 58780 7785 58800
rect 7477 58778 7483 58780
rect 7539 58778 7563 58780
rect 7619 58778 7643 58780
rect 7699 58778 7723 58780
rect 7779 58778 7785 58780
rect 7539 58726 7541 58778
rect 7721 58726 7723 58778
rect 7477 58724 7483 58726
rect 7539 58724 7563 58726
rect 7619 58724 7643 58726
rect 7699 58724 7723 58726
rect 7779 58724 7785 58726
rect 7477 58704 7785 58724
rect 7477 57692 7785 57712
rect 7477 57690 7483 57692
rect 7539 57690 7563 57692
rect 7619 57690 7643 57692
rect 7699 57690 7723 57692
rect 7779 57690 7785 57692
rect 7539 57638 7541 57690
rect 7721 57638 7723 57690
rect 7477 57636 7483 57638
rect 7539 57636 7563 57638
rect 7619 57636 7643 57638
rect 7699 57636 7723 57638
rect 7779 57636 7785 57638
rect 7477 57616 7785 57636
rect 7477 56604 7785 56624
rect 7477 56602 7483 56604
rect 7539 56602 7563 56604
rect 7619 56602 7643 56604
rect 7699 56602 7723 56604
rect 7779 56602 7785 56604
rect 7539 56550 7541 56602
rect 7721 56550 7723 56602
rect 7477 56548 7483 56550
rect 7539 56548 7563 56550
rect 7619 56548 7643 56550
rect 7699 56548 7723 56550
rect 7779 56548 7785 56550
rect 7477 56528 7785 56548
rect 7748 56160 7800 56166
rect 7748 56102 7800 56108
rect 7760 55706 7788 56102
rect 7852 55842 7880 70382
rect 7944 68882 7972 70450
rect 8392 69420 8444 69426
rect 8392 69362 8444 69368
rect 7932 68876 7984 68882
rect 7932 68818 7984 68824
rect 8206 68776 8262 68785
rect 7932 68740 7984 68746
rect 8206 68711 8262 68720
rect 7932 68682 7984 68688
rect 7944 55978 7972 68682
rect 8220 68678 8248 68711
rect 8208 68672 8260 68678
rect 8208 68614 8260 68620
rect 8208 68332 8260 68338
rect 8208 68274 8260 68280
rect 8024 66564 8076 66570
rect 8024 66506 8076 66512
rect 8036 56166 8064 66506
rect 8116 65068 8168 65074
rect 8116 65010 8168 65016
rect 8128 62762 8156 65010
rect 8116 62756 8168 62762
rect 8116 62698 8168 62704
rect 8128 60858 8156 62698
rect 8220 62234 8248 68274
rect 8300 67584 8352 67590
rect 8300 67526 8352 67532
rect 8312 67425 8340 67526
rect 8298 67416 8354 67425
rect 8404 67386 8432 69362
rect 8576 68672 8628 68678
rect 8576 68614 8628 68620
rect 8298 67351 8354 67360
rect 8392 67380 8444 67386
rect 8392 67322 8444 67328
rect 8300 67244 8352 67250
rect 8300 67186 8352 67192
rect 8312 66337 8340 67186
rect 8298 66328 8354 66337
rect 8298 66263 8354 66272
rect 8392 64456 8444 64462
rect 8392 64398 8444 64404
rect 8220 62206 8340 62234
rect 8208 62144 8260 62150
rect 8208 62086 8260 62092
rect 8116 60852 8168 60858
rect 8116 60794 8168 60800
rect 8114 60752 8170 60761
rect 8114 60687 8170 60696
rect 8024 56160 8076 56166
rect 8024 56102 8076 56108
rect 7944 55950 8064 55978
rect 7852 55814 7972 55842
rect 7760 55678 7880 55706
rect 7477 55516 7785 55536
rect 7477 55514 7483 55516
rect 7539 55514 7563 55516
rect 7619 55514 7643 55516
rect 7699 55514 7723 55516
rect 7779 55514 7785 55516
rect 7539 55462 7541 55514
rect 7721 55462 7723 55514
rect 7477 55460 7483 55462
rect 7539 55460 7563 55462
rect 7619 55460 7643 55462
rect 7699 55460 7723 55462
rect 7779 55460 7785 55462
rect 7477 55440 7785 55460
rect 7477 54428 7785 54448
rect 7477 54426 7483 54428
rect 7539 54426 7563 54428
rect 7619 54426 7643 54428
rect 7699 54426 7723 54428
rect 7779 54426 7785 54428
rect 7539 54374 7541 54426
rect 7721 54374 7723 54426
rect 7477 54372 7483 54374
rect 7539 54372 7563 54374
rect 7619 54372 7643 54374
rect 7699 54372 7723 54374
rect 7779 54372 7785 54374
rect 7477 54352 7785 54372
rect 7477 53340 7785 53360
rect 7477 53338 7483 53340
rect 7539 53338 7563 53340
rect 7619 53338 7643 53340
rect 7699 53338 7723 53340
rect 7779 53338 7785 53340
rect 7539 53286 7541 53338
rect 7721 53286 7723 53338
rect 7477 53284 7483 53286
rect 7539 53284 7563 53286
rect 7619 53284 7643 53286
rect 7699 53284 7723 53286
rect 7779 53284 7785 53286
rect 7477 53264 7785 53284
rect 7477 52252 7785 52272
rect 7477 52250 7483 52252
rect 7539 52250 7563 52252
rect 7619 52250 7643 52252
rect 7699 52250 7723 52252
rect 7779 52250 7785 52252
rect 7539 52198 7541 52250
rect 7721 52198 7723 52250
rect 7477 52196 7483 52198
rect 7539 52196 7563 52198
rect 7619 52196 7643 52198
rect 7699 52196 7723 52198
rect 7779 52196 7785 52198
rect 7477 52176 7785 52196
rect 7477 51164 7785 51184
rect 7477 51162 7483 51164
rect 7539 51162 7563 51164
rect 7619 51162 7643 51164
rect 7699 51162 7723 51164
rect 7779 51162 7785 51164
rect 7539 51110 7541 51162
rect 7721 51110 7723 51162
rect 7477 51108 7483 51110
rect 7539 51108 7563 51110
rect 7619 51108 7643 51110
rect 7699 51108 7723 51110
rect 7779 51108 7785 51110
rect 7477 51088 7785 51108
rect 7288 51060 7340 51066
rect 7288 51002 7340 51008
rect 7380 51060 7432 51066
rect 7380 51002 7432 51008
rect 7196 50856 7248 50862
rect 7196 50798 7248 50804
rect 7288 50856 7340 50862
rect 7288 50798 7340 50804
rect 7380 50856 7432 50862
rect 7380 50798 7432 50804
rect 7208 49638 7236 50798
rect 7196 49632 7248 49638
rect 7196 49574 7248 49580
rect 7196 49292 7248 49298
rect 7196 49234 7248 49240
rect 7208 46345 7236 49234
rect 7194 46336 7250 46345
rect 7194 46271 7250 46280
rect 7012 46164 7064 46170
rect 7116 46158 7236 46186
rect 7012 46106 7064 46112
rect 6932 46022 7144 46050
rect 6920 45960 6972 45966
rect 6920 45902 6972 45908
rect 7012 45960 7064 45966
rect 7012 45902 7064 45908
rect 6932 43450 6960 45902
rect 6920 43444 6972 43450
rect 6920 43386 6972 43392
rect 6828 42900 6880 42906
rect 6828 42842 6880 42848
rect 6826 42800 6882 42809
rect 6826 42735 6828 42744
rect 6880 42735 6882 42744
rect 6920 42764 6972 42770
rect 6828 42706 6880 42712
rect 6920 42706 6972 42712
rect 6932 42673 6960 42706
rect 6918 42664 6974 42673
rect 6918 42599 6974 42608
rect 6920 42560 6972 42566
rect 6840 42508 6920 42514
rect 6840 42502 6972 42508
rect 6840 42486 6960 42502
rect 6840 41138 6868 42486
rect 6920 42288 6972 42294
rect 6920 42230 6972 42236
rect 6932 41478 6960 42230
rect 6920 41472 6972 41478
rect 6920 41414 6972 41420
rect 6828 41132 6880 41138
rect 6828 41074 6880 41080
rect 6828 40996 6880 41002
rect 6828 40938 6880 40944
rect 6840 39386 6868 40938
rect 6920 40928 6972 40934
rect 6920 40870 6972 40876
rect 6932 39522 6960 40870
rect 7024 39642 7052 45902
rect 7012 39636 7064 39642
rect 7012 39578 7064 39584
rect 6932 39494 7052 39522
rect 6840 39358 6960 39386
rect 6828 39024 6880 39030
rect 6828 38966 6880 38972
rect 6840 28994 6868 38966
rect 6932 38332 6960 39358
rect 7024 38457 7052 39494
rect 7116 38554 7144 46022
rect 7208 41002 7236 46158
rect 7300 45286 7328 50798
rect 7288 45280 7340 45286
rect 7288 45222 7340 45228
rect 7288 44736 7340 44742
rect 7288 44678 7340 44684
rect 7300 43897 7328 44678
rect 7286 43888 7342 43897
rect 7286 43823 7342 43832
rect 7288 43648 7340 43654
rect 7288 43590 7340 43596
rect 7196 40996 7248 41002
rect 7196 40938 7248 40944
rect 7196 40724 7248 40730
rect 7196 40666 7248 40672
rect 7104 38548 7156 38554
rect 7104 38490 7156 38496
rect 7010 38448 7066 38457
rect 7010 38383 7066 38392
rect 6932 38304 7144 38332
rect 7010 38176 7066 38185
rect 7010 38111 7066 38120
rect 6920 37256 6972 37262
rect 6920 37198 6972 37204
rect 6932 36718 6960 37198
rect 6920 36712 6972 36718
rect 6920 36654 6972 36660
rect 7024 32910 7052 38111
rect 7116 33998 7144 38304
rect 7208 35698 7236 40666
rect 7196 35692 7248 35698
rect 7196 35634 7248 35640
rect 7196 35556 7248 35562
rect 7196 35498 7248 35504
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 7012 32904 7064 32910
rect 7012 32846 7064 32852
rect 7104 32836 7156 32842
rect 7104 32778 7156 32784
rect 6840 28966 7052 28994
rect 7024 27470 7052 28966
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 6736 26036 6788 26042
rect 6736 25978 6788 25984
rect 7116 24818 7144 32778
rect 7208 28558 7236 35498
rect 7300 29170 7328 43590
rect 7392 30734 7420 50798
rect 7477 50076 7785 50096
rect 7477 50074 7483 50076
rect 7539 50074 7563 50076
rect 7619 50074 7643 50076
rect 7699 50074 7723 50076
rect 7779 50074 7785 50076
rect 7539 50022 7541 50074
rect 7721 50022 7723 50074
rect 7477 50020 7483 50022
rect 7539 50020 7563 50022
rect 7619 50020 7643 50022
rect 7699 50020 7723 50022
rect 7779 50020 7785 50022
rect 7477 50000 7785 50020
rect 7477 48988 7785 49008
rect 7477 48986 7483 48988
rect 7539 48986 7563 48988
rect 7619 48986 7643 48988
rect 7699 48986 7723 48988
rect 7779 48986 7785 48988
rect 7539 48934 7541 48986
rect 7721 48934 7723 48986
rect 7477 48932 7483 48934
rect 7539 48932 7563 48934
rect 7619 48932 7643 48934
rect 7699 48932 7723 48934
rect 7779 48932 7785 48934
rect 7477 48912 7785 48932
rect 7746 48784 7802 48793
rect 7746 48719 7802 48728
rect 7760 48113 7788 48719
rect 7746 48104 7802 48113
rect 7746 48039 7802 48048
rect 7477 47900 7785 47920
rect 7477 47898 7483 47900
rect 7539 47898 7563 47900
rect 7619 47898 7643 47900
rect 7699 47898 7723 47900
rect 7779 47898 7785 47900
rect 7539 47846 7541 47898
rect 7721 47846 7723 47898
rect 7477 47844 7483 47846
rect 7539 47844 7563 47846
rect 7619 47844 7643 47846
rect 7699 47844 7723 47846
rect 7779 47844 7785 47846
rect 7477 47824 7785 47844
rect 7477 46812 7785 46832
rect 7477 46810 7483 46812
rect 7539 46810 7563 46812
rect 7619 46810 7643 46812
rect 7699 46810 7723 46812
rect 7779 46810 7785 46812
rect 7539 46758 7541 46810
rect 7721 46758 7723 46810
rect 7477 46756 7483 46758
rect 7539 46756 7563 46758
rect 7619 46756 7643 46758
rect 7699 46756 7723 46758
rect 7779 46756 7785 46758
rect 7477 46736 7785 46756
rect 7477 45724 7785 45744
rect 7477 45722 7483 45724
rect 7539 45722 7563 45724
rect 7619 45722 7643 45724
rect 7699 45722 7723 45724
rect 7779 45722 7785 45724
rect 7539 45670 7541 45722
rect 7721 45670 7723 45722
rect 7477 45668 7483 45670
rect 7539 45668 7563 45670
rect 7619 45668 7643 45670
rect 7699 45668 7723 45670
rect 7779 45668 7785 45670
rect 7477 45648 7785 45668
rect 7477 44636 7785 44656
rect 7477 44634 7483 44636
rect 7539 44634 7563 44636
rect 7619 44634 7643 44636
rect 7699 44634 7723 44636
rect 7779 44634 7785 44636
rect 7539 44582 7541 44634
rect 7721 44582 7723 44634
rect 7477 44580 7483 44582
rect 7539 44580 7563 44582
rect 7619 44580 7643 44582
rect 7699 44580 7723 44582
rect 7779 44580 7785 44582
rect 7477 44560 7785 44580
rect 7562 44296 7618 44305
rect 7562 44231 7618 44240
rect 7576 43994 7604 44231
rect 7564 43988 7616 43994
rect 7564 43930 7616 43936
rect 7477 43548 7785 43568
rect 7477 43546 7483 43548
rect 7539 43546 7563 43548
rect 7619 43546 7643 43548
rect 7699 43546 7723 43548
rect 7779 43546 7785 43548
rect 7539 43494 7541 43546
rect 7721 43494 7723 43546
rect 7477 43492 7483 43494
rect 7539 43492 7563 43494
rect 7619 43492 7643 43494
rect 7699 43492 7723 43494
rect 7779 43492 7785 43494
rect 7477 43472 7785 43492
rect 7477 42460 7785 42480
rect 7477 42458 7483 42460
rect 7539 42458 7563 42460
rect 7619 42458 7643 42460
rect 7699 42458 7723 42460
rect 7779 42458 7785 42460
rect 7539 42406 7541 42458
rect 7721 42406 7723 42458
rect 7477 42404 7483 42406
rect 7539 42404 7563 42406
rect 7619 42404 7643 42406
rect 7699 42404 7723 42406
rect 7779 42404 7785 42406
rect 7477 42384 7785 42404
rect 7477 41372 7785 41392
rect 7477 41370 7483 41372
rect 7539 41370 7563 41372
rect 7619 41370 7643 41372
rect 7699 41370 7723 41372
rect 7779 41370 7785 41372
rect 7539 41318 7541 41370
rect 7721 41318 7723 41370
rect 7477 41316 7483 41318
rect 7539 41316 7563 41318
rect 7619 41316 7643 41318
rect 7699 41316 7723 41318
rect 7779 41316 7785 41318
rect 7477 41296 7785 41316
rect 7472 41200 7524 41206
rect 7472 41142 7524 41148
rect 7484 40458 7512 41142
rect 7852 40934 7880 55678
rect 7840 40928 7892 40934
rect 7840 40870 7892 40876
rect 7944 40730 7972 55814
rect 8036 46442 8064 55950
rect 8128 51074 8156 60687
rect 8220 60178 8248 62086
rect 8312 61033 8340 62206
rect 8298 61024 8354 61033
rect 8298 60959 8354 60968
rect 8300 60852 8352 60858
rect 8300 60794 8352 60800
rect 8208 60172 8260 60178
rect 8208 60114 8260 60120
rect 8220 59770 8248 60114
rect 8208 59764 8260 59770
rect 8208 59706 8260 59712
rect 8312 59650 8340 60794
rect 8220 59622 8340 59650
rect 8220 51270 8248 59622
rect 8300 58676 8352 58682
rect 8300 58618 8352 58624
rect 8312 51377 8340 58618
rect 8298 51368 8354 51377
rect 8298 51303 8354 51312
rect 8208 51264 8260 51270
rect 8208 51206 8260 51212
rect 8298 51232 8354 51241
rect 8298 51167 8354 51176
rect 8128 51046 8248 51074
rect 8312 51066 8340 51167
rect 8116 50312 8168 50318
rect 8114 50280 8116 50289
rect 8168 50280 8170 50289
rect 8114 50215 8170 50224
rect 8220 49314 8248 51046
rect 8300 51060 8352 51066
rect 8300 51002 8352 51008
rect 8300 50924 8352 50930
rect 8300 50866 8352 50872
rect 8128 49286 8248 49314
rect 8128 46730 8156 49286
rect 8208 49224 8260 49230
rect 8208 49166 8260 49172
rect 8220 48929 8248 49166
rect 8206 48920 8262 48929
rect 8206 48855 8262 48864
rect 8208 48748 8260 48754
rect 8208 48690 8260 48696
rect 8220 48657 8248 48690
rect 8206 48648 8262 48657
rect 8206 48583 8262 48592
rect 8208 48136 8260 48142
rect 8208 48078 8260 48084
rect 8220 47977 8248 48078
rect 8206 47968 8262 47977
rect 8206 47903 8262 47912
rect 8208 47048 8260 47054
rect 8206 47016 8208 47025
rect 8260 47016 8262 47025
rect 8206 46951 8262 46960
rect 8128 46702 8248 46730
rect 8116 46640 8168 46646
rect 8116 46582 8168 46588
rect 8024 46436 8076 46442
rect 8024 46378 8076 46384
rect 8022 46336 8078 46345
rect 8022 46271 8078 46280
rect 7932 40724 7984 40730
rect 7932 40666 7984 40672
rect 8036 40610 8064 46271
rect 8128 43790 8156 46582
rect 8220 45966 8248 46702
rect 8208 45960 8260 45966
rect 8208 45902 8260 45908
rect 8208 45484 8260 45490
rect 8208 45426 8260 45432
rect 8220 44713 8248 45426
rect 8206 44704 8262 44713
rect 8206 44639 8262 44648
rect 8208 44464 8260 44470
rect 8208 44406 8260 44412
rect 8220 43858 8248 44406
rect 8208 43852 8260 43858
rect 8208 43794 8260 43800
rect 8116 43784 8168 43790
rect 8116 43726 8168 43732
rect 7852 40582 8064 40610
rect 7472 40452 7524 40458
rect 7472 40394 7524 40400
rect 7477 40284 7785 40304
rect 7477 40282 7483 40284
rect 7539 40282 7563 40284
rect 7619 40282 7643 40284
rect 7699 40282 7723 40284
rect 7779 40282 7785 40284
rect 7539 40230 7541 40282
rect 7721 40230 7723 40282
rect 7477 40228 7483 40230
rect 7539 40228 7563 40230
rect 7619 40228 7643 40230
rect 7699 40228 7723 40230
rect 7779 40228 7785 40230
rect 7477 40208 7785 40228
rect 7472 39908 7524 39914
rect 7472 39850 7524 39856
rect 7484 39409 7512 39850
rect 7470 39400 7526 39409
rect 7470 39335 7526 39344
rect 7477 39196 7785 39216
rect 7477 39194 7483 39196
rect 7539 39194 7563 39196
rect 7619 39194 7643 39196
rect 7699 39194 7723 39196
rect 7779 39194 7785 39196
rect 7539 39142 7541 39194
rect 7721 39142 7723 39194
rect 7477 39140 7483 39142
rect 7539 39140 7563 39142
rect 7619 39140 7643 39142
rect 7699 39140 7723 39142
rect 7779 39140 7785 39142
rect 7477 39120 7785 39140
rect 7748 38412 7800 38418
rect 7748 38354 7800 38360
rect 7760 38321 7788 38354
rect 7746 38312 7802 38321
rect 7746 38247 7802 38256
rect 7477 38108 7785 38128
rect 7477 38106 7483 38108
rect 7539 38106 7563 38108
rect 7619 38106 7643 38108
rect 7699 38106 7723 38108
rect 7779 38106 7785 38108
rect 7539 38054 7541 38106
rect 7721 38054 7723 38106
rect 7477 38052 7483 38054
rect 7539 38052 7563 38054
rect 7619 38052 7643 38054
rect 7699 38052 7723 38054
rect 7779 38052 7785 38054
rect 7477 38032 7785 38052
rect 7748 37732 7800 37738
rect 7748 37674 7800 37680
rect 7760 37466 7788 37674
rect 7748 37460 7800 37466
rect 7748 37402 7800 37408
rect 7477 37020 7785 37040
rect 7477 37018 7483 37020
rect 7539 37018 7563 37020
rect 7619 37018 7643 37020
rect 7699 37018 7723 37020
rect 7779 37018 7785 37020
rect 7539 36966 7541 37018
rect 7721 36966 7723 37018
rect 7477 36964 7483 36966
rect 7539 36964 7563 36966
rect 7619 36964 7643 36966
rect 7699 36964 7723 36966
rect 7779 36964 7785 36966
rect 7477 36944 7785 36964
rect 7852 36310 7880 40582
rect 7932 40452 7984 40458
rect 7932 40394 7984 40400
rect 7840 36304 7892 36310
rect 7840 36246 7892 36252
rect 7477 35932 7785 35952
rect 7477 35930 7483 35932
rect 7539 35930 7563 35932
rect 7619 35930 7643 35932
rect 7699 35930 7723 35932
rect 7779 35930 7785 35932
rect 7539 35878 7541 35930
rect 7721 35878 7723 35930
rect 7477 35876 7483 35878
rect 7539 35876 7563 35878
rect 7619 35876 7643 35878
rect 7699 35876 7723 35878
rect 7779 35876 7785 35878
rect 7477 35856 7785 35876
rect 7477 34844 7785 34864
rect 7477 34842 7483 34844
rect 7539 34842 7563 34844
rect 7619 34842 7643 34844
rect 7699 34842 7723 34844
rect 7779 34842 7785 34844
rect 7539 34790 7541 34842
rect 7721 34790 7723 34842
rect 7477 34788 7483 34790
rect 7539 34788 7563 34790
rect 7619 34788 7643 34790
rect 7699 34788 7723 34790
rect 7779 34788 7785 34790
rect 7477 34768 7785 34788
rect 7840 34536 7892 34542
rect 7840 34478 7892 34484
rect 7477 33756 7785 33776
rect 7477 33754 7483 33756
rect 7539 33754 7563 33756
rect 7619 33754 7643 33756
rect 7699 33754 7723 33756
rect 7779 33754 7785 33756
rect 7539 33702 7541 33754
rect 7721 33702 7723 33754
rect 7477 33700 7483 33702
rect 7539 33700 7563 33702
rect 7619 33700 7643 33702
rect 7699 33700 7723 33702
rect 7779 33700 7785 33702
rect 7477 33680 7785 33700
rect 7477 32668 7785 32688
rect 7477 32666 7483 32668
rect 7539 32666 7563 32668
rect 7619 32666 7643 32668
rect 7699 32666 7723 32668
rect 7779 32666 7785 32668
rect 7539 32614 7541 32666
rect 7721 32614 7723 32666
rect 7477 32612 7483 32614
rect 7539 32612 7563 32614
rect 7619 32612 7643 32614
rect 7699 32612 7723 32614
rect 7779 32612 7785 32614
rect 7477 32592 7785 32612
rect 7477 31580 7785 31600
rect 7477 31578 7483 31580
rect 7539 31578 7563 31580
rect 7619 31578 7643 31580
rect 7699 31578 7723 31580
rect 7779 31578 7785 31580
rect 7539 31526 7541 31578
rect 7721 31526 7723 31578
rect 7477 31524 7483 31526
rect 7539 31524 7563 31526
rect 7619 31524 7643 31526
rect 7699 31524 7723 31526
rect 7779 31524 7785 31526
rect 7477 31504 7785 31524
rect 7380 30728 7432 30734
rect 7380 30670 7432 30676
rect 7477 30492 7785 30512
rect 7477 30490 7483 30492
rect 7539 30490 7563 30492
rect 7619 30490 7643 30492
rect 7699 30490 7723 30492
rect 7779 30490 7785 30492
rect 7539 30438 7541 30490
rect 7721 30438 7723 30490
rect 7477 30436 7483 30438
rect 7539 30436 7563 30438
rect 7619 30436 7643 30438
rect 7699 30436 7723 30438
rect 7779 30436 7785 30438
rect 7477 30416 7785 30436
rect 7477 29404 7785 29424
rect 7477 29402 7483 29404
rect 7539 29402 7563 29404
rect 7619 29402 7643 29404
rect 7699 29402 7723 29404
rect 7779 29402 7785 29404
rect 7539 29350 7541 29402
rect 7721 29350 7723 29402
rect 7477 29348 7483 29350
rect 7539 29348 7563 29350
rect 7619 29348 7643 29350
rect 7699 29348 7723 29350
rect 7779 29348 7785 29350
rect 7477 29328 7785 29348
rect 7380 29300 7432 29306
rect 7380 29242 7432 29248
rect 7288 29164 7340 29170
rect 7288 29106 7340 29112
rect 7288 29028 7340 29034
rect 7288 28970 7340 28976
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 6736 23588 6788 23594
rect 6736 23530 6788 23536
rect 6564 22066 6684 22094
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6472 17202 6500 17478
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 5845 16892 6153 16912
rect 5845 16890 5851 16892
rect 5907 16890 5931 16892
rect 5987 16890 6011 16892
rect 6067 16890 6091 16892
rect 6147 16890 6153 16892
rect 5907 16838 5909 16890
rect 6089 16838 6091 16890
rect 5845 16836 5851 16838
rect 5907 16836 5931 16838
rect 5987 16836 6011 16838
rect 6067 16836 6091 16838
rect 6147 16836 6153 16838
rect 5845 16816 6153 16836
rect 5845 15804 6153 15824
rect 5845 15802 5851 15804
rect 5907 15802 5931 15804
rect 5987 15802 6011 15804
rect 6067 15802 6091 15804
rect 6147 15802 6153 15804
rect 5907 15750 5909 15802
rect 6089 15750 6091 15802
rect 5845 15748 5851 15750
rect 5907 15748 5931 15750
rect 5987 15748 6011 15750
rect 6067 15748 6091 15750
rect 6147 15748 6153 15750
rect 5845 15728 6153 15748
rect 5845 14716 6153 14736
rect 5845 14714 5851 14716
rect 5907 14714 5931 14716
rect 5987 14714 6011 14716
rect 6067 14714 6091 14716
rect 6147 14714 6153 14716
rect 5907 14662 5909 14714
rect 6089 14662 6091 14714
rect 5845 14660 5851 14662
rect 5907 14660 5931 14662
rect 5987 14660 6011 14662
rect 6067 14660 6091 14662
rect 6147 14660 6153 14662
rect 5845 14640 6153 14660
rect 6182 14512 6238 14521
rect 6182 14447 6238 14456
rect 5845 13628 6153 13648
rect 5845 13626 5851 13628
rect 5907 13626 5931 13628
rect 5987 13626 6011 13628
rect 6067 13626 6091 13628
rect 6147 13626 6153 13628
rect 5907 13574 5909 13626
rect 6089 13574 6091 13626
rect 5845 13572 5851 13574
rect 5907 13572 5931 13574
rect 5987 13572 6011 13574
rect 6067 13572 6091 13574
rect 6147 13572 6153 13574
rect 5845 13552 6153 13572
rect 6196 13512 6224 14447
rect 6288 14278 6316 16934
rect 6366 14784 6422 14793
rect 6366 14719 6422 14728
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6380 14074 6408 14719
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6564 13920 6592 22066
rect 6748 20466 6776 23530
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6932 19378 6960 21286
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7024 17762 7052 19654
rect 7116 18426 7144 22578
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 6932 17734 7052 17762
rect 6932 16454 6960 17734
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7024 16658 7052 17614
rect 7208 17320 7236 26930
rect 7300 18970 7328 28970
rect 7392 21554 7420 29242
rect 7477 28316 7785 28336
rect 7477 28314 7483 28316
rect 7539 28314 7563 28316
rect 7619 28314 7643 28316
rect 7699 28314 7723 28316
rect 7779 28314 7785 28316
rect 7539 28262 7541 28314
rect 7721 28262 7723 28314
rect 7477 28260 7483 28262
rect 7539 28260 7563 28262
rect 7619 28260 7643 28262
rect 7699 28260 7723 28262
rect 7779 28260 7785 28262
rect 7477 28240 7785 28260
rect 7477 27228 7785 27248
rect 7477 27226 7483 27228
rect 7539 27226 7563 27228
rect 7619 27226 7643 27228
rect 7699 27226 7723 27228
rect 7779 27226 7785 27228
rect 7539 27174 7541 27226
rect 7721 27174 7723 27226
rect 7477 27172 7483 27174
rect 7539 27172 7563 27174
rect 7619 27172 7643 27174
rect 7699 27172 7723 27174
rect 7779 27172 7785 27174
rect 7477 27152 7785 27172
rect 7852 26602 7880 34478
rect 7944 26994 7972 40394
rect 8024 40384 8076 40390
rect 8024 40326 8076 40332
rect 8036 39030 8064 40326
rect 8024 39024 8076 39030
rect 8024 38966 8076 38972
rect 8128 38842 8156 43726
rect 8312 43602 8340 50866
rect 8404 50425 8432 64398
rect 8484 62824 8536 62830
rect 8484 62766 8536 62772
rect 8496 62354 8524 62766
rect 8484 62348 8536 62354
rect 8484 62290 8536 62296
rect 8496 60178 8524 62290
rect 8484 60172 8536 60178
rect 8484 60114 8536 60120
rect 8484 59424 8536 59430
rect 8484 59366 8536 59372
rect 8390 50416 8446 50425
rect 8390 50351 8446 50360
rect 8392 50176 8444 50182
rect 8392 50118 8444 50124
rect 8404 44742 8432 50118
rect 8392 44736 8444 44742
rect 8392 44678 8444 44684
rect 8392 44192 8444 44198
rect 8392 44134 8444 44140
rect 8220 43574 8340 43602
rect 8220 42634 8248 43574
rect 8300 43444 8352 43450
rect 8300 43386 8352 43392
rect 8208 42628 8260 42634
rect 8208 42570 8260 42576
rect 8208 42084 8260 42090
rect 8208 42026 8260 42032
rect 8220 40458 8248 42026
rect 8208 40452 8260 40458
rect 8208 40394 8260 40400
rect 8206 40352 8262 40361
rect 8206 40287 8262 40296
rect 8036 38814 8156 38842
rect 8036 37890 8064 38814
rect 8116 38752 8168 38758
rect 8116 38694 8168 38700
rect 8128 38457 8156 38694
rect 8114 38448 8170 38457
rect 8114 38383 8170 38392
rect 8116 38208 8168 38214
rect 8116 38150 8168 38156
rect 8128 38049 8156 38150
rect 8114 38040 8170 38049
rect 8114 37975 8170 37984
rect 8036 37862 8156 37890
rect 8024 37800 8076 37806
rect 8024 37742 8076 37748
rect 8036 36378 8064 37742
rect 8128 37398 8156 37862
rect 8116 37392 8168 37398
rect 8116 37334 8168 37340
rect 8116 37256 8168 37262
rect 8114 37224 8116 37233
rect 8168 37224 8170 37233
rect 8114 37159 8170 37168
rect 8116 37120 8168 37126
rect 8114 37088 8116 37097
rect 8168 37088 8170 37097
rect 8114 37023 8170 37032
rect 8114 36680 8170 36689
rect 8114 36615 8116 36624
rect 8168 36615 8170 36624
rect 8116 36586 8168 36592
rect 8024 36372 8076 36378
rect 8024 36314 8076 36320
rect 8024 36236 8076 36242
rect 8024 36178 8076 36184
rect 8036 34202 8064 36178
rect 8116 35488 8168 35494
rect 8116 35430 8168 35436
rect 8128 35193 8156 35430
rect 8114 35184 8170 35193
rect 8114 35119 8170 35128
rect 8116 35012 8168 35018
rect 8116 34954 8168 34960
rect 8024 34196 8076 34202
rect 8024 34138 8076 34144
rect 8024 33312 8076 33318
rect 8024 33254 8076 33260
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 8036 26738 8064 33254
rect 8128 33114 8156 34954
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 8116 32972 8168 32978
rect 8116 32914 8168 32920
rect 8128 27062 8156 32914
rect 8116 27056 8168 27062
rect 8116 26998 8168 27004
rect 8036 26710 8156 26738
rect 7852 26574 8064 26602
rect 7932 26512 7984 26518
rect 7932 26454 7984 26460
rect 7477 26140 7785 26160
rect 7477 26138 7483 26140
rect 7539 26138 7563 26140
rect 7619 26138 7643 26140
rect 7699 26138 7723 26140
rect 7779 26138 7785 26140
rect 7539 26086 7541 26138
rect 7721 26086 7723 26138
rect 7477 26084 7483 26086
rect 7539 26084 7563 26086
rect 7619 26084 7643 26086
rect 7699 26084 7723 26086
rect 7779 26084 7785 26086
rect 7477 26064 7785 26084
rect 7477 25052 7785 25072
rect 7477 25050 7483 25052
rect 7539 25050 7563 25052
rect 7619 25050 7643 25052
rect 7699 25050 7723 25052
rect 7779 25050 7785 25052
rect 7539 24998 7541 25050
rect 7721 24998 7723 25050
rect 7477 24996 7483 24998
rect 7539 24996 7563 24998
rect 7619 24996 7643 24998
rect 7699 24996 7723 24998
rect 7779 24996 7785 24998
rect 7477 24976 7785 24996
rect 7477 23964 7785 23984
rect 7477 23962 7483 23964
rect 7539 23962 7563 23964
rect 7619 23962 7643 23964
rect 7699 23962 7723 23964
rect 7779 23962 7785 23964
rect 7539 23910 7541 23962
rect 7721 23910 7723 23962
rect 7477 23908 7483 23910
rect 7539 23908 7563 23910
rect 7619 23908 7643 23910
rect 7699 23908 7723 23910
rect 7779 23908 7785 23910
rect 7477 23888 7785 23908
rect 7477 22876 7785 22896
rect 7477 22874 7483 22876
rect 7539 22874 7563 22876
rect 7619 22874 7643 22876
rect 7699 22874 7723 22876
rect 7779 22874 7785 22876
rect 7539 22822 7541 22874
rect 7721 22822 7723 22874
rect 7477 22820 7483 22822
rect 7539 22820 7563 22822
rect 7619 22820 7643 22822
rect 7699 22820 7723 22822
rect 7779 22820 7785 22822
rect 7477 22800 7785 22820
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7477 21788 7785 21808
rect 7477 21786 7483 21788
rect 7539 21786 7563 21788
rect 7619 21786 7643 21788
rect 7699 21786 7723 21788
rect 7779 21786 7785 21788
rect 7539 21734 7541 21786
rect 7721 21734 7723 21786
rect 7477 21732 7483 21734
rect 7539 21732 7563 21734
rect 7619 21732 7643 21734
rect 7699 21732 7723 21734
rect 7779 21732 7785 21734
rect 7477 21712 7785 21732
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7477 20700 7785 20720
rect 7477 20698 7483 20700
rect 7539 20698 7563 20700
rect 7619 20698 7643 20700
rect 7699 20698 7723 20700
rect 7779 20698 7785 20700
rect 7539 20646 7541 20698
rect 7721 20646 7723 20698
rect 7477 20644 7483 20646
rect 7539 20644 7563 20646
rect 7619 20644 7643 20646
rect 7699 20644 7723 20646
rect 7779 20644 7785 20646
rect 7477 20624 7785 20644
rect 7852 19854 7880 22374
rect 7944 20058 7972 26454
rect 8036 20602 8064 26574
rect 8128 26518 8156 26710
rect 8116 26512 8168 26518
rect 8116 26454 8168 26460
rect 8114 21992 8170 22001
rect 8114 21927 8116 21936
rect 8168 21927 8170 21936
rect 8116 21898 8168 21904
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 8128 20369 8156 20402
rect 8114 20360 8170 20369
rect 8114 20295 8170 20304
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 7477 19612 7785 19632
rect 7477 19610 7483 19612
rect 7539 19610 7563 19612
rect 7619 19610 7643 19612
rect 7699 19610 7723 19612
rect 7779 19610 7785 19612
rect 7539 19558 7541 19610
rect 7721 19558 7723 19610
rect 7477 19556 7483 19558
rect 7539 19556 7563 19558
rect 7619 19556 7643 19558
rect 7699 19556 7723 19558
rect 7779 19556 7785 19558
rect 7477 19536 7785 19556
rect 8128 19553 8156 19790
rect 8114 19544 8170 19553
rect 8114 19479 8170 19488
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7477 18524 7785 18544
rect 7477 18522 7483 18524
rect 7539 18522 7563 18524
rect 7619 18522 7643 18524
rect 7699 18522 7723 18524
rect 7779 18522 7785 18524
rect 7539 18470 7541 18522
rect 7721 18470 7723 18522
rect 7477 18468 7483 18470
rect 7539 18468 7563 18470
rect 7619 18468 7643 18470
rect 7699 18468 7723 18470
rect 7779 18468 7785 18470
rect 7477 18448 7785 18468
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7116 17292 7236 17320
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6736 16040 6788 16046
rect 6932 16017 6960 16050
rect 6736 15982 6788 15988
rect 6918 16008 6974 16017
rect 6644 15428 6696 15434
rect 6644 15370 6696 15376
rect 6104 13484 6224 13512
rect 6472 13892 6592 13920
rect 6104 13326 6132 13484
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 5845 12540 6153 12560
rect 5845 12538 5851 12540
rect 5907 12538 5931 12540
rect 5987 12538 6011 12540
rect 6067 12538 6091 12540
rect 6147 12538 6153 12540
rect 5907 12486 5909 12538
rect 6089 12486 6091 12538
rect 5845 12484 5851 12486
rect 5907 12484 5931 12486
rect 5987 12484 6011 12486
rect 6067 12484 6091 12486
rect 6147 12484 6153 12486
rect 5845 12464 6153 12484
rect 6196 12442 6224 13262
rect 6274 13016 6330 13025
rect 6274 12951 6330 12960
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 5816 12232 5868 12238
rect 5908 12232 5960 12238
rect 5816 12174 5868 12180
rect 5906 12200 5908 12209
rect 5960 12200 5962 12209
rect 5828 11898 5856 12174
rect 5906 12135 5962 12144
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5845 11452 6153 11472
rect 5845 11450 5851 11452
rect 5907 11450 5931 11452
rect 5987 11450 6011 11452
rect 6067 11450 6091 11452
rect 6147 11450 6153 11452
rect 5907 11398 5909 11450
rect 6089 11398 6091 11450
rect 5845 11396 5851 11398
rect 5907 11396 5931 11398
rect 5987 11396 6011 11398
rect 6067 11396 6091 11398
rect 6147 11396 6153 11398
rect 5845 11376 6153 11396
rect 5845 10364 6153 10384
rect 5845 10362 5851 10364
rect 5907 10362 5931 10364
rect 5987 10362 6011 10364
rect 6067 10362 6091 10364
rect 6147 10362 6153 10364
rect 5907 10310 5909 10362
rect 6089 10310 6091 10362
rect 5845 10308 5851 10310
rect 5907 10308 5931 10310
rect 5987 10308 6011 10310
rect 6067 10308 6091 10310
rect 6147 10308 6153 10310
rect 5845 10288 6153 10308
rect 5845 9276 6153 9296
rect 5845 9274 5851 9276
rect 5907 9274 5931 9276
rect 5987 9274 6011 9276
rect 6067 9274 6091 9276
rect 6147 9274 6153 9276
rect 5907 9222 5909 9274
rect 6089 9222 6091 9274
rect 5845 9220 5851 9222
rect 5907 9220 5931 9222
rect 5987 9220 6011 9222
rect 6067 9220 6091 9222
rect 6147 9220 6153 9222
rect 5845 9200 6153 9220
rect 5845 8188 6153 8208
rect 5845 8186 5851 8188
rect 5907 8186 5931 8188
rect 5987 8186 6011 8188
rect 6067 8186 6091 8188
rect 6147 8186 6153 8188
rect 5907 8134 5909 8186
rect 6089 8134 6091 8186
rect 5845 8132 5851 8134
rect 5907 8132 5931 8134
rect 5987 8132 6011 8134
rect 6067 8132 6091 8134
rect 6147 8132 6153 8134
rect 5845 8112 6153 8132
rect 5845 7100 6153 7120
rect 5845 7098 5851 7100
rect 5907 7098 5931 7100
rect 5987 7098 6011 7100
rect 6067 7098 6091 7100
rect 6147 7098 6153 7100
rect 5907 7046 5909 7098
rect 6089 7046 6091 7098
rect 5845 7044 5851 7046
rect 5907 7044 5931 7046
rect 5987 7044 6011 7046
rect 6067 7044 6091 7046
rect 6147 7044 6153 7046
rect 5845 7024 6153 7044
rect 6196 6322 6224 12378
rect 6288 12322 6316 12951
rect 6472 12442 6500 13892
rect 6656 13274 6684 15370
rect 6748 15366 6776 15982
rect 6918 15943 6974 15952
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6748 13410 6776 13874
rect 6840 13530 6868 15438
rect 6918 14920 6974 14929
rect 6918 14855 6974 14864
rect 6932 14550 6960 14855
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6932 13841 6960 14350
rect 6918 13832 6974 13841
rect 6918 13767 6974 13776
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6748 13382 6868 13410
rect 6564 13246 6684 13274
rect 6840 13274 6868 13382
rect 6736 13252 6788 13258
rect 6564 13190 6592 13246
rect 6840 13246 6960 13274
rect 6736 13194 6788 13200
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6288 12294 6408 12322
rect 6380 12238 6408 12294
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 11626 6592 12174
rect 6656 11762 6684 12582
rect 6748 12434 6776 13194
rect 6932 12753 6960 13246
rect 7024 12986 7052 16594
rect 7116 16538 7144 17292
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7208 16794 7236 17138
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7300 16697 7328 18226
rect 7852 18193 7880 18702
rect 7838 18184 7894 18193
rect 7838 18119 7894 18128
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7286 16688 7342 16697
rect 7392 16658 7420 17614
rect 7477 17436 7785 17456
rect 7477 17434 7483 17436
rect 7539 17434 7563 17436
rect 7619 17434 7643 17436
rect 7699 17434 7723 17436
rect 7779 17434 7785 17436
rect 7539 17382 7541 17434
rect 7721 17382 7723 17434
rect 7477 17380 7483 17382
rect 7539 17380 7563 17382
rect 7619 17380 7643 17382
rect 7699 17380 7723 17382
rect 7779 17380 7785 17382
rect 7477 17360 7785 17380
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7668 16794 7696 17206
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7286 16623 7342 16632
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7116 16510 7420 16538
rect 7760 16522 7788 17206
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7208 16114 7236 16390
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7116 15473 7144 16050
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15570 7328 15846
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7102 15464 7158 15473
rect 7102 15399 7158 15408
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 14074 7144 14758
rect 7208 14385 7236 15506
rect 7392 14822 7420 16510
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7477 16348 7785 16368
rect 7477 16346 7483 16348
rect 7539 16346 7563 16348
rect 7619 16346 7643 16348
rect 7699 16346 7723 16348
rect 7779 16346 7785 16348
rect 7539 16294 7541 16346
rect 7721 16294 7723 16346
rect 7477 16292 7483 16294
rect 7539 16292 7563 16294
rect 7619 16292 7643 16294
rect 7699 16292 7723 16294
rect 7779 16292 7785 16294
rect 7477 16272 7785 16292
rect 7852 16182 7880 18022
rect 7944 17241 7972 19382
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 7930 17232 7986 17241
rect 7930 17167 7986 17176
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 7944 15910 7972 16594
rect 8036 16454 8064 17478
rect 8128 16658 8156 17478
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7477 15260 7785 15280
rect 7477 15258 7483 15260
rect 7539 15258 7563 15260
rect 7619 15258 7643 15260
rect 7699 15258 7723 15260
rect 7779 15258 7785 15260
rect 7539 15206 7541 15258
rect 7721 15206 7723 15258
rect 7477 15204 7483 15206
rect 7539 15204 7563 15206
rect 7619 15204 7643 15206
rect 7699 15204 7723 15206
rect 7779 15204 7785 15206
rect 7477 15184 7785 15204
rect 7930 15192 7986 15201
rect 7930 15127 7932 15136
rect 7984 15127 7986 15136
rect 7932 15098 7984 15104
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7484 14906 7512 14962
rect 7484 14878 7788 14906
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7286 14648 7342 14657
rect 7286 14583 7342 14592
rect 7300 14482 7328 14583
rect 7668 14521 7696 14758
rect 7760 14550 7788 14878
rect 7840 14884 7892 14890
rect 7840 14826 7892 14832
rect 7748 14544 7800 14550
rect 7654 14512 7710 14521
rect 7288 14476 7340 14482
rect 7748 14486 7800 14492
rect 7654 14447 7710 14456
rect 7288 14418 7340 14424
rect 7668 14414 7696 14447
rect 7656 14408 7708 14414
rect 7194 14376 7250 14385
rect 7656 14350 7708 14356
rect 7194 14311 7250 14320
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7116 13977 7144 14010
rect 7102 13968 7158 13977
rect 7102 13903 7158 13912
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7208 12889 7236 13806
rect 7300 13734 7328 14214
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7392 12986 7420 14282
rect 7477 14172 7785 14192
rect 7477 14170 7483 14172
rect 7539 14170 7563 14172
rect 7619 14170 7643 14172
rect 7699 14170 7723 14172
rect 7779 14170 7785 14172
rect 7539 14118 7541 14170
rect 7721 14118 7723 14170
rect 7477 14116 7483 14118
rect 7539 14116 7563 14118
rect 7619 14116 7643 14118
rect 7699 14116 7723 14118
rect 7779 14116 7785 14118
rect 7477 14096 7785 14116
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 13394 7604 13806
rect 7668 13802 7696 13942
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7654 13560 7710 13569
rect 7654 13495 7656 13504
rect 7708 13495 7710 13504
rect 7656 13466 7708 13472
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7477 13084 7785 13104
rect 7477 13082 7483 13084
rect 7539 13082 7563 13084
rect 7619 13082 7643 13084
rect 7699 13082 7723 13084
rect 7779 13082 7785 13084
rect 7539 13030 7541 13082
rect 7721 13030 7723 13082
rect 7477 13028 7483 13030
rect 7539 13028 7563 13030
rect 7619 13028 7643 13030
rect 7699 13028 7723 13030
rect 7779 13028 7785 13030
rect 7477 13008 7785 13028
rect 7852 12986 7880 14826
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7194 12880 7250 12889
rect 7104 12844 7156 12850
rect 7194 12815 7250 12824
rect 7380 12844 7432 12850
rect 7104 12786 7156 12792
rect 7380 12786 7432 12792
rect 6918 12744 6974 12753
rect 6918 12679 6974 12688
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6748 12406 6868 12434
rect 6840 11914 6868 12406
rect 7024 12306 7052 12650
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6748 11886 6868 11914
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6564 11286 6592 11562
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 5845 6012 6153 6032
rect 5845 6010 5851 6012
rect 5907 6010 5931 6012
rect 5987 6010 6011 6012
rect 6067 6010 6091 6012
rect 6147 6010 6153 6012
rect 5907 5958 5909 6010
rect 6089 5958 6091 6010
rect 5845 5956 5851 5958
rect 5907 5956 5931 5958
rect 5987 5956 6011 5958
rect 6067 5956 6091 5958
rect 6147 5956 6153 5958
rect 5845 5936 6153 5956
rect 6748 5710 6776 11886
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11354 6868 11698
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7116 10538 7144 12786
rect 7286 11248 7342 11257
rect 7286 11183 7342 11192
rect 7300 11150 7328 11183
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7392 11082 7420 12786
rect 7477 11996 7785 12016
rect 7477 11994 7483 11996
rect 7539 11994 7563 11996
rect 7619 11994 7643 11996
rect 7699 11994 7723 11996
rect 7779 11994 7785 11996
rect 7539 11942 7541 11994
rect 7721 11942 7723 11994
rect 7477 11940 7483 11942
rect 7539 11940 7563 11942
rect 7619 11940 7643 11942
rect 7699 11940 7723 11942
rect 7779 11940 7785 11942
rect 7477 11920 7785 11940
rect 7944 11354 7972 14350
rect 8036 14074 8064 16390
rect 8128 15502 8156 16458
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8128 13433 8156 14486
rect 8114 13424 8170 13433
rect 8114 13359 8170 13368
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12442 8064 13262
rect 8220 12918 8248 40287
rect 8312 37346 8340 43386
rect 8404 37466 8432 44134
rect 8496 41414 8524 59366
rect 8588 55865 8616 68614
rect 8680 62490 8708 73714
rect 9496 73568 9548 73574
rect 9494 73536 9496 73545
rect 9548 73536 9550 73545
rect 9109 73468 9417 73488
rect 9494 73471 9550 73480
rect 9109 73466 9115 73468
rect 9171 73466 9195 73468
rect 9251 73466 9275 73468
rect 9331 73466 9355 73468
rect 9411 73466 9417 73468
rect 9171 73414 9173 73466
rect 9353 73414 9355 73466
rect 9109 73412 9115 73414
rect 9171 73412 9195 73414
rect 9251 73412 9275 73414
rect 9331 73412 9355 73414
rect 9411 73412 9417 73414
rect 9109 73392 9417 73412
rect 9876 73166 9904 75890
rect 10060 75449 10088 76230
rect 10046 75440 10102 75449
rect 10046 75375 10102 75384
rect 10140 75200 10192 75206
rect 10140 75142 10192 75148
rect 10048 74656 10100 74662
rect 10048 74598 10100 74604
rect 9956 74180 10008 74186
rect 9956 74122 10008 74128
rect 9864 73160 9916 73166
rect 9864 73102 9916 73108
rect 9968 73098 9996 74122
rect 10060 73953 10088 74598
rect 10152 74497 10180 75142
rect 10968 74928 11020 74934
rect 10966 74896 10968 74905
rect 11020 74896 11022 74905
rect 10966 74831 11022 74840
rect 10138 74488 10194 74497
rect 10138 74423 10194 74432
rect 10232 74316 10284 74322
rect 10232 74258 10284 74264
rect 10140 74112 10192 74118
rect 10140 74054 10192 74060
rect 10046 73944 10102 73953
rect 10046 73879 10102 73888
rect 10048 73568 10100 73574
rect 10048 73510 10100 73516
rect 9956 73092 10008 73098
rect 9956 73034 10008 73040
rect 10060 73001 10088 73510
rect 10152 73234 10180 74054
rect 10140 73228 10192 73234
rect 10140 73170 10192 73176
rect 10244 73166 10272 74258
rect 10232 73160 10284 73166
rect 10232 73102 10284 73108
rect 10046 72992 10102 73001
rect 10046 72927 10102 72936
rect 9036 72684 9088 72690
rect 9036 72626 9088 72632
rect 9048 70106 9076 72626
rect 9310 72584 9366 72593
rect 9310 72519 9312 72528
rect 9364 72519 9366 72528
rect 9312 72490 9364 72496
rect 10140 72480 10192 72486
rect 10140 72422 10192 72428
rect 9109 72380 9417 72400
rect 9109 72378 9115 72380
rect 9171 72378 9195 72380
rect 9251 72378 9275 72380
rect 9331 72378 9355 72380
rect 9411 72378 9417 72380
rect 9171 72326 9173 72378
rect 9353 72326 9355 72378
rect 9109 72324 9115 72326
rect 9171 72324 9195 72326
rect 9251 72324 9275 72326
rect 9331 72324 9355 72326
rect 9411 72324 9417 72326
rect 9109 72304 9417 72324
rect 9310 72040 9366 72049
rect 9310 71975 9366 71984
rect 9324 71942 9352 71975
rect 9312 71936 9364 71942
rect 9312 71878 9364 71884
rect 10048 71936 10100 71942
rect 10048 71878 10100 71884
rect 9772 71392 9824 71398
rect 9772 71334 9824 71340
rect 9109 71292 9417 71312
rect 9109 71290 9115 71292
rect 9171 71290 9195 71292
rect 9251 71290 9275 71292
rect 9331 71290 9355 71292
rect 9411 71290 9417 71292
rect 9171 71238 9173 71290
rect 9353 71238 9355 71290
rect 9109 71236 9115 71238
rect 9171 71236 9195 71238
rect 9251 71236 9275 71238
rect 9331 71236 9355 71238
rect 9411 71236 9417 71238
rect 9109 71216 9417 71236
rect 9109 70204 9417 70224
rect 9109 70202 9115 70204
rect 9171 70202 9195 70204
rect 9251 70202 9275 70204
rect 9331 70202 9355 70204
rect 9411 70202 9417 70204
rect 9171 70150 9173 70202
rect 9353 70150 9355 70202
rect 9109 70148 9115 70150
rect 9171 70148 9195 70150
rect 9251 70148 9275 70150
rect 9331 70148 9355 70150
rect 9411 70148 9417 70150
rect 9109 70128 9417 70148
rect 9036 70100 9088 70106
rect 9036 70042 9088 70048
rect 8852 69760 8904 69766
rect 8852 69702 8904 69708
rect 8864 69358 8892 69702
rect 9588 69556 9640 69562
rect 9588 69498 9640 69504
rect 9036 69420 9088 69426
rect 9036 69362 9088 69368
rect 8852 69352 8904 69358
rect 9048 69329 9076 69362
rect 8852 69294 8904 69300
rect 9034 69320 9090 69329
rect 8864 68134 8892 69294
rect 9034 69255 9090 69264
rect 9496 69284 9548 69290
rect 9496 69226 9548 69232
rect 9508 69193 9536 69226
rect 9494 69184 9550 69193
rect 9109 69116 9417 69136
rect 9494 69119 9550 69128
rect 9109 69114 9115 69116
rect 9171 69114 9195 69116
rect 9251 69114 9275 69116
rect 9331 69114 9355 69116
rect 9411 69114 9417 69116
rect 9171 69062 9173 69114
rect 9353 69062 9355 69114
rect 9109 69060 9115 69062
rect 9171 69060 9195 69062
rect 9251 69060 9275 69062
rect 9331 69060 9355 69062
rect 9411 69060 9417 69062
rect 9109 69040 9417 69060
rect 9496 68672 9548 68678
rect 9496 68614 9548 68620
rect 9508 68406 9536 68614
rect 9496 68400 9548 68406
rect 9600 68377 9628 69498
rect 9784 69426 9812 71334
rect 10060 71097 10088 71878
rect 10152 71641 10180 72422
rect 10138 71632 10194 71641
rect 10138 71567 10194 71576
rect 10140 71392 10192 71398
rect 10140 71334 10192 71340
rect 10046 71088 10102 71097
rect 10046 71023 10102 71032
rect 10048 70848 10100 70854
rect 10048 70790 10100 70796
rect 9864 70440 9916 70446
rect 9864 70382 9916 70388
rect 9876 69766 9904 70382
rect 10060 70145 10088 70790
rect 10152 70689 10180 71334
rect 10138 70680 10194 70689
rect 10138 70615 10194 70624
rect 10046 70136 10102 70145
rect 10046 70071 10102 70080
rect 10244 69970 10272 73102
rect 10232 69964 10284 69970
rect 10232 69906 10284 69912
rect 9956 69828 10008 69834
rect 9956 69770 10008 69776
rect 9864 69760 9916 69766
rect 9864 69702 9916 69708
rect 9772 69420 9824 69426
rect 9772 69362 9824 69368
rect 9496 68342 9548 68348
rect 9586 68368 9642 68377
rect 9586 68303 9642 68312
rect 8760 68128 8812 68134
rect 8760 68070 8812 68076
rect 8852 68128 8904 68134
rect 8852 68070 8904 68076
rect 8772 67833 8800 68070
rect 8758 67824 8814 67833
rect 8758 67759 8814 67768
rect 8864 67658 8892 68070
rect 9109 68028 9417 68048
rect 9109 68026 9115 68028
rect 9171 68026 9195 68028
rect 9251 68026 9275 68028
rect 9331 68026 9355 68028
rect 9411 68026 9417 68028
rect 9171 67974 9173 68026
rect 9353 67974 9355 68026
rect 9109 67972 9115 67974
rect 9171 67972 9195 67974
rect 9251 67972 9275 67974
rect 9331 67972 9355 67974
rect 9411 67972 9417 67974
rect 9109 67952 9417 67972
rect 9404 67856 9456 67862
rect 9404 67798 9456 67804
rect 9416 67697 9444 67798
rect 9402 67688 9458 67697
rect 8852 67652 8904 67658
rect 9784 67658 9812 69362
rect 9876 68678 9904 69702
rect 9864 68672 9916 68678
rect 9864 68614 9916 68620
rect 9968 68474 9996 69770
rect 10244 69442 10272 69906
rect 10414 69728 10470 69737
rect 10414 69663 10470 69672
rect 10428 69562 10456 69663
rect 10416 69556 10468 69562
rect 10416 69498 10468 69504
rect 10152 69414 10272 69442
rect 10152 69358 10180 69414
rect 10140 69352 10192 69358
rect 10140 69294 10192 69300
rect 9956 68468 10008 68474
rect 9956 68410 10008 68416
rect 10152 68406 10180 69294
rect 10140 68400 10192 68406
rect 10140 68342 10192 68348
rect 10152 67794 10180 68342
rect 10140 67788 10192 67794
rect 10140 67730 10192 67736
rect 9402 67623 9458 67632
rect 9772 67652 9824 67658
rect 8852 67594 8904 67600
rect 9772 67594 9824 67600
rect 8864 65226 8892 67594
rect 10152 67386 10180 67730
rect 10140 67380 10192 67386
rect 10140 67322 10192 67328
rect 8944 67244 8996 67250
rect 8944 67186 8996 67192
rect 8956 66570 8984 67186
rect 9128 67176 9180 67182
rect 9048 67136 9128 67164
rect 9048 66638 9076 67136
rect 9128 67118 9180 67124
rect 9680 67176 9732 67182
rect 9680 67118 9732 67124
rect 9496 67108 9548 67114
rect 9496 67050 9548 67056
rect 9109 66940 9417 66960
rect 9109 66938 9115 66940
rect 9171 66938 9195 66940
rect 9251 66938 9275 66940
rect 9331 66938 9355 66940
rect 9411 66938 9417 66940
rect 9171 66886 9173 66938
rect 9353 66886 9355 66938
rect 9109 66884 9115 66886
rect 9171 66884 9195 66886
rect 9251 66884 9275 66886
rect 9331 66884 9355 66886
rect 9411 66884 9417 66886
rect 9109 66864 9417 66884
rect 9508 66881 9536 67050
rect 9494 66872 9550 66881
rect 9494 66807 9550 66816
rect 9692 66638 9720 67118
rect 10048 67040 10100 67046
rect 10048 66982 10100 66988
rect 9036 66632 9088 66638
rect 9404 66632 9456 66638
rect 9036 66574 9088 66580
rect 9402 66600 9404 66609
rect 9680 66632 9732 66638
rect 9456 66600 9458 66609
rect 8944 66564 8996 66570
rect 9402 66535 9458 66544
rect 9600 66592 9680 66620
rect 8944 66506 8996 66512
rect 8956 65414 8984 66506
rect 9496 65952 9548 65958
rect 9494 65920 9496 65929
rect 9548 65920 9550 65929
rect 9109 65852 9417 65872
rect 9494 65855 9550 65864
rect 9109 65850 9115 65852
rect 9171 65850 9195 65852
rect 9251 65850 9275 65852
rect 9331 65850 9355 65852
rect 9411 65850 9417 65852
rect 9171 65798 9173 65850
rect 9353 65798 9355 65850
rect 9109 65796 9115 65798
rect 9171 65796 9195 65798
rect 9251 65796 9275 65798
rect 9331 65796 9355 65798
rect 9411 65796 9417 65798
rect 9109 65776 9417 65796
rect 9036 65680 9088 65686
rect 9036 65622 9088 65628
rect 8944 65408 8996 65414
rect 8944 65350 8996 65356
rect 8864 65198 8984 65226
rect 8760 65068 8812 65074
rect 8760 65010 8812 65016
rect 8772 64569 8800 65010
rect 8758 64560 8814 64569
rect 8758 64495 8814 64504
rect 8852 64320 8904 64326
rect 8852 64262 8904 64268
rect 8668 62484 8720 62490
rect 8668 62426 8720 62432
rect 8668 60784 8720 60790
rect 8668 60726 8720 60732
rect 8680 60217 8708 60726
rect 8760 60512 8812 60518
rect 8760 60454 8812 60460
rect 8666 60208 8722 60217
rect 8666 60143 8722 60152
rect 8668 57928 8720 57934
rect 8668 57870 8720 57876
rect 8574 55856 8630 55865
rect 8574 55791 8630 55800
rect 8680 55706 8708 57870
rect 8588 55678 8708 55706
rect 8588 53553 8616 55678
rect 8668 53984 8720 53990
rect 8668 53926 8720 53932
rect 8574 53544 8630 53553
rect 8574 53479 8630 53488
rect 8576 53440 8628 53446
rect 8576 53382 8628 53388
rect 8588 46442 8616 53382
rect 8680 49994 8708 53926
rect 8772 50182 8800 60454
rect 8864 58682 8892 64262
rect 8852 58676 8904 58682
rect 8852 58618 8904 58624
rect 8852 58540 8904 58546
rect 8852 58482 8904 58488
rect 8864 51610 8892 58482
rect 8852 51604 8904 51610
rect 8852 51546 8904 51552
rect 8956 51105 8984 65198
rect 9048 64122 9076 65622
rect 9600 65618 9628 66592
rect 9680 66574 9732 66580
rect 10060 66473 10088 66982
rect 10140 66564 10192 66570
rect 10140 66506 10192 66512
rect 10046 66464 10102 66473
rect 10046 66399 10102 66408
rect 10048 65952 10100 65958
rect 10048 65894 10100 65900
rect 9588 65612 9640 65618
rect 9588 65554 9640 65560
rect 9496 65544 9548 65550
rect 9496 65486 9548 65492
rect 9508 65210 9536 65486
rect 9600 65226 9628 65554
rect 10060 65521 10088 65894
rect 10046 65512 10102 65521
rect 9864 65476 9916 65482
rect 10046 65447 10102 65456
rect 9864 65418 9916 65424
rect 9496 65204 9548 65210
rect 9600 65198 9720 65226
rect 9496 65146 9548 65152
rect 9588 65068 9640 65074
rect 9588 65010 9640 65016
rect 9496 64864 9548 64870
rect 9496 64806 9548 64812
rect 9109 64764 9417 64784
rect 9109 64762 9115 64764
rect 9171 64762 9195 64764
rect 9251 64762 9275 64764
rect 9331 64762 9355 64764
rect 9411 64762 9417 64764
rect 9171 64710 9173 64762
rect 9353 64710 9355 64762
rect 9109 64708 9115 64710
rect 9171 64708 9195 64710
rect 9251 64708 9275 64710
rect 9331 64708 9355 64710
rect 9411 64708 9417 64710
rect 9109 64688 9417 64708
rect 9508 64462 9536 64806
rect 9496 64456 9548 64462
rect 9496 64398 9548 64404
rect 9496 64320 9548 64326
rect 9496 64262 9548 64268
rect 9036 64116 9088 64122
rect 9036 64058 9088 64064
rect 9048 63034 9076 64058
rect 9508 63900 9536 64262
rect 9600 64025 9628 65010
rect 9692 64938 9720 65198
rect 9876 65074 9904 65418
rect 9864 65068 9916 65074
rect 9864 65010 9916 65016
rect 10046 64968 10102 64977
rect 9680 64932 9732 64938
rect 10046 64903 10048 64912
rect 9680 64874 9732 64880
rect 10100 64903 10102 64912
rect 10048 64874 10100 64880
rect 9692 64462 9720 64874
rect 9680 64456 9732 64462
rect 9680 64398 9732 64404
rect 10152 64138 10180 66506
rect 11704 66156 11756 66162
rect 11704 66098 11756 66104
rect 10600 65476 10652 65482
rect 10600 65418 10652 65424
rect 10416 64388 10468 64394
rect 10416 64330 10468 64336
rect 10060 64110 10180 64138
rect 9586 64016 9642 64025
rect 9586 63951 9642 63960
rect 9588 63912 9640 63918
rect 9508 63872 9588 63900
rect 9588 63854 9640 63860
rect 9109 63676 9417 63696
rect 9109 63674 9115 63676
rect 9171 63674 9195 63676
rect 9251 63674 9275 63676
rect 9331 63674 9355 63676
rect 9411 63674 9417 63676
rect 9171 63622 9173 63674
rect 9353 63622 9355 63674
rect 9109 63620 9115 63622
rect 9171 63620 9195 63622
rect 9251 63620 9275 63622
rect 9331 63620 9355 63622
rect 9411 63620 9417 63622
rect 9109 63600 9417 63620
rect 9494 63608 9550 63617
rect 9494 63543 9550 63552
rect 9508 63374 9536 63543
rect 9496 63368 9548 63374
rect 9496 63310 9548 63316
rect 9496 63232 9548 63238
rect 9496 63174 9548 63180
rect 9036 63028 9088 63034
rect 9036 62970 9088 62976
rect 9109 62588 9417 62608
rect 9109 62586 9115 62588
rect 9171 62586 9195 62588
rect 9251 62586 9275 62588
rect 9331 62586 9355 62588
rect 9411 62586 9417 62588
rect 9171 62534 9173 62586
rect 9353 62534 9355 62586
rect 9109 62532 9115 62534
rect 9171 62532 9195 62534
rect 9251 62532 9275 62534
rect 9331 62532 9355 62534
rect 9411 62532 9417 62534
rect 9109 62512 9417 62532
rect 9312 62280 9364 62286
rect 9312 62222 9364 62228
rect 9324 61713 9352 62222
rect 9310 61704 9366 61713
rect 9310 61639 9366 61648
rect 9109 61500 9417 61520
rect 9109 61498 9115 61500
rect 9171 61498 9195 61500
rect 9251 61498 9275 61500
rect 9331 61498 9355 61500
rect 9411 61498 9417 61500
rect 9171 61446 9173 61498
rect 9353 61446 9355 61498
rect 9109 61444 9115 61446
rect 9171 61444 9195 61446
rect 9251 61444 9275 61446
rect 9331 61444 9355 61446
rect 9411 61444 9417 61446
rect 9109 61424 9417 61444
rect 9508 61198 9536 63174
rect 9600 62898 9628 63854
rect 9588 62892 9640 62898
rect 9588 62834 9640 62840
rect 9600 61690 9628 62834
rect 9600 61662 9720 61690
rect 9588 61600 9640 61606
rect 9588 61542 9640 61548
rect 9404 61192 9456 61198
rect 9404 61134 9456 61140
rect 9496 61192 9548 61198
rect 9600 61169 9628 61542
rect 9692 61198 9720 61662
rect 9680 61192 9732 61198
rect 9496 61134 9548 61140
rect 9586 61160 9642 61169
rect 9310 60752 9366 60761
rect 9416 60734 9444 61134
rect 9680 61134 9732 61140
rect 9586 61095 9642 61104
rect 10060 60734 10088 64110
rect 10140 63980 10192 63986
rect 10140 63922 10192 63928
rect 10152 63073 10180 63922
rect 10232 63368 10284 63374
rect 10232 63310 10284 63316
rect 10138 63064 10194 63073
rect 10138 62999 10194 63008
rect 10140 62892 10192 62898
rect 10140 62834 10192 62840
rect 10152 62121 10180 62834
rect 10244 62665 10272 63310
rect 10230 62656 10286 62665
rect 10230 62591 10286 62600
rect 10138 62112 10194 62121
rect 10138 62047 10194 62056
rect 9416 60706 9536 60734
rect 10060 60706 10180 60734
rect 9310 60687 9312 60696
rect 9364 60687 9366 60696
rect 9312 60658 9364 60664
rect 9109 60412 9417 60432
rect 9109 60410 9115 60412
rect 9171 60410 9195 60412
rect 9251 60410 9275 60412
rect 9331 60410 9355 60412
rect 9411 60410 9417 60412
rect 9171 60358 9173 60410
rect 9353 60358 9355 60410
rect 9109 60356 9115 60358
rect 9171 60356 9195 60358
rect 9251 60356 9275 60358
rect 9331 60356 9355 60358
rect 9411 60356 9417 60358
rect 9109 60336 9417 60356
rect 9218 59800 9274 59809
rect 9218 59735 9274 59744
rect 9232 59702 9260 59735
rect 9220 59696 9272 59702
rect 9220 59638 9272 59644
rect 9109 59324 9417 59344
rect 9109 59322 9115 59324
rect 9171 59322 9195 59324
rect 9251 59322 9275 59324
rect 9331 59322 9355 59324
rect 9411 59322 9417 59324
rect 9171 59270 9173 59322
rect 9353 59270 9355 59322
rect 9109 59268 9115 59270
rect 9171 59268 9195 59270
rect 9251 59268 9275 59270
rect 9331 59268 9355 59270
rect 9411 59268 9417 59270
rect 9109 59248 9417 59268
rect 9109 58236 9417 58256
rect 9109 58234 9115 58236
rect 9171 58234 9195 58236
rect 9251 58234 9275 58236
rect 9331 58234 9355 58236
rect 9411 58234 9417 58236
rect 9171 58182 9173 58234
rect 9353 58182 9355 58234
rect 9109 58180 9115 58182
rect 9171 58180 9195 58182
rect 9251 58180 9275 58182
rect 9331 58180 9355 58182
rect 9411 58180 9417 58182
rect 9109 58160 9417 58180
rect 9036 57452 9088 57458
rect 9036 57394 9088 57400
rect 9220 57452 9272 57458
rect 9220 57394 9272 57400
rect 8942 51096 8998 51105
rect 8942 51031 8998 51040
rect 8944 50924 8996 50930
rect 8944 50866 8996 50872
rect 8852 50856 8904 50862
rect 8852 50798 8904 50804
rect 8760 50176 8812 50182
rect 8760 50118 8812 50124
rect 8680 49966 8800 49994
rect 8666 49872 8722 49881
rect 8666 49807 8668 49816
rect 8720 49807 8722 49816
rect 8668 49778 8720 49784
rect 8668 49700 8720 49706
rect 8668 49642 8720 49648
rect 8680 47546 8708 49642
rect 8772 48210 8800 49966
rect 8864 48686 8892 50798
rect 8956 49434 8984 50866
rect 9048 50522 9076 57394
rect 9232 57361 9260 57394
rect 9218 57352 9274 57361
rect 9218 57287 9274 57296
rect 9109 57148 9417 57168
rect 9109 57146 9115 57148
rect 9171 57146 9195 57148
rect 9251 57146 9275 57148
rect 9331 57146 9355 57148
rect 9411 57146 9417 57148
rect 9171 57094 9173 57146
rect 9353 57094 9355 57146
rect 9109 57092 9115 57094
rect 9171 57092 9195 57094
rect 9251 57092 9275 57094
rect 9331 57092 9355 57094
rect 9411 57092 9417 57094
rect 9109 57072 9417 57092
rect 9508 56352 9536 60706
rect 10048 60104 10100 60110
rect 10048 60046 10100 60052
rect 9956 59628 10008 59634
rect 9956 59570 10008 59576
rect 9968 58857 9996 59570
rect 10060 59265 10088 60046
rect 10046 59256 10102 59265
rect 10046 59191 10102 59200
rect 9954 58848 10010 58857
rect 9954 58783 10010 58792
rect 9956 58540 10008 58546
rect 9956 58482 10008 58488
rect 9968 57905 9996 58482
rect 9954 57896 10010 57905
rect 9954 57831 10010 57840
rect 9588 57452 9640 57458
rect 9588 57394 9640 57400
rect 9600 56545 9628 57394
rect 10048 56772 10100 56778
rect 10048 56714 10100 56720
rect 9586 56536 9642 56545
rect 9586 56471 9642 56480
rect 9864 56364 9916 56370
rect 9508 56324 9628 56352
rect 9109 56060 9417 56080
rect 9109 56058 9115 56060
rect 9171 56058 9195 56060
rect 9251 56058 9275 56060
rect 9331 56058 9355 56060
rect 9411 56058 9417 56060
rect 9171 56006 9173 56058
rect 9353 56006 9355 56058
rect 9109 56004 9115 56006
rect 9171 56004 9195 56006
rect 9251 56004 9275 56006
rect 9331 56004 9355 56006
rect 9411 56004 9417 56006
rect 9109 55984 9417 56004
rect 9109 54972 9417 54992
rect 9109 54970 9115 54972
rect 9171 54970 9195 54972
rect 9251 54970 9275 54972
rect 9331 54970 9355 54972
rect 9411 54970 9417 54972
rect 9171 54918 9173 54970
rect 9353 54918 9355 54970
rect 9109 54916 9115 54918
rect 9171 54916 9195 54918
rect 9251 54916 9275 54918
rect 9331 54916 9355 54918
rect 9411 54916 9417 54918
rect 9109 54896 9417 54916
rect 9600 54210 9628 56324
rect 9864 56306 9916 56312
rect 9876 56001 9904 56306
rect 9862 55992 9918 56001
rect 9862 55927 9918 55936
rect 9864 55752 9916 55758
rect 9864 55694 9916 55700
rect 9876 55593 9904 55694
rect 9862 55584 9918 55593
rect 9862 55519 9918 55528
rect 9864 55276 9916 55282
rect 9864 55218 9916 55224
rect 9876 55049 9904 55218
rect 9862 55040 9918 55049
rect 9862 54975 9918 54984
rect 9954 54632 10010 54641
rect 9954 54567 9956 54576
rect 10008 54567 10010 54576
rect 9956 54538 10008 54544
rect 9496 54188 9548 54194
rect 9600 54182 9720 54210
rect 9496 54130 9548 54136
rect 9109 53884 9417 53904
rect 9109 53882 9115 53884
rect 9171 53882 9195 53884
rect 9251 53882 9275 53884
rect 9331 53882 9355 53884
rect 9411 53882 9417 53884
rect 9171 53830 9173 53882
rect 9353 53830 9355 53882
rect 9109 53828 9115 53830
rect 9171 53828 9195 53830
rect 9251 53828 9275 53830
rect 9331 53828 9355 53830
rect 9411 53828 9417 53830
rect 9109 53808 9417 53828
rect 9508 53689 9536 54130
rect 9586 54088 9642 54097
rect 9586 54023 9642 54032
rect 9494 53680 9550 53689
rect 9494 53615 9550 53624
rect 9600 53582 9628 54023
rect 9588 53576 9640 53582
rect 9588 53518 9640 53524
rect 9692 53394 9720 54182
rect 9956 54188 10008 54194
rect 9956 54130 10008 54136
rect 9864 53576 9916 53582
rect 9864 53518 9916 53524
rect 9600 53366 9720 53394
rect 9109 52796 9417 52816
rect 9109 52794 9115 52796
rect 9171 52794 9195 52796
rect 9251 52794 9275 52796
rect 9331 52794 9355 52796
rect 9411 52794 9417 52796
rect 9171 52742 9173 52794
rect 9353 52742 9355 52794
rect 9109 52740 9115 52742
rect 9171 52740 9195 52742
rect 9251 52740 9275 52742
rect 9331 52740 9355 52742
rect 9411 52740 9417 52742
rect 9109 52720 9417 52740
rect 9128 52488 9180 52494
rect 9128 52430 9180 52436
rect 9140 52193 9168 52430
rect 9126 52184 9182 52193
rect 9126 52119 9182 52128
rect 9496 52012 9548 52018
rect 9496 51954 9548 51960
rect 9508 51785 9536 51954
rect 9494 51776 9550 51785
rect 9109 51708 9417 51728
rect 9494 51711 9550 51720
rect 9109 51706 9115 51708
rect 9171 51706 9195 51708
rect 9251 51706 9275 51708
rect 9331 51706 9355 51708
rect 9411 51706 9417 51708
rect 9171 51654 9173 51706
rect 9353 51654 9355 51706
rect 9109 51652 9115 51654
rect 9171 51652 9195 51654
rect 9251 51652 9275 51654
rect 9331 51652 9355 51654
rect 9411 51652 9417 51654
rect 9109 51632 9417 51652
rect 9600 51542 9628 53366
rect 9772 53100 9824 53106
rect 9772 53042 9824 53048
rect 9588 51536 9640 51542
rect 9588 51478 9640 51484
rect 9496 51332 9548 51338
rect 9496 51274 9548 51280
rect 9508 50810 9536 51274
rect 9680 51264 9732 51270
rect 9680 51206 9732 51212
rect 9692 50810 9720 51206
rect 9784 50998 9812 53042
rect 9876 52737 9904 53518
rect 9968 53145 9996 54130
rect 10060 53530 10088 56714
rect 10152 53650 10180 60706
rect 10232 60648 10284 60654
rect 10230 60616 10232 60625
rect 10284 60616 10286 60625
rect 10230 60551 10286 60560
rect 10232 58948 10284 58954
rect 10232 58890 10284 58896
rect 10244 58313 10272 58890
rect 10230 58304 10286 58313
rect 10230 58239 10286 58248
rect 10324 57860 10376 57866
rect 10324 57802 10376 57808
rect 10336 56953 10364 57802
rect 10322 56944 10378 56953
rect 10232 56908 10284 56914
rect 10322 56879 10378 56888
rect 10232 56850 10284 56856
rect 10244 53990 10272 56850
rect 10428 55842 10456 64330
rect 10508 61124 10560 61130
rect 10508 61066 10560 61072
rect 10336 55814 10456 55842
rect 10232 53984 10284 53990
rect 10232 53926 10284 53932
rect 10140 53644 10192 53650
rect 10140 53586 10192 53592
rect 10060 53502 10272 53530
rect 10048 53440 10100 53446
rect 10048 53382 10100 53388
rect 10140 53440 10192 53446
rect 10140 53382 10192 53388
rect 9954 53136 10010 53145
rect 9954 53071 10010 53080
rect 10060 52850 10088 53382
rect 9968 52822 10088 52850
rect 9862 52728 9918 52737
rect 9862 52663 9918 52672
rect 9864 52012 9916 52018
rect 9864 51954 9916 51960
rect 9772 50992 9824 50998
rect 9772 50934 9824 50940
rect 9876 50833 9904 51954
rect 9862 50824 9918 50833
rect 9508 50782 9628 50810
rect 9692 50782 9812 50810
rect 9600 50726 9628 50782
rect 9496 50720 9548 50726
rect 9496 50662 9548 50668
rect 9588 50720 9640 50726
rect 9588 50662 9640 50668
rect 9109 50620 9417 50640
rect 9109 50618 9115 50620
rect 9171 50618 9195 50620
rect 9251 50618 9275 50620
rect 9331 50618 9355 50620
rect 9411 50618 9417 50620
rect 9171 50566 9173 50618
rect 9353 50566 9355 50618
rect 9109 50564 9115 50566
rect 9171 50564 9195 50566
rect 9251 50564 9275 50566
rect 9331 50564 9355 50566
rect 9411 50564 9417 50566
rect 9109 50544 9417 50564
rect 9036 50516 9088 50522
rect 9036 50458 9088 50464
rect 9126 50416 9182 50425
rect 9508 50386 9536 50662
rect 9126 50351 9182 50360
rect 9496 50380 9548 50386
rect 9036 50176 9088 50182
rect 9036 50118 9088 50124
rect 8944 49428 8996 49434
rect 8944 49370 8996 49376
rect 8956 48754 8984 49370
rect 8944 48748 8996 48754
rect 8944 48690 8996 48696
rect 8852 48680 8904 48686
rect 9048 48634 9076 50118
rect 9140 49706 9168 50351
rect 9496 50322 9548 50328
rect 9496 50176 9548 50182
rect 9496 50118 9548 50124
rect 9128 49700 9180 49706
rect 9128 49642 9180 49648
rect 9109 49532 9417 49552
rect 9109 49530 9115 49532
rect 9171 49530 9195 49532
rect 9251 49530 9275 49532
rect 9331 49530 9355 49532
rect 9411 49530 9417 49532
rect 9171 49478 9173 49530
rect 9353 49478 9355 49530
rect 9109 49476 9115 49478
rect 9171 49476 9195 49478
rect 9251 49476 9275 49478
rect 9331 49476 9355 49478
rect 9411 49476 9417 49478
rect 9109 49456 9417 49476
rect 9404 49224 9456 49230
rect 9404 49166 9456 49172
rect 9416 48754 9444 49166
rect 9508 48890 9536 50118
rect 9600 49298 9628 50662
rect 9680 50176 9732 50182
rect 9680 50118 9732 50124
rect 9588 49292 9640 49298
rect 9588 49234 9640 49240
rect 9692 49178 9720 50118
rect 9784 49366 9812 50782
rect 9862 50759 9918 50768
rect 9968 50454 9996 52822
rect 10048 51808 10100 51814
rect 10048 51750 10100 51756
rect 9956 50448 10008 50454
rect 9956 50390 10008 50396
rect 9864 50380 9916 50386
rect 9864 50322 9916 50328
rect 9876 49842 9904 50322
rect 9954 50144 10010 50153
rect 9954 50079 10010 50088
rect 9968 49978 9996 50079
rect 9956 49972 10008 49978
rect 9956 49914 10008 49920
rect 9864 49836 9916 49842
rect 9864 49778 9916 49784
rect 9876 49722 9904 49778
rect 9876 49694 9996 49722
rect 9772 49360 9824 49366
rect 9772 49302 9824 49308
rect 9600 49150 9720 49178
rect 9496 48884 9548 48890
rect 9496 48826 9548 48832
rect 9404 48748 9456 48754
rect 9404 48690 9456 48696
rect 8852 48622 8904 48628
rect 8956 48606 9076 48634
rect 8850 48512 8906 48521
rect 8850 48447 8906 48456
rect 8864 48346 8892 48447
rect 8852 48340 8904 48346
rect 8852 48282 8904 48288
rect 8760 48204 8812 48210
rect 8760 48146 8812 48152
rect 8852 48136 8904 48142
rect 8852 48078 8904 48084
rect 8680 47518 8800 47546
rect 8668 47456 8720 47462
rect 8668 47398 8720 47404
rect 8680 46986 8708 47398
rect 8668 46980 8720 46986
rect 8668 46922 8720 46928
rect 8576 46436 8628 46442
rect 8576 46378 8628 46384
rect 8772 46186 8800 47518
rect 8864 47122 8892 48078
rect 8852 47116 8904 47122
rect 8852 47058 8904 47064
rect 8852 46436 8904 46442
rect 8852 46378 8904 46384
rect 8588 46158 8800 46186
rect 8588 43382 8616 46158
rect 8668 46096 8720 46102
rect 8668 46038 8720 46044
rect 8576 43376 8628 43382
rect 8576 43318 8628 43324
rect 8576 43104 8628 43110
rect 8576 43046 8628 43052
rect 8588 42809 8616 43046
rect 8574 42800 8630 42809
rect 8574 42735 8630 42744
rect 8576 42628 8628 42634
rect 8576 42570 8628 42576
rect 8588 41546 8616 42570
rect 8576 41540 8628 41546
rect 8576 41482 8628 41488
rect 8496 41386 8616 41414
rect 8482 41304 8538 41313
rect 8482 41239 8538 41248
rect 8392 37460 8444 37466
rect 8392 37402 8444 37408
rect 8312 37318 8432 37346
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 8312 22098 8340 37198
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8312 19514 8340 20266
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8312 18601 8340 19314
rect 8298 18592 8354 18601
rect 8298 18527 8354 18536
rect 8404 18465 8432 37318
rect 8496 37262 8524 41239
rect 8588 40934 8616 41386
rect 8576 40928 8628 40934
rect 8576 40870 8628 40876
rect 8574 40760 8630 40769
rect 8574 40695 8630 40704
rect 8588 40118 8616 40695
rect 8576 40112 8628 40118
rect 8576 40054 8628 40060
rect 8680 39930 8708 46038
rect 8760 45348 8812 45354
rect 8760 45290 8812 45296
rect 8772 41585 8800 45290
rect 8758 41576 8814 41585
rect 8758 41511 8814 41520
rect 8760 41472 8812 41478
rect 8760 41414 8812 41420
rect 8864 41414 8892 46378
rect 8956 41750 8984 48606
rect 9109 48444 9417 48464
rect 9109 48442 9115 48444
rect 9171 48442 9195 48444
rect 9251 48442 9275 48444
rect 9331 48442 9355 48444
rect 9411 48442 9417 48444
rect 9171 48390 9173 48442
rect 9353 48390 9355 48442
rect 9109 48388 9115 48390
rect 9171 48388 9195 48390
rect 9251 48388 9275 48390
rect 9331 48388 9355 48390
rect 9411 48388 9417 48390
rect 9109 48368 9417 48388
rect 9036 48340 9088 48346
rect 9088 48288 9168 48314
rect 9036 48286 9168 48288
rect 9036 48282 9088 48286
rect 9036 48204 9088 48210
rect 9036 48146 9088 48152
rect 8944 41744 8996 41750
rect 8944 41686 8996 41692
rect 8588 39902 8708 39930
rect 8588 37618 8616 39902
rect 8668 39840 8720 39846
rect 8668 39782 8720 39788
rect 8680 39409 8708 39782
rect 8666 39400 8722 39409
rect 8666 39335 8722 39344
rect 8668 39024 8720 39030
rect 8668 38966 8720 38972
rect 8680 37874 8708 38966
rect 8668 37868 8720 37874
rect 8668 37810 8720 37816
rect 8588 37590 8708 37618
rect 8576 37460 8628 37466
rect 8576 37402 8628 37408
rect 8484 37256 8536 37262
rect 8484 37198 8536 37204
rect 8484 37120 8536 37126
rect 8484 37062 8536 37068
rect 8496 33300 8524 37062
rect 8588 33425 8616 37402
rect 8680 34610 8708 37590
rect 8772 34898 8800 41414
rect 8864 41386 8984 41414
rect 8852 40996 8904 41002
rect 8852 40938 8904 40944
rect 8864 36922 8892 40938
rect 8852 36916 8904 36922
rect 8852 36858 8904 36864
rect 8852 36576 8904 36582
rect 8852 36518 8904 36524
rect 8864 36145 8892 36518
rect 8850 36136 8906 36145
rect 8850 36071 8906 36080
rect 8852 36032 8904 36038
rect 8850 36000 8852 36009
rect 8904 36000 8906 36009
rect 8850 35935 8906 35944
rect 8850 35592 8906 35601
rect 8850 35527 8906 35536
rect 8864 35290 8892 35527
rect 8852 35284 8904 35290
rect 8852 35226 8904 35232
rect 8772 34870 8892 34898
rect 8864 34728 8892 34870
rect 8772 34700 8892 34728
rect 8668 34604 8720 34610
rect 8668 34546 8720 34552
rect 8666 34504 8722 34513
rect 8666 34439 8722 34448
rect 8680 33522 8708 34439
rect 8668 33516 8720 33522
rect 8668 33458 8720 33464
rect 8574 33416 8630 33425
rect 8574 33351 8630 33360
rect 8496 33272 8708 33300
rect 8574 33144 8630 33153
rect 8484 33108 8536 33114
rect 8574 33079 8630 33088
rect 8484 33050 8536 33056
rect 8496 25906 8524 33050
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 8496 20942 8524 25094
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8390 18456 8446 18465
rect 8390 18391 8446 18400
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8312 15638 8340 17138
rect 8404 16454 8432 18226
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8496 16266 8524 16594
rect 8404 16238 8524 16266
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8312 15094 8340 15438
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8404 14958 8432 16238
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8298 14784 8354 14793
rect 8298 14719 8354 14728
rect 8312 14346 8340 14719
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8404 14226 8432 14894
rect 8312 14198 8432 14226
rect 8312 13852 8340 14198
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8404 13977 8432 14010
rect 8390 13968 8446 13977
rect 8390 13903 8446 13912
rect 8312 13824 8432 13852
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8312 13462 8340 13670
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8404 13308 8432 13824
rect 8312 13280 8432 13308
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8128 11150 8156 11494
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7477 10908 7785 10928
rect 7477 10906 7483 10908
rect 7539 10906 7563 10908
rect 7619 10906 7643 10908
rect 7699 10906 7723 10908
rect 7779 10906 7785 10908
rect 7539 10854 7541 10906
rect 7721 10854 7723 10906
rect 7477 10852 7483 10854
rect 7539 10852 7563 10854
rect 7619 10852 7643 10854
rect 7699 10852 7723 10854
rect 7779 10852 7785 10854
rect 7477 10832 7785 10852
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7116 10062 7144 10474
rect 7208 10266 7236 10610
rect 8036 10577 8064 10610
rect 8022 10568 8078 10577
rect 8022 10503 8078 10512
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 4213 5468 4521 5488
rect 4213 5466 4219 5468
rect 4275 5466 4299 5468
rect 4355 5466 4379 5468
rect 4435 5466 4459 5468
rect 4515 5466 4521 5468
rect 4275 5414 4277 5466
rect 4457 5414 4459 5466
rect 4213 5412 4219 5414
rect 4275 5412 4299 5414
rect 4355 5412 4379 5414
rect 4435 5412 4459 5414
rect 4515 5412 4521 5414
rect 4213 5392 4521 5412
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 1584 5024 1636 5030
rect 1582 4992 1584 5001
rect 1636 4992 1638 5001
rect 1582 4927 1638 4936
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 1412 4678 1532 4706
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 1601 1440 2790
rect 1504 2446 1532 4678
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4321 1624 4422
rect 4213 4380 4521 4400
rect 4213 4378 4219 4380
rect 4275 4378 4299 4380
rect 4355 4378 4379 4380
rect 4435 4378 4459 4380
rect 4515 4378 4521 4380
rect 4275 4326 4277 4378
rect 4457 4326 4459 4378
rect 4213 4324 4219 4326
rect 4275 4324 4299 4326
rect 4355 4324 4379 4326
rect 4435 4324 4459 4326
rect 4515 4324 4521 4326
rect 1582 4312 1638 4321
rect 4213 4304 4521 4324
rect 1582 4247 1638 4256
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3641 1624 3878
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 2961 1624 3334
rect 4213 3292 4521 3312
rect 4213 3290 4219 3292
rect 4275 3290 4299 3292
rect 4355 3290 4379 3292
rect 4435 3290 4459 3292
rect 4515 3290 4521 3292
rect 4275 3238 4277 3290
rect 4457 3238 4459 3290
rect 4213 3236 4219 3238
rect 4275 3236 4299 3238
rect 4355 3236 4379 3238
rect 4435 3236 4459 3238
rect 4515 3236 4521 3238
rect 4213 3216 4521 3236
rect 1582 2952 1638 2961
rect 1582 2887 1638 2896
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 5552 2514 5580 5034
rect 5845 4924 6153 4944
rect 5845 4922 5851 4924
rect 5907 4922 5931 4924
rect 5987 4922 6011 4924
rect 6067 4922 6091 4924
rect 6147 4922 6153 4924
rect 5907 4870 5909 4922
rect 6089 4870 6091 4922
rect 5845 4868 5851 4870
rect 5907 4868 5931 4870
rect 5987 4868 6011 4870
rect 6067 4868 6091 4870
rect 6147 4868 6153 4870
rect 5845 4848 6153 4868
rect 5845 3836 6153 3856
rect 5845 3834 5851 3836
rect 5907 3834 5931 3836
rect 5987 3834 6011 3836
rect 6067 3834 6091 3836
rect 6147 3834 6153 3836
rect 5907 3782 5909 3834
rect 6089 3782 6091 3834
rect 5845 3780 5851 3782
rect 5907 3780 5931 3782
rect 5987 3780 6011 3782
rect 6067 3780 6091 3782
rect 6147 3780 6153 3782
rect 5845 3760 6153 3780
rect 5845 2748 6153 2768
rect 5845 2746 5851 2748
rect 5907 2746 5931 2748
rect 5987 2746 6011 2748
rect 6067 2746 6091 2748
rect 6147 2746 6153 2748
rect 5907 2694 5909 2746
rect 6089 2694 6091 2746
rect 5845 2692 5851 2694
rect 5907 2692 5931 2694
rect 5987 2692 6011 2694
rect 6067 2692 6091 2694
rect 6147 2692 6153 2694
rect 5845 2672 6153 2692
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 7116 2446 7144 9998
rect 7477 9820 7785 9840
rect 7477 9818 7483 9820
rect 7539 9818 7563 9820
rect 7619 9818 7643 9820
rect 7699 9818 7723 9820
rect 7779 9818 7785 9820
rect 7539 9766 7541 9818
rect 7721 9766 7723 9818
rect 7477 9764 7483 9766
rect 7539 9764 7563 9766
rect 7619 9764 7643 9766
rect 7699 9764 7723 9766
rect 7779 9764 7785 9766
rect 7477 9744 7785 9764
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 9489 7880 9522
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7477 8732 7785 8752
rect 7477 8730 7483 8732
rect 7539 8730 7563 8732
rect 7619 8730 7643 8732
rect 7699 8730 7723 8732
rect 7779 8730 7785 8732
rect 7539 8678 7541 8730
rect 7721 8678 7723 8730
rect 7477 8676 7483 8678
rect 7539 8676 7563 8678
rect 7619 8676 7643 8678
rect 7699 8676 7723 8678
rect 7779 8676 7785 8678
rect 7477 8656 7785 8676
rect 7477 7644 7785 7664
rect 7477 7642 7483 7644
rect 7539 7642 7563 7644
rect 7619 7642 7643 7644
rect 7699 7642 7723 7644
rect 7779 7642 7785 7644
rect 7539 7590 7541 7642
rect 7721 7590 7723 7642
rect 7477 7588 7483 7590
rect 7539 7588 7563 7590
rect 7619 7588 7643 7590
rect 7699 7588 7723 7590
rect 7779 7588 7785 7590
rect 7477 7568 7785 7588
rect 7477 6556 7785 6576
rect 7477 6554 7483 6556
rect 7539 6554 7563 6556
rect 7619 6554 7643 6556
rect 7699 6554 7723 6556
rect 7779 6554 7785 6556
rect 7539 6502 7541 6554
rect 7721 6502 7723 6554
rect 7477 6500 7483 6502
rect 7539 6500 7563 6502
rect 7619 6500 7643 6502
rect 7699 6500 7723 6502
rect 7779 6500 7785 6502
rect 7477 6480 7785 6500
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7477 5468 7785 5488
rect 7477 5466 7483 5468
rect 7539 5466 7563 5468
rect 7619 5466 7643 5468
rect 7699 5466 7723 5468
rect 7779 5466 7785 5468
rect 7539 5414 7541 5466
rect 7721 5414 7723 5466
rect 7477 5412 7483 5414
rect 7539 5412 7563 5414
rect 7619 5412 7643 5414
rect 7699 5412 7723 5414
rect 7779 5412 7785 5414
rect 7477 5392 7785 5412
rect 7477 4380 7785 4400
rect 7477 4378 7483 4380
rect 7539 4378 7563 4380
rect 7619 4378 7643 4380
rect 7699 4378 7723 4380
rect 7779 4378 7785 4380
rect 7539 4326 7541 4378
rect 7721 4326 7723 4378
rect 7477 4324 7483 4326
rect 7539 4324 7563 4326
rect 7619 4324 7643 4326
rect 7699 4324 7723 4326
rect 7779 4324 7785 4326
rect 7477 4304 7785 4324
rect 8036 4282 8064 5646
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8128 5137 8156 5170
rect 8114 5128 8170 5137
rect 8114 5063 8170 5072
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8116 3528 8168 3534
rect 8114 3496 8116 3505
rect 8168 3496 8170 3505
rect 8114 3431 8170 3440
rect 7477 3292 7785 3312
rect 7477 3290 7483 3292
rect 7539 3290 7563 3292
rect 7619 3290 7643 3292
rect 7699 3290 7723 3292
rect 7779 3290 7785 3292
rect 7539 3238 7541 3290
rect 7721 3238 7723 3290
rect 7477 3236 7483 3238
rect 7539 3236 7563 3238
rect 7619 3236 7643 3238
rect 7699 3236 7723 3238
rect 7779 3236 7785 3238
rect 7477 3216 7785 3236
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7838 2952 7894 2961
rect 7838 2887 7840 2896
rect 7892 2887 7894 2896
rect 7840 2858 7892 2864
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 1584 2304 1636 2310
rect 2320 2304 2372 2310
rect 1584 2246 1636 2252
rect 2318 2272 2320 2281
rect 2872 2304 2924 2310
rect 2372 2272 2374 2281
rect 1398 1592 1454 1601
rect 1398 1527 1454 1536
rect 1596 921 1624 2246
rect 2872 2246 2924 2252
rect 2318 2207 2374 2216
rect 1582 912 1638 921
rect 1582 847 1638 856
rect 2884 377 2912 2246
rect 4213 2204 4521 2224
rect 4213 2202 4219 2204
rect 4275 2202 4299 2204
rect 4355 2202 4379 2204
rect 4435 2202 4459 2204
rect 4515 2202 4521 2204
rect 4275 2150 4277 2202
rect 4457 2150 4459 2202
rect 4213 2148 4219 2150
rect 4275 2148 4299 2150
rect 4355 2148 4379 2150
rect 4435 2148 4459 2150
rect 4515 2148 4521 2150
rect 4213 2128 4521 2148
rect 7477 2204 7785 2224
rect 7477 2202 7483 2204
rect 7539 2202 7563 2204
rect 7619 2202 7643 2204
rect 7699 2202 7723 2204
rect 7779 2202 7785 2204
rect 7539 2150 7541 2202
rect 7721 2150 7723 2202
rect 7477 2148 7483 2150
rect 7539 2148 7563 2150
rect 7619 2148 7643 2150
rect 7699 2148 7723 2150
rect 7779 2148 7785 2150
rect 7477 2128 7785 2148
rect 7944 1601 7972 2450
rect 7930 1592 7986 1601
rect 7930 1527 7986 1536
rect 2870 368 2926 377
rect 2870 303 2926 312
rect 8128 241 8156 2994
rect 8220 649 8248 11698
rect 8312 2922 8340 13280
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 8404 11898 8432 12106
rect 8496 11898 8524 14962
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8390 11112 8446 11121
rect 8390 11047 8446 11056
rect 8404 10062 8432 11047
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8496 9654 8524 11834
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8404 4622 8432 7210
rect 8588 7206 8616 33079
rect 8680 28558 8708 33272
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8680 20534 8708 26930
rect 8772 23866 8800 34700
rect 8852 34604 8904 34610
rect 8852 34546 8904 34552
rect 8864 32978 8892 34546
rect 8852 32972 8904 32978
rect 8852 32914 8904 32920
rect 8852 32224 8904 32230
rect 8852 32166 8904 32172
rect 8864 31929 8892 32166
rect 8850 31920 8906 31929
rect 8850 31855 8906 31864
rect 8852 31136 8904 31142
rect 8852 31078 8904 31084
rect 8864 27062 8892 31078
rect 8852 27056 8904 27062
rect 8852 26998 8904 27004
rect 8956 26994 8984 41386
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 9048 26874 9076 48146
rect 9140 47569 9168 48286
rect 9508 48142 9536 48826
rect 9600 48278 9628 49150
rect 9968 48754 9996 49694
rect 9956 48748 10008 48754
rect 9956 48690 10008 48696
rect 9588 48272 9640 48278
rect 9588 48214 9640 48220
rect 9968 48142 9996 48690
rect 9496 48136 9548 48142
rect 9496 48078 9548 48084
rect 9956 48136 10008 48142
rect 9956 48078 10008 48084
rect 9680 48000 9732 48006
rect 9680 47942 9732 47948
rect 9220 47796 9272 47802
rect 9220 47738 9272 47744
rect 9232 47705 9260 47738
rect 9692 47734 9720 47942
rect 9680 47728 9732 47734
rect 9218 47696 9274 47705
rect 9680 47670 9732 47676
rect 9218 47631 9274 47640
rect 9588 47660 9640 47666
rect 9588 47602 9640 47608
rect 9864 47660 9916 47666
rect 9864 47602 9916 47608
rect 9496 47592 9548 47598
rect 9126 47560 9182 47569
rect 9496 47534 9548 47540
rect 9126 47495 9182 47504
rect 9508 47433 9536 47534
rect 9494 47424 9550 47433
rect 9109 47356 9417 47376
rect 9494 47359 9550 47368
rect 9109 47354 9115 47356
rect 9171 47354 9195 47356
rect 9251 47354 9275 47356
rect 9331 47354 9355 47356
rect 9411 47354 9417 47356
rect 9171 47302 9173 47354
rect 9353 47302 9355 47354
rect 9109 47300 9115 47302
rect 9171 47300 9195 47302
rect 9251 47300 9275 47302
rect 9331 47300 9355 47302
rect 9411 47300 9417 47302
rect 9109 47280 9417 47300
rect 9404 47116 9456 47122
rect 9404 47058 9456 47064
rect 9416 46510 9444 47058
rect 9600 46617 9628 47602
rect 9772 47184 9824 47190
rect 9772 47126 9824 47132
rect 9680 46912 9732 46918
rect 9680 46854 9732 46860
rect 9586 46608 9642 46617
rect 9586 46543 9642 46552
rect 9404 46504 9456 46510
rect 9496 46504 9548 46510
rect 9404 46446 9456 46452
rect 9494 46472 9496 46481
rect 9548 46472 9550 46481
rect 9494 46407 9550 46416
rect 9588 46436 9640 46442
rect 9588 46378 9640 46384
rect 9109 46268 9417 46288
rect 9109 46266 9115 46268
rect 9171 46266 9195 46268
rect 9251 46266 9275 46268
rect 9331 46266 9355 46268
rect 9411 46266 9417 46268
rect 9171 46214 9173 46266
rect 9353 46214 9355 46266
rect 9109 46212 9115 46214
rect 9171 46212 9195 46214
rect 9251 46212 9275 46214
rect 9331 46212 9355 46214
rect 9411 46212 9417 46214
rect 9109 46192 9417 46212
rect 9494 46200 9550 46209
rect 9494 46135 9550 46144
rect 9109 45180 9417 45200
rect 9109 45178 9115 45180
rect 9171 45178 9195 45180
rect 9251 45178 9275 45180
rect 9331 45178 9355 45180
rect 9411 45178 9417 45180
rect 9171 45126 9173 45178
rect 9353 45126 9355 45178
rect 9109 45124 9115 45126
rect 9171 45124 9195 45126
rect 9251 45124 9275 45126
rect 9331 45124 9355 45126
rect 9411 45124 9417 45126
rect 9109 45104 9417 45124
rect 9404 44872 9456 44878
rect 9402 44840 9404 44849
rect 9508 44860 9536 46135
rect 9600 46034 9628 46378
rect 9588 46028 9640 46034
rect 9588 45970 9640 45976
rect 9588 45892 9640 45898
rect 9588 45834 9640 45840
rect 9600 45354 9628 45834
rect 9588 45348 9640 45354
rect 9588 45290 9640 45296
rect 9588 45076 9640 45082
rect 9588 45018 9640 45024
rect 9456 44840 9536 44860
rect 9458 44832 9536 44840
rect 9600 44792 9628 45018
rect 9402 44775 9458 44784
rect 9508 44764 9628 44792
rect 9402 44568 9458 44577
rect 9508 44554 9536 44764
rect 9458 44526 9536 44554
rect 9588 44532 9640 44538
rect 9402 44503 9458 44512
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9232 44305 9260 44338
rect 9416 44334 9444 44503
rect 9588 44474 9640 44480
rect 9404 44328 9456 44334
rect 9218 44296 9274 44305
rect 9404 44270 9456 44276
rect 9218 44231 9274 44240
rect 9109 44092 9417 44112
rect 9109 44090 9115 44092
rect 9171 44090 9195 44092
rect 9251 44090 9275 44092
rect 9331 44090 9355 44092
rect 9411 44090 9417 44092
rect 9171 44038 9173 44090
rect 9353 44038 9355 44090
rect 9109 44036 9115 44038
rect 9171 44036 9195 44038
rect 9251 44036 9275 44038
rect 9331 44036 9355 44038
rect 9411 44036 9417 44038
rect 9109 44016 9417 44036
rect 9600 43976 9628 44474
rect 9508 43948 9628 43976
rect 9126 43752 9182 43761
rect 9126 43687 9182 43696
rect 9140 43314 9168 43687
rect 9128 43308 9180 43314
rect 9128 43250 9180 43256
rect 9109 43004 9417 43024
rect 9109 43002 9115 43004
rect 9171 43002 9195 43004
rect 9251 43002 9275 43004
rect 9331 43002 9355 43004
rect 9411 43002 9417 43004
rect 9171 42950 9173 43002
rect 9353 42950 9355 43002
rect 9109 42948 9115 42950
rect 9171 42948 9195 42950
rect 9251 42948 9275 42950
rect 9331 42948 9355 42950
rect 9411 42948 9417 42950
rect 9109 42928 9417 42948
rect 9126 42256 9182 42265
rect 9126 42191 9128 42200
rect 9180 42191 9182 42200
rect 9128 42162 9180 42168
rect 9109 41916 9417 41936
rect 9109 41914 9115 41916
rect 9171 41914 9195 41916
rect 9251 41914 9275 41916
rect 9331 41914 9355 41916
rect 9411 41914 9417 41916
rect 9171 41862 9173 41914
rect 9353 41862 9355 41914
rect 9109 41860 9115 41862
rect 9171 41860 9195 41862
rect 9251 41860 9275 41862
rect 9331 41860 9355 41862
rect 9411 41860 9417 41862
rect 9109 41840 9417 41860
rect 9404 41744 9456 41750
rect 9404 41686 9456 41692
rect 9416 41002 9444 41686
rect 9508 41070 9536 43948
rect 9586 43888 9642 43897
rect 9586 43823 9642 43832
rect 9496 41064 9548 41070
rect 9496 41006 9548 41012
rect 9404 40996 9456 41002
rect 9404 40938 9456 40944
rect 9496 40928 9548 40934
rect 9496 40870 9548 40876
rect 9109 40828 9417 40848
rect 9109 40826 9115 40828
rect 9171 40826 9195 40828
rect 9251 40826 9275 40828
rect 9331 40826 9355 40828
rect 9411 40826 9417 40828
rect 9171 40774 9173 40826
rect 9353 40774 9355 40826
rect 9109 40772 9115 40774
rect 9171 40772 9195 40774
rect 9251 40772 9275 40774
rect 9331 40772 9355 40774
rect 9411 40772 9417 40774
rect 9109 40752 9417 40772
rect 9128 40656 9180 40662
rect 9128 40598 9180 40604
rect 9140 39914 9168 40598
rect 9312 40384 9364 40390
rect 9312 40326 9364 40332
rect 9324 39953 9352 40326
rect 9310 39944 9366 39953
rect 9128 39908 9180 39914
rect 9310 39879 9366 39888
rect 9128 39850 9180 39856
rect 9109 39740 9417 39760
rect 9109 39738 9115 39740
rect 9171 39738 9195 39740
rect 9251 39738 9275 39740
rect 9331 39738 9355 39740
rect 9411 39738 9417 39740
rect 9171 39686 9173 39738
rect 9353 39686 9355 39738
rect 9109 39684 9115 39686
rect 9171 39684 9195 39686
rect 9251 39684 9275 39686
rect 9331 39684 9355 39686
rect 9411 39684 9417 39686
rect 9109 39664 9417 39684
rect 9402 39536 9458 39545
rect 9508 39506 9536 40870
rect 9402 39471 9458 39480
rect 9496 39500 9548 39506
rect 9416 39370 9444 39471
rect 9496 39442 9548 39448
rect 9404 39364 9456 39370
rect 9404 39306 9456 39312
rect 9496 38888 9548 38894
rect 9126 38856 9182 38865
rect 9496 38830 9548 38836
rect 9126 38791 9128 38800
rect 9180 38791 9182 38800
rect 9128 38762 9180 38768
rect 9109 38652 9417 38672
rect 9109 38650 9115 38652
rect 9171 38650 9195 38652
rect 9251 38650 9275 38652
rect 9331 38650 9355 38652
rect 9411 38650 9417 38652
rect 9171 38598 9173 38650
rect 9353 38598 9355 38650
rect 9109 38596 9115 38598
rect 9171 38596 9195 38598
rect 9251 38596 9275 38598
rect 9331 38596 9355 38598
rect 9411 38596 9417 38598
rect 9109 38576 9417 38596
rect 9312 38480 9364 38486
rect 9312 38422 9364 38428
rect 9126 38312 9182 38321
rect 9126 38247 9182 38256
rect 9140 37738 9168 38247
rect 9220 38208 9272 38214
rect 9218 38176 9220 38185
rect 9272 38176 9274 38185
rect 9218 38111 9274 38120
rect 9324 37913 9352 38422
rect 9508 38010 9536 38830
rect 9600 38554 9628 43823
rect 9692 43654 9720 46854
rect 9784 46714 9812 47126
rect 9772 46708 9824 46714
rect 9772 46650 9824 46656
rect 9784 44946 9812 46650
rect 9876 45082 9904 47602
rect 9968 47598 9996 48078
rect 10060 47802 10088 51750
rect 10048 47796 10100 47802
rect 10048 47738 10100 47744
rect 9956 47592 10008 47598
rect 9956 47534 10008 47540
rect 9968 47122 9996 47534
rect 10048 47456 10100 47462
rect 10048 47398 10100 47404
rect 9956 47116 10008 47122
rect 9956 47058 10008 47064
rect 9956 46368 10008 46374
rect 9954 46336 9956 46345
rect 10008 46336 10010 46345
rect 9954 46271 10010 46280
rect 9956 45824 10008 45830
rect 9956 45766 10008 45772
rect 9968 45626 9996 45766
rect 9956 45620 10008 45626
rect 9956 45562 10008 45568
rect 10060 45558 10088 47398
rect 10048 45552 10100 45558
rect 10048 45494 10100 45500
rect 9864 45076 9916 45082
rect 9864 45018 9916 45024
rect 10152 44962 10180 53382
rect 10244 53038 10272 53502
rect 10232 53032 10284 53038
rect 10232 52974 10284 52980
rect 10244 51474 10272 52974
rect 10232 51468 10284 51474
rect 10232 51410 10284 51416
rect 10244 50862 10272 51410
rect 10232 50856 10284 50862
rect 10232 50798 10284 50804
rect 10232 47660 10284 47666
rect 10232 47602 10284 47608
rect 10244 46345 10272 47602
rect 10230 46336 10286 46345
rect 10230 46271 10286 46280
rect 10232 46164 10284 46170
rect 10232 46106 10284 46112
rect 9772 44940 9824 44946
rect 9772 44882 9824 44888
rect 9876 44934 10180 44962
rect 9876 44826 9904 44934
rect 9784 44798 9904 44826
rect 9956 44872 10008 44878
rect 9956 44814 10008 44820
rect 9680 43648 9732 43654
rect 9680 43590 9732 43596
rect 9680 43444 9732 43450
rect 9680 43386 9732 43392
rect 9588 38548 9640 38554
rect 9588 38490 9640 38496
rect 9588 38412 9640 38418
rect 9588 38354 9640 38360
rect 9496 38004 9548 38010
rect 9496 37946 9548 37952
rect 9310 37904 9366 37913
rect 9310 37839 9366 37848
rect 9600 37806 9628 38354
rect 9692 38298 9720 43386
rect 9784 38593 9812 44798
rect 9862 44432 9918 44441
rect 9968 44402 9996 44814
rect 10140 44804 10192 44810
rect 10140 44746 10192 44752
rect 10152 44538 10180 44746
rect 10140 44532 10192 44538
rect 10140 44474 10192 44480
rect 9862 44367 9918 44376
rect 9956 44396 10008 44402
rect 9876 43450 9904 44367
rect 9956 44338 10008 44344
rect 10048 44328 10100 44334
rect 10048 44270 10100 44276
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9864 43308 9916 43314
rect 9864 43250 9916 43256
rect 9956 43308 10008 43314
rect 9956 43250 10008 43256
rect 9876 43217 9904 43250
rect 9862 43208 9918 43217
rect 9862 43143 9918 43152
rect 9968 42634 9996 43250
rect 9956 42628 10008 42634
rect 9956 42570 10008 42576
rect 9956 42220 10008 42226
rect 9956 42162 10008 42168
rect 9968 41857 9996 42162
rect 9954 41848 10010 41857
rect 9954 41783 10010 41792
rect 9864 41608 9916 41614
rect 9864 41550 9916 41556
rect 9876 40526 9904 41550
rect 9956 41540 10008 41546
rect 9956 41482 10008 41488
rect 9968 41313 9996 41482
rect 9954 41304 10010 41313
rect 9954 41239 10010 41248
rect 9956 41132 10008 41138
rect 9956 41074 10008 41080
rect 9968 40905 9996 41074
rect 9954 40896 10010 40905
rect 9954 40831 10010 40840
rect 9864 40520 9916 40526
rect 10060 40474 10088 44270
rect 10140 43716 10192 43722
rect 10140 43658 10192 43664
rect 10152 43178 10180 43658
rect 10140 43172 10192 43178
rect 10140 43114 10192 43120
rect 10140 42832 10192 42838
rect 10140 42774 10192 42780
rect 10152 42673 10180 42774
rect 10138 42664 10194 42673
rect 10138 42599 10194 42608
rect 10138 42392 10194 42401
rect 10138 42327 10194 42336
rect 10152 42226 10180 42327
rect 10140 42220 10192 42226
rect 10140 42162 10192 42168
rect 10138 42120 10194 42129
rect 10138 42055 10194 42064
rect 10152 41682 10180 42055
rect 10140 41676 10192 41682
rect 10140 41618 10192 41624
rect 10140 41540 10192 41546
rect 10140 41482 10192 41488
rect 10152 40594 10180 41482
rect 10140 40588 10192 40594
rect 10140 40530 10192 40536
rect 9864 40462 9916 40468
rect 9968 40446 10088 40474
rect 10138 40488 10194 40497
rect 9864 40112 9916 40118
rect 9864 40054 9916 40060
rect 9876 39681 9904 40054
rect 9862 39672 9918 39681
rect 9968 39642 9996 40446
rect 10138 40423 10194 40432
rect 10048 40384 10100 40390
rect 10048 40326 10100 40332
rect 9862 39607 9918 39616
rect 9956 39636 10008 39642
rect 9956 39578 10008 39584
rect 9956 39500 10008 39506
rect 9956 39442 10008 39448
rect 9864 39296 9916 39302
rect 9864 39238 9916 39244
rect 9770 38584 9826 38593
rect 9770 38519 9826 38528
rect 9692 38270 9812 38298
rect 9588 37800 9640 37806
rect 9640 37760 9720 37788
rect 9588 37742 9640 37748
rect 9128 37732 9180 37738
rect 9128 37674 9180 37680
rect 9588 37664 9640 37670
rect 9588 37606 9640 37612
rect 9109 37564 9417 37584
rect 9109 37562 9115 37564
rect 9171 37562 9195 37564
rect 9251 37562 9275 37564
rect 9331 37562 9355 37564
rect 9411 37562 9417 37564
rect 9171 37510 9173 37562
rect 9353 37510 9355 37562
rect 9109 37508 9115 37510
rect 9171 37508 9195 37510
rect 9251 37508 9275 37510
rect 9331 37508 9355 37510
rect 9411 37508 9417 37510
rect 9109 37488 9417 37508
rect 9600 37505 9628 37606
rect 9586 37496 9642 37505
rect 9586 37431 9642 37440
rect 9692 37330 9720 37760
rect 9680 37324 9732 37330
rect 9600 37272 9680 37274
rect 9600 37266 9732 37272
rect 9600 37246 9720 37266
rect 9600 36854 9628 37246
rect 9588 36848 9640 36854
rect 9588 36790 9640 36796
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9496 36576 9548 36582
rect 9496 36518 9548 36524
rect 9109 36476 9417 36496
rect 9109 36474 9115 36476
rect 9171 36474 9195 36476
rect 9251 36474 9275 36476
rect 9331 36474 9355 36476
rect 9411 36474 9417 36476
rect 9171 36422 9173 36474
rect 9353 36422 9355 36474
rect 9109 36420 9115 36422
rect 9171 36420 9195 36422
rect 9251 36420 9275 36422
rect 9331 36420 9355 36422
rect 9411 36420 9417 36422
rect 9109 36400 9417 36420
rect 9402 36272 9458 36281
rect 9402 36207 9404 36216
rect 9456 36207 9458 36216
rect 9404 36178 9456 36184
rect 9109 35388 9417 35408
rect 9109 35386 9115 35388
rect 9171 35386 9195 35388
rect 9251 35386 9275 35388
rect 9331 35386 9355 35388
rect 9411 35386 9417 35388
rect 9171 35334 9173 35386
rect 9353 35334 9355 35386
rect 9109 35332 9115 35334
rect 9171 35332 9195 35334
rect 9251 35332 9275 35334
rect 9331 35332 9355 35334
rect 9411 35332 9417 35334
rect 9109 35312 9417 35332
rect 9312 35148 9364 35154
rect 9312 35090 9364 35096
rect 9324 34678 9352 35090
rect 9312 34672 9364 34678
rect 9312 34614 9364 34620
rect 9109 34300 9417 34320
rect 9109 34298 9115 34300
rect 9171 34298 9195 34300
rect 9251 34298 9275 34300
rect 9331 34298 9355 34300
rect 9411 34298 9417 34300
rect 9171 34246 9173 34298
rect 9353 34246 9355 34298
rect 9109 34244 9115 34246
rect 9171 34244 9195 34246
rect 9251 34244 9275 34246
rect 9331 34244 9355 34246
rect 9411 34244 9417 34246
rect 9109 34224 9417 34244
rect 9312 33856 9364 33862
rect 9310 33824 9312 33833
rect 9364 33824 9366 33833
rect 9310 33759 9366 33768
rect 9109 33212 9417 33232
rect 9109 33210 9115 33212
rect 9171 33210 9195 33212
rect 9251 33210 9275 33212
rect 9331 33210 9355 33212
rect 9411 33210 9417 33212
rect 9171 33158 9173 33210
rect 9353 33158 9355 33210
rect 9109 33156 9115 33158
rect 9171 33156 9195 33158
rect 9251 33156 9275 33158
rect 9331 33156 9355 33158
rect 9411 33156 9417 33158
rect 9109 33136 9417 33156
rect 9508 32842 9536 36518
rect 9692 36242 9720 36790
rect 9588 36236 9640 36242
rect 9588 36178 9640 36184
rect 9680 36236 9732 36242
rect 9680 36178 9732 36184
rect 9600 34474 9628 36178
rect 9784 35086 9812 38270
rect 9876 37126 9904 39238
rect 9968 38162 9996 39442
rect 10060 39001 10088 40326
rect 10152 40050 10180 40423
rect 10140 40044 10192 40050
rect 10140 39986 10192 39992
rect 10140 39432 10192 39438
rect 10140 39374 10192 39380
rect 10046 38992 10102 39001
rect 10046 38927 10102 38936
rect 10048 38888 10100 38894
rect 10048 38830 10100 38836
rect 10060 38418 10088 38830
rect 10048 38412 10100 38418
rect 10048 38354 10100 38360
rect 9968 38134 10088 38162
rect 9956 37936 10008 37942
rect 9956 37878 10008 37884
rect 9864 37120 9916 37126
rect 9864 37062 9916 37068
rect 9864 35828 9916 35834
rect 9864 35770 9916 35776
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9588 34468 9640 34474
rect 9588 34410 9640 34416
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9586 33552 9642 33561
rect 9642 33510 9720 33538
rect 9586 33487 9642 33496
rect 9588 33380 9640 33386
rect 9588 33322 9640 33328
rect 9600 33289 9628 33322
rect 9586 33280 9642 33289
rect 9586 33215 9642 33224
rect 9692 33130 9720 33510
rect 9600 33102 9720 33130
rect 9496 32836 9548 32842
rect 9496 32778 9548 32784
rect 9220 32768 9272 32774
rect 9220 32710 9272 32716
rect 9404 32768 9456 32774
rect 9404 32710 9456 32716
rect 9232 32337 9260 32710
rect 9416 32366 9444 32710
rect 9404 32360 9456 32366
rect 9218 32328 9274 32337
rect 9404 32302 9456 32308
rect 9218 32263 9274 32272
rect 9416 32212 9444 32302
rect 9416 32184 9536 32212
rect 9109 32124 9417 32144
rect 9109 32122 9115 32124
rect 9171 32122 9195 32124
rect 9251 32122 9275 32124
rect 9331 32122 9355 32124
rect 9411 32122 9417 32124
rect 9171 32070 9173 32122
rect 9353 32070 9355 32122
rect 9109 32068 9115 32070
rect 9171 32068 9195 32070
rect 9251 32068 9275 32070
rect 9331 32068 9355 32070
rect 9411 32068 9417 32070
rect 9109 32048 9417 32068
rect 9508 32008 9536 32184
rect 9416 31980 9536 32008
rect 9416 31226 9444 31980
rect 9416 31198 9536 31226
rect 9109 31036 9417 31056
rect 9109 31034 9115 31036
rect 9171 31034 9195 31036
rect 9251 31034 9275 31036
rect 9331 31034 9355 31036
rect 9411 31034 9417 31036
rect 9171 30982 9173 31034
rect 9353 30982 9355 31034
rect 9109 30980 9115 30982
rect 9171 30980 9195 30982
rect 9251 30980 9275 30982
rect 9331 30980 9355 30982
rect 9411 30980 9417 30982
rect 9109 30960 9417 30980
rect 9109 29948 9417 29968
rect 9109 29946 9115 29948
rect 9171 29946 9195 29948
rect 9251 29946 9275 29948
rect 9331 29946 9355 29948
rect 9411 29946 9417 29948
rect 9171 29894 9173 29946
rect 9353 29894 9355 29946
rect 9109 29892 9115 29894
rect 9171 29892 9195 29894
rect 9251 29892 9275 29894
rect 9331 29892 9355 29894
rect 9411 29892 9417 29894
rect 9109 29872 9417 29892
rect 9312 29504 9364 29510
rect 9310 29472 9312 29481
rect 9364 29472 9366 29481
rect 9310 29407 9366 29416
rect 9126 29064 9182 29073
rect 9126 28999 9128 29008
rect 9180 28999 9182 29008
rect 9128 28970 9180 28976
rect 9109 28860 9417 28880
rect 9109 28858 9115 28860
rect 9171 28858 9195 28860
rect 9251 28858 9275 28860
rect 9331 28858 9355 28860
rect 9411 28858 9417 28860
rect 9171 28806 9173 28858
rect 9353 28806 9355 28858
rect 9109 28804 9115 28806
rect 9171 28804 9195 28806
rect 9251 28804 9275 28806
rect 9331 28804 9355 28806
rect 9411 28804 9417 28806
rect 9109 28784 9417 28804
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 9324 28121 9352 28358
rect 9310 28112 9366 28121
rect 9310 28047 9366 28056
rect 9109 27772 9417 27792
rect 9109 27770 9115 27772
rect 9171 27770 9195 27772
rect 9251 27770 9275 27772
rect 9331 27770 9355 27772
rect 9411 27770 9417 27772
rect 9171 27718 9173 27770
rect 9353 27718 9355 27770
rect 9109 27716 9115 27718
rect 9171 27716 9195 27718
rect 9251 27716 9275 27718
rect 9331 27716 9355 27718
rect 9411 27716 9417 27718
rect 9109 27696 9417 27716
rect 8864 26846 9076 26874
rect 8760 23860 8812 23866
rect 8760 23802 8812 23808
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8772 22953 8800 23666
rect 8758 22944 8814 22953
rect 8758 22879 8814 22888
rect 8760 22568 8812 22574
rect 8760 22510 8812 22516
rect 8772 21486 8800 22510
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 8772 19990 8800 21286
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8680 17649 8708 18702
rect 8864 18426 8892 26846
rect 9036 26784 9088 26790
rect 9036 26726 9088 26732
rect 8944 26580 8996 26586
rect 8944 26522 8996 26528
rect 8956 20330 8984 26522
rect 9048 23118 9076 26726
rect 9109 26684 9417 26704
rect 9109 26682 9115 26684
rect 9171 26682 9195 26684
rect 9251 26682 9275 26684
rect 9331 26682 9355 26684
rect 9411 26682 9417 26684
rect 9171 26630 9173 26682
rect 9353 26630 9355 26682
rect 9109 26628 9115 26630
rect 9171 26628 9195 26630
rect 9251 26628 9275 26630
rect 9331 26628 9355 26630
rect 9411 26628 9417 26630
rect 9109 26608 9417 26628
rect 9508 26586 9536 31198
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9496 25696 9548 25702
rect 9494 25664 9496 25673
rect 9548 25664 9550 25673
rect 9109 25596 9417 25616
rect 9494 25599 9550 25608
rect 9109 25594 9115 25596
rect 9171 25594 9195 25596
rect 9251 25594 9275 25596
rect 9331 25594 9355 25596
rect 9411 25594 9417 25596
rect 9171 25542 9173 25594
rect 9353 25542 9355 25594
rect 9109 25540 9115 25542
rect 9171 25540 9195 25542
rect 9251 25540 9275 25542
rect 9331 25540 9355 25542
rect 9411 25540 9417 25542
rect 9109 25520 9417 25540
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9109 24508 9417 24528
rect 9109 24506 9115 24508
rect 9171 24506 9195 24508
rect 9251 24506 9275 24508
rect 9331 24506 9355 24508
rect 9411 24506 9417 24508
rect 9171 24454 9173 24506
rect 9353 24454 9355 24506
rect 9109 24452 9115 24454
rect 9171 24452 9195 24454
rect 9251 24452 9275 24454
rect 9331 24452 9355 24454
rect 9411 24452 9417 24454
rect 9109 24432 9417 24452
rect 9508 24313 9536 24754
rect 9494 24304 9550 24313
rect 9494 24239 9550 24248
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9140 23769 9168 24142
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 9126 23760 9182 23769
rect 9126 23695 9182 23704
rect 9109 23420 9417 23440
rect 9109 23418 9115 23420
rect 9171 23418 9195 23420
rect 9251 23418 9275 23420
rect 9331 23418 9355 23420
rect 9411 23418 9417 23420
rect 9171 23366 9173 23418
rect 9353 23366 9355 23418
rect 9109 23364 9115 23366
rect 9171 23364 9195 23366
rect 9251 23364 9275 23366
rect 9331 23364 9355 23366
rect 9411 23364 9417 23366
rect 9109 23344 9417 23364
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 9109 22332 9417 22352
rect 9109 22330 9115 22332
rect 9171 22330 9195 22332
rect 9251 22330 9275 22332
rect 9331 22330 9355 22332
rect 9411 22330 9417 22332
rect 9171 22278 9173 22330
rect 9353 22278 9355 22330
rect 9109 22276 9115 22278
rect 9171 22276 9195 22278
rect 9251 22276 9275 22278
rect 9331 22276 9355 22278
rect 9411 22276 9417 22278
rect 9109 22256 9417 22276
rect 9508 22094 9536 24074
rect 9048 22066 9536 22094
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 9048 19530 9076 22066
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9324 21457 9352 21966
rect 9496 21480 9548 21486
rect 9310 21448 9366 21457
rect 9496 21422 9548 21428
rect 9310 21383 9366 21392
rect 9109 21244 9417 21264
rect 9109 21242 9115 21244
rect 9171 21242 9195 21244
rect 9251 21242 9275 21244
rect 9331 21242 9355 21244
rect 9411 21242 9417 21244
rect 9171 21190 9173 21242
rect 9353 21190 9355 21242
rect 9109 21188 9115 21190
rect 9171 21188 9195 21190
rect 9251 21188 9275 21190
rect 9331 21188 9355 21190
rect 9411 21188 9417 21190
rect 9109 21168 9417 21188
rect 9508 21049 9536 21422
rect 9600 21350 9628 33102
rect 9680 33040 9732 33046
rect 9680 32982 9732 32988
rect 9692 27470 9720 32982
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9784 26994 9812 34138
rect 9876 33046 9904 35770
rect 9864 33040 9916 33046
rect 9864 32982 9916 32988
rect 9968 32178 9996 37878
rect 10060 35154 10088 38134
rect 10152 35834 10180 39374
rect 10244 36530 10272 46106
rect 10336 38654 10364 55814
rect 10416 53984 10468 53990
rect 10416 53926 10468 53932
rect 10428 46170 10456 53926
rect 10416 46164 10468 46170
rect 10416 46106 10468 46112
rect 10416 45892 10468 45898
rect 10416 45834 10468 45840
rect 10428 44878 10456 45834
rect 10416 44872 10468 44878
rect 10416 44814 10468 44820
rect 10416 43648 10468 43654
rect 10416 43590 10468 43596
rect 10428 40390 10456 43590
rect 10416 40384 10468 40390
rect 10416 40326 10468 40332
rect 10416 39976 10468 39982
rect 10416 39918 10468 39924
rect 10428 39370 10456 39918
rect 10416 39364 10468 39370
rect 10416 39306 10468 39312
rect 10428 39030 10456 39306
rect 10416 39024 10468 39030
rect 10416 38966 10468 38972
rect 10336 38626 10456 38654
rect 10244 36502 10364 36530
rect 10232 36304 10284 36310
rect 10232 36246 10284 36252
rect 10140 35828 10192 35834
rect 10140 35770 10192 35776
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 10048 35148 10100 35154
rect 10048 35090 10100 35096
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 10060 34241 10088 34886
rect 10152 34649 10180 35430
rect 10138 34640 10194 34649
rect 10138 34575 10194 34584
rect 10140 34536 10192 34542
rect 10140 34478 10192 34484
rect 10046 34232 10102 34241
rect 10046 34167 10102 34176
rect 10048 33856 10100 33862
rect 10048 33798 10100 33804
rect 10060 32881 10088 33798
rect 10152 33454 10180 34478
rect 10140 33448 10192 33454
rect 10140 33390 10192 33396
rect 10152 32978 10180 33390
rect 10140 32972 10192 32978
rect 10140 32914 10192 32920
rect 10046 32872 10102 32881
rect 10046 32807 10102 32816
rect 10048 32564 10100 32570
rect 10048 32506 10100 32512
rect 9876 32150 9996 32178
rect 9876 29646 9904 32150
rect 9956 31748 10008 31754
rect 9956 31690 10008 31696
rect 9968 31482 9996 31690
rect 9956 31476 10008 31482
rect 9956 31418 10008 31424
rect 10060 31362 10088 32506
rect 10140 32496 10192 32502
rect 10140 32438 10192 32444
rect 10152 31754 10180 32438
rect 10140 31748 10192 31754
rect 10140 31690 10192 31696
rect 9968 31334 10088 31362
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 9862 29336 9918 29345
rect 9862 29271 9864 29280
rect 9916 29271 9918 29280
rect 9864 29242 9916 29248
rect 9864 29096 9916 29102
rect 9864 29038 9916 29044
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9876 26058 9904 29038
rect 9968 26382 9996 31334
rect 10048 31272 10100 31278
rect 10048 31214 10100 31220
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 10060 30734 10088 31214
rect 10152 30802 10180 31214
rect 10140 30796 10192 30802
rect 10140 30738 10192 30744
rect 10048 30728 10100 30734
rect 10048 30670 10100 30676
rect 10048 30592 10100 30598
rect 10048 30534 10100 30540
rect 10138 30560 10194 30569
rect 10060 30433 10088 30534
rect 10138 30495 10194 30504
rect 10046 30424 10102 30433
rect 10046 30359 10102 30368
rect 10152 30326 10180 30495
rect 10140 30320 10192 30326
rect 10140 30262 10192 30268
rect 10048 30048 10100 30054
rect 10046 30016 10048 30025
rect 10100 30016 10102 30025
rect 10046 29951 10102 29960
rect 10046 29744 10102 29753
rect 10046 29679 10048 29688
rect 10100 29679 10102 29688
rect 10048 29650 10100 29656
rect 10138 29608 10194 29617
rect 10138 29543 10140 29552
rect 10192 29543 10194 29552
rect 10140 29514 10192 29520
rect 10048 29504 10100 29510
rect 10048 29446 10100 29452
rect 10060 28529 10088 29446
rect 10244 28558 10272 36246
rect 10232 28552 10284 28558
rect 10046 28520 10102 28529
rect 10232 28494 10284 28500
rect 10046 28455 10102 28464
rect 10140 28416 10192 28422
rect 10140 28358 10192 28364
rect 10048 27872 10100 27878
rect 10048 27814 10100 27820
rect 10060 27169 10088 27814
rect 10152 27577 10180 28358
rect 10230 28248 10286 28257
rect 10230 28183 10232 28192
rect 10284 28183 10286 28192
rect 10232 28154 10284 28160
rect 10138 27568 10194 27577
rect 10138 27503 10194 27512
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 10046 27160 10102 27169
rect 10046 27095 10102 27104
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 10060 26217 10088 26726
rect 10152 26625 10180 27270
rect 10138 26616 10194 26625
rect 10138 26551 10194 26560
rect 10046 26208 10102 26217
rect 10046 26143 10102 26152
rect 9876 26030 9996 26058
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9494 21040 9550 21049
rect 9494 20975 9550 20984
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 20505 9352 20878
rect 9588 20528 9640 20534
rect 9310 20496 9366 20505
rect 9588 20470 9640 20476
rect 9310 20431 9366 20440
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9109 20156 9417 20176
rect 9109 20154 9115 20156
rect 9171 20154 9195 20156
rect 9251 20154 9275 20156
rect 9331 20154 9355 20156
rect 9411 20154 9417 20156
rect 9171 20102 9173 20154
rect 9353 20102 9355 20154
rect 9109 20100 9115 20102
rect 9171 20100 9195 20102
rect 9251 20100 9275 20102
rect 9331 20100 9355 20102
rect 9411 20100 9417 20102
rect 9109 20080 9417 20100
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 8956 19502 9076 19530
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 8666 17640 8722 17649
rect 8666 17575 8722 17584
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8680 15162 8708 15302
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8680 7018 8708 13194
rect 8772 10742 8800 17478
rect 8956 16674 8984 19502
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 17882 9076 19314
rect 9324 19258 9352 19926
rect 9508 19802 9536 20402
rect 9600 19922 9628 20470
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9508 19774 9628 19802
rect 9324 19230 9536 19258
rect 9109 19068 9417 19088
rect 9109 19066 9115 19068
rect 9171 19066 9195 19068
rect 9251 19066 9275 19068
rect 9331 19066 9355 19068
rect 9411 19066 9417 19068
rect 9171 19014 9173 19066
rect 9353 19014 9355 19066
rect 9109 19012 9115 19014
rect 9171 19012 9195 19014
rect 9251 19012 9275 19014
rect 9331 19012 9355 19014
rect 9411 19012 9417 19014
rect 9109 18992 9417 19012
rect 9109 17980 9417 18000
rect 9109 17978 9115 17980
rect 9171 17978 9195 17980
rect 9251 17978 9275 17980
rect 9331 17978 9355 17980
rect 9411 17978 9417 17980
rect 9171 17926 9173 17978
rect 9353 17926 9355 17978
rect 9109 17924 9115 17926
rect 9171 17924 9195 17926
rect 9251 17924 9275 17926
rect 9331 17924 9355 17926
rect 9411 17924 9417 17926
rect 9109 17904 9417 17924
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9140 17338 9168 17546
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9109 16892 9417 16912
rect 9109 16890 9115 16892
rect 9171 16890 9195 16892
rect 9251 16890 9275 16892
rect 9331 16890 9355 16892
rect 9411 16890 9417 16892
rect 9171 16838 9173 16890
rect 9353 16838 9355 16890
rect 9109 16836 9115 16838
rect 9171 16836 9195 16838
rect 9251 16836 9275 16838
rect 9331 16836 9355 16838
rect 9411 16836 9417 16838
rect 9109 16816 9417 16836
rect 8956 16646 9260 16674
rect 8956 15366 8984 16646
rect 9232 16590 9260 16646
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9109 15804 9417 15824
rect 9109 15802 9115 15804
rect 9171 15802 9195 15804
rect 9251 15802 9275 15804
rect 9331 15802 9355 15804
rect 9411 15802 9417 15804
rect 9171 15750 9173 15802
rect 9353 15750 9355 15802
rect 9109 15748 9115 15750
rect 9171 15748 9195 15750
rect 9251 15748 9275 15750
rect 9331 15748 9355 15750
rect 9411 15748 9417 15750
rect 9109 15728 9417 15748
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 15366 9444 15438
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 8850 15192 8906 15201
rect 8850 15127 8852 15136
rect 8904 15127 8906 15136
rect 8852 15098 8904 15104
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8956 14618 8984 14758
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9048 14498 9076 14962
rect 9109 14716 9417 14736
rect 9109 14714 9115 14716
rect 9171 14714 9195 14716
rect 9251 14714 9275 14716
rect 9331 14714 9355 14716
rect 9411 14714 9417 14716
rect 9171 14662 9173 14714
rect 9353 14662 9355 14714
rect 9109 14660 9115 14662
rect 9171 14660 9195 14662
rect 9251 14660 9275 14662
rect 9331 14660 9355 14662
rect 9411 14660 9417 14662
rect 9109 14640 9417 14660
rect 8944 14476 8996 14482
rect 9048 14470 9168 14498
rect 8944 14418 8996 14424
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 12918 8892 14214
rect 8956 12986 8984 14418
rect 9140 14414 9168 14470
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8864 12442 8892 12718
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8956 11354 8984 12786
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8772 10266 8800 10542
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8864 9654 8892 10610
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8496 6990 8708 7018
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8496 3074 8524 6990
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8588 3126 8616 5510
rect 8680 3602 8708 6598
rect 8772 5166 8800 7142
rect 8864 6866 8892 9386
rect 8956 8634 8984 10542
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8956 7313 8984 7346
rect 8942 7304 8998 7313
rect 8942 7239 8998 7248
rect 9048 7154 9076 13874
rect 9140 13870 9168 14350
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9416 14006 9444 14214
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9109 13628 9417 13648
rect 9109 13626 9115 13628
rect 9171 13626 9195 13628
rect 9251 13626 9275 13628
rect 9331 13626 9355 13628
rect 9411 13626 9417 13628
rect 9171 13574 9173 13626
rect 9353 13574 9355 13626
rect 9109 13572 9115 13574
rect 9171 13572 9195 13574
rect 9251 13572 9275 13574
rect 9331 13572 9355 13574
rect 9411 13572 9417 13574
rect 9109 13552 9417 13572
rect 9508 13274 9536 19230
rect 9600 19145 9628 19774
rect 9692 19446 9720 23666
rect 9784 22794 9812 25094
rect 9876 24721 9904 25842
rect 9968 25362 9996 26030
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 9968 25242 9996 25298
rect 9968 25214 10180 25242
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 9862 24712 9918 24721
rect 9862 24647 9918 24656
rect 9968 23361 9996 24754
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 9954 23352 10010 23361
rect 9954 23287 10010 23296
rect 9784 22766 9904 22794
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9784 21894 9812 22578
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9876 19530 9904 22766
rect 10060 22409 10088 24142
rect 10152 23662 10180 25214
rect 10336 24818 10364 36502
rect 10428 33538 10456 38626
rect 10520 36689 10548 61066
rect 10612 36825 10640 65418
rect 11428 62824 11480 62830
rect 11428 62766 11480 62772
rect 11244 62416 11296 62422
rect 11244 62358 11296 62364
rect 10968 60988 11020 60994
rect 10968 60930 11020 60936
rect 10980 60654 11008 60930
rect 11256 60790 11284 62358
rect 11336 61056 11388 61062
rect 11336 60998 11388 61004
rect 11244 60784 11296 60790
rect 11244 60726 11296 60732
rect 10968 60648 11020 60654
rect 10968 60590 11020 60596
rect 10784 59492 10836 59498
rect 10784 59434 10836 59440
rect 10692 56160 10744 56166
rect 10692 56102 10744 56108
rect 10704 52465 10732 56102
rect 10690 52456 10746 52465
rect 10690 52391 10746 52400
rect 10692 52352 10744 52358
rect 10692 52294 10744 52300
rect 10704 50998 10732 52294
rect 10796 51270 10824 59434
rect 11244 57792 11296 57798
rect 11244 57734 11296 57740
rect 11256 57338 11284 57734
rect 11348 57526 11376 60998
rect 11440 60858 11468 62766
rect 11428 60852 11480 60858
rect 11428 60794 11480 60800
rect 11520 60308 11572 60314
rect 11520 60250 11572 60256
rect 11336 57520 11388 57526
rect 11336 57462 11388 57468
rect 11256 57310 11376 57338
rect 11152 57248 11204 57254
rect 11152 57190 11204 57196
rect 10968 56092 11020 56098
rect 10968 56034 11020 56040
rect 10876 55208 10928 55214
rect 10876 55150 10928 55156
rect 10888 51610 10916 55150
rect 10980 53281 11008 56034
rect 10966 53272 11022 53281
rect 10966 53207 11022 53216
rect 10968 53168 11020 53174
rect 10968 53110 11020 53116
rect 10876 51604 10928 51610
rect 10876 51546 10928 51552
rect 10980 51513 11008 53110
rect 10966 51504 11022 51513
rect 10876 51468 10928 51474
rect 10966 51439 11022 51448
rect 10876 51410 10928 51416
rect 10784 51264 10836 51270
rect 10784 51206 10836 51212
rect 10782 51096 10838 51105
rect 10782 51031 10838 51040
rect 10692 50992 10744 50998
rect 10692 50934 10744 50940
rect 10796 50844 10824 51031
rect 10704 50816 10824 50844
rect 10704 43314 10732 50816
rect 10784 50720 10836 50726
rect 10784 50662 10836 50668
rect 10796 50164 10824 50662
rect 10888 50266 10916 51410
rect 10968 51400 11020 51406
rect 10966 51368 10968 51377
rect 11060 51400 11112 51406
rect 11020 51368 11022 51377
rect 11060 51342 11112 51348
rect 10966 51303 11022 51312
rect 10968 51196 11020 51202
rect 10968 51138 11020 51144
rect 10980 51066 11008 51138
rect 10968 51060 11020 51066
rect 10968 51002 11020 51008
rect 11072 50708 11100 51342
rect 11164 50862 11192 57190
rect 11244 52896 11296 52902
rect 11244 52838 11296 52844
rect 11152 50856 11204 50862
rect 11152 50798 11204 50804
rect 10980 50680 11100 50708
rect 10980 50368 11008 50680
rect 10980 50340 11192 50368
rect 10888 50238 11100 50266
rect 10796 50136 10916 50164
rect 10784 48680 10836 48686
rect 10784 48622 10836 48628
rect 10692 43308 10744 43314
rect 10692 43250 10744 43256
rect 10692 42900 10744 42906
rect 10692 42842 10744 42848
rect 10704 41721 10732 42842
rect 10690 41712 10746 41721
rect 10690 41647 10746 41656
rect 10692 41608 10744 41614
rect 10692 41550 10744 41556
rect 10704 39930 10732 41550
rect 10796 41546 10824 48622
rect 10888 47546 10916 50136
rect 10968 49360 11020 49366
rect 10966 49328 10968 49337
rect 11020 49328 11022 49337
rect 10966 49263 11022 49272
rect 10888 47518 11008 47546
rect 10876 47252 10928 47258
rect 10876 47194 10928 47200
rect 10784 41540 10836 41546
rect 10784 41482 10836 41488
rect 10782 41440 10838 41449
rect 10782 41375 10838 41384
rect 10796 40458 10824 41375
rect 10888 40934 10916 47194
rect 10980 45490 11008 47518
rect 10968 45484 11020 45490
rect 10968 45426 11020 45432
rect 11072 43246 11100 50238
rect 11164 49094 11192 50340
rect 11256 49842 11284 52838
rect 11348 51474 11376 57310
rect 11532 53242 11560 60250
rect 11716 57934 11744 66098
rect 11796 60852 11848 60858
rect 11796 60794 11848 60800
rect 11704 57928 11756 57934
rect 11704 57870 11756 57876
rect 11704 56976 11756 56982
rect 11704 56918 11756 56924
rect 11716 56273 11744 56918
rect 11808 56846 11836 60794
rect 11888 58404 11940 58410
rect 11888 58346 11940 58352
rect 11796 56840 11848 56846
rect 11796 56782 11848 56788
rect 11702 56264 11758 56273
rect 11702 56199 11758 56208
rect 11796 55888 11848 55894
rect 11796 55830 11848 55836
rect 11808 54369 11836 55830
rect 11794 54360 11850 54369
rect 11794 54295 11850 54304
rect 11520 53236 11572 53242
rect 11520 53178 11572 53184
rect 11520 53100 11572 53106
rect 11520 53042 11572 53048
rect 11428 52692 11480 52698
rect 11428 52634 11480 52640
rect 11336 51468 11388 51474
rect 11336 51410 11388 51416
rect 11440 51218 11468 52634
rect 11532 51388 11560 53042
rect 11900 53038 11928 58346
rect 11888 53032 11940 53038
rect 11888 52974 11940 52980
rect 11796 51400 11848 51406
rect 11532 51360 11652 51388
rect 11440 51190 11560 51218
rect 11336 51128 11388 51134
rect 11336 51070 11388 51076
rect 11348 50658 11376 51070
rect 11428 50720 11480 50726
rect 11428 50662 11480 50668
rect 11336 50652 11388 50658
rect 11336 50594 11388 50600
rect 11334 50552 11390 50561
rect 11334 50487 11390 50496
rect 11244 49836 11296 49842
rect 11244 49778 11296 49784
rect 11152 49088 11204 49094
rect 11152 49030 11204 49036
rect 11244 48136 11296 48142
rect 11244 48078 11296 48084
rect 11256 46578 11284 48078
rect 11244 46572 11296 46578
rect 11244 46514 11296 46520
rect 11256 45370 11284 46514
rect 11164 45342 11284 45370
rect 11164 43994 11192 45342
rect 11244 45280 11296 45286
rect 11244 45222 11296 45228
rect 11152 43988 11204 43994
rect 11152 43930 11204 43936
rect 10968 43240 11020 43246
rect 10968 43182 11020 43188
rect 11060 43240 11112 43246
rect 11060 43182 11112 43188
rect 10980 41138 11008 43182
rect 11060 43104 11112 43110
rect 11060 43046 11112 43052
rect 11072 41342 11100 43046
rect 11152 42764 11204 42770
rect 11152 42706 11204 42712
rect 11164 42294 11192 42706
rect 11152 42288 11204 42294
rect 11152 42230 11204 42236
rect 11256 42106 11284 45222
rect 11348 43722 11376 50487
rect 11336 43716 11388 43722
rect 11336 43658 11388 43664
rect 11440 43489 11468 50662
rect 11426 43480 11482 43489
rect 11426 43415 11482 43424
rect 11336 43240 11388 43246
rect 11336 43182 11388 43188
rect 11164 42078 11284 42106
rect 11164 41614 11192 42078
rect 11348 41886 11376 43182
rect 11532 42537 11560 51190
rect 11624 48142 11652 51360
rect 11796 51342 11848 51348
rect 11704 50992 11756 50998
rect 11704 50934 11756 50940
rect 11612 48136 11664 48142
rect 11612 48078 11664 48084
rect 11612 48000 11664 48006
rect 11612 47942 11664 47948
rect 11624 43790 11652 47942
rect 11716 45626 11744 50934
rect 11808 50386 11836 51342
rect 11888 50448 11940 50454
rect 11888 50390 11940 50396
rect 11796 50380 11848 50386
rect 11796 50322 11848 50328
rect 11796 49768 11848 49774
rect 11796 49710 11848 49716
rect 11704 45620 11756 45626
rect 11704 45562 11756 45568
rect 11704 45484 11756 45490
rect 11704 45426 11756 45432
rect 11612 43784 11664 43790
rect 11612 43726 11664 43732
rect 11612 43648 11664 43654
rect 11612 43590 11664 43596
rect 11518 42528 11574 42537
rect 11518 42463 11574 42472
rect 11624 42242 11652 43590
rect 11716 42770 11744 45426
rect 11704 42764 11756 42770
rect 11704 42706 11756 42712
rect 11704 42560 11756 42566
rect 11704 42502 11756 42508
rect 11532 42214 11652 42242
rect 11336 41880 11388 41886
rect 11336 41822 11388 41828
rect 11532 41800 11560 42214
rect 11612 41880 11664 41886
rect 11612 41822 11664 41828
rect 11440 41772 11560 41800
rect 11336 41744 11388 41750
rect 11336 41686 11388 41692
rect 11152 41608 11204 41614
rect 11152 41550 11204 41556
rect 11244 41472 11296 41478
rect 11244 41414 11296 41420
rect 11060 41336 11112 41342
rect 11060 41278 11112 41284
rect 11152 41336 11204 41342
rect 11152 41278 11204 41284
rect 11060 41200 11112 41206
rect 11060 41142 11112 41148
rect 10968 41132 11020 41138
rect 10968 41074 11020 41080
rect 10968 40996 11020 41002
rect 10968 40938 11020 40944
rect 10876 40928 10928 40934
rect 10876 40870 10928 40876
rect 10876 40724 10928 40730
rect 10876 40666 10928 40672
rect 10784 40452 10836 40458
rect 10784 40394 10836 40400
rect 10782 40216 10838 40225
rect 10782 40151 10838 40160
rect 10796 40118 10824 40151
rect 10784 40112 10836 40118
rect 10784 40054 10836 40060
rect 10704 39902 10824 39930
rect 10692 39840 10744 39846
rect 10692 39782 10744 39788
rect 10598 36816 10654 36825
rect 10598 36751 10654 36760
rect 10506 36680 10562 36689
rect 10506 36615 10562 36624
rect 10704 33538 10732 39782
rect 10796 33658 10824 39902
rect 10888 33998 10916 40666
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10428 33510 10548 33538
rect 10704 33510 10916 33538
rect 10414 33416 10470 33425
rect 10414 33351 10470 33360
rect 10428 31278 10456 33351
rect 10520 32065 10548 33510
rect 10692 33312 10744 33318
rect 10692 33254 10744 33260
rect 10598 33144 10654 33153
rect 10598 33079 10600 33088
rect 10652 33079 10654 33088
rect 10600 33050 10652 33056
rect 10600 32972 10652 32978
rect 10600 32914 10652 32920
rect 10506 32056 10562 32065
rect 10506 31991 10562 32000
rect 10612 31906 10640 32914
rect 10520 31878 10640 31906
rect 10416 31272 10468 31278
rect 10416 31214 10468 31220
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10428 30977 10456 31078
rect 10414 30968 10470 30977
rect 10414 30903 10470 30912
rect 10414 30832 10470 30841
rect 10414 30767 10416 30776
rect 10468 30767 10470 30776
rect 10416 30738 10468 30744
rect 10416 30660 10468 30666
rect 10416 30602 10468 30608
rect 10428 29102 10456 30602
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10152 23202 10180 23598
rect 10152 23186 10272 23202
rect 10140 23180 10272 23186
rect 10192 23174 10272 23180
rect 10140 23122 10192 23128
rect 10140 23044 10192 23050
rect 10140 22986 10192 22992
rect 10046 22400 10102 22409
rect 10046 22335 10102 22344
rect 9956 21412 10008 21418
rect 9956 21354 10008 21360
rect 9968 19922 9996 21354
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9784 19502 9904 19530
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9586 19136 9642 19145
rect 9586 19071 9642 19080
rect 9784 18970 9812 19502
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9600 17338 9628 18362
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9692 16182 9720 18566
rect 9876 17746 9904 19314
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9968 17626 9996 19382
rect 9784 17598 9996 17626
rect 9784 17542 9812 17598
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 13462 9628 15982
rect 9784 15502 9812 17478
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9784 15162 9812 15302
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9876 14482 9904 17478
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9968 14074 9996 16730
rect 10060 15978 10088 19654
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10152 15638 10180 22986
rect 10244 22574 10272 23174
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10336 22098 10364 22646
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10428 22030 10456 25366
rect 10520 24342 10548 31878
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10612 31362 10640 31758
rect 10704 31482 10732 33254
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10692 31476 10744 31482
rect 10692 31418 10744 31424
rect 10612 31334 10732 31362
rect 10598 31240 10654 31249
rect 10704 31210 10732 31334
rect 10598 31175 10654 31184
rect 10692 31204 10744 31210
rect 10612 30258 10640 31175
rect 10692 31146 10744 31152
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10508 24336 10560 24342
rect 10508 24278 10560 24284
rect 10612 22386 10640 26318
rect 10520 22358 10640 22386
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 10244 18970 10272 21558
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10336 19446 10364 19858
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10336 18834 10364 19382
rect 10520 19378 10548 22358
rect 10704 22094 10732 31146
rect 10796 22506 10824 31962
rect 10888 31906 10916 33510
rect 10980 32008 11008 40938
rect 11072 32502 11100 41142
rect 11060 32496 11112 32502
rect 11060 32438 11112 32444
rect 11164 32298 11192 41278
rect 11152 32292 11204 32298
rect 11152 32234 11204 32240
rect 11256 32026 11284 41414
rect 11348 37126 11376 41686
rect 11336 37120 11388 37126
rect 11336 37062 11388 37068
rect 11336 36984 11388 36990
rect 11336 36926 11388 36932
rect 11348 33046 11376 36926
rect 11336 33040 11388 33046
rect 11336 32982 11388 32988
rect 11336 32700 11388 32706
rect 11336 32642 11388 32648
rect 11348 32026 11376 32642
rect 11440 32434 11468 41772
rect 11624 41290 11652 41822
rect 11532 41262 11652 41290
rect 11532 41154 11560 41262
rect 11532 41126 11652 41154
rect 11520 41064 11572 41070
rect 11520 41006 11572 41012
rect 11532 32978 11560 41006
rect 11624 40662 11652 41126
rect 11612 40656 11664 40662
rect 11612 40598 11664 40604
rect 11610 38720 11666 38729
rect 11610 38655 11666 38664
rect 11624 36990 11652 38655
rect 11612 36984 11664 36990
rect 11612 36926 11664 36932
rect 11612 36848 11664 36854
rect 11610 36816 11612 36825
rect 11664 36816 11666 36825
rect 11610 36751 11666 36760
rect 11612 36576 11664 36582
rect 11612 36518 11664 36524
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11428 32428 11480 32434
rect 11428 32370 11480 32376
rect 11624 32280 11652 36518
rect 11716 32774 11744 42502
rect 11808 41070 11836 49710
rect 11900 42022 11928 50390
rect 11888 42016 11940 42022
rect 11888 41958 11940 41964
rect 11888 41540 11940 41546
rect 11888 41482 11940 41488
rect 11796 41064 11848 41070
rect 11796 41006 11848 41012
rect 11796 40384 11848 40390
rect 11796 40326 11848 40332
rect 11704 32768 11756 32774
rect 11704 32710 11756 32716
rect 11808 32586 11836 40326
rect 11900 39681 11928 41482
rect 11886 39672 11942 39681
rect 11886 39607 11942 39616
rect 11888 39568 11940 39574
rect 11888 39510 11940 39516
rect 11900 32706 11928 39510
rect 11888 32700 11940 32706
rect 11888 32642 11940 32648
rect 11440 32252 11652 32280
rect 11716 32558 11836 32586
rect 11886 32600 11942 32609
rect 11244 32020 11296 32026
rect 10980 31980 11192 32008
rect 10888 31878 11100 31906
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 10888 31657 10916 31758
rect 10874 31648 10930 31657
rect 10874 31583 10930 31592
rect 10968 31272 11020 31278
rect 10968 31214 11020 31220
rect 10980 25430 11008 31214
rect 10968 25424 11020 25430
rect 10968 25366 11020 25372
rect 10968 25288 11020 25294
rect 10966 25256 10968 25265
rect 11020 25256 11022 25265
rect 10966 25191 11022 25200
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 11072 22386 11100 31878
rect 11164 31498 11192 31980
rect 11244 31962 11296 31968
rect 11336 32020 11388 32026
rect 11336 31962 11388 31968
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 11164 31470 11284 31498
rect 11256 28218 11284 31470
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 10612 22066 10732 22094
rect 10796 22358 11100 22386
rect 10612 20602 10640 22066
rect 10796 21554 10824 22358
rect 11060 22296 11112 22302
rect 10966 22264 11022 22273
rect 11060 22238 11112 22244
rect 10966 22199 11022 22208
rect 10980 22166 11008 22199
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 11072 21758 11100 22238
rect 11060 21752 11112 21758
rect 11060 21694 11112 21700
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 11164 20874 11192 22714
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11256 21962 11284 22374
rect 11348 22302 11376 31758
rect 11440 31618 11468 32252
rect 11612 31952 11664 31958
rect 11612 31894 11664 31900
rect 11428 31612 11480 31618
rect 11428 31554 11480 31560
rect 11520 31544 11572 31550
rect 11520 31486 11572 31492
rect 11532 23866 11560 31486
rect 11624 31362 11652 31894
rect 11716 31618 11744 32558
rect 11886 32535 11942 32544
rect 11796 32088 11848 32094
rect 11796 32030 11848 32036
rect 11704 31612 11756 31618
rect 11704 31554 11756 31560
rect 11624 31334 11744 31362
rect 11612 31272 11664 31278
rect 11612 31214 11664 31220
rect 11624 25974 11652 31214
rect 11612 25968 11664 25974
rect 11612 25910 11664 25916
rect 11716 24138 11744 31334
rect 11808 24682 11836 32030
rect 11900 31822 11928 32535
rect 11888 31816 11940 31822
rect 11888 31758 11940 31764
rect 11886 29744 11942 29753
rect 11886 29679 11888 29688
rect 11940 29679 11942 29688
rect 11888 29650 11940 29656
rect 11888 28212 11940 28218
rect 11888 28154 11940 28160
rect 11796 24676 11848 24682
rect 11796 24618 11848 24624
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11336 22296 11388 22302
rect 11336 22238 11388 22244
rect 11704 22296 11756 22302
rect 11704 22238 11756 22244
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10336 17746 10364 18770
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 16250 10272 17138
rect 10336 17134 10364 17682
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10336 16658 10364 17070
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10336 16046 10364 16594
rect 11060 16312 11112 16318
rect 11058 16280 11060 16289
rect 11112 16280 11114 16289
rect 11058 16215 11114 16224
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10336 15570 10364 15982
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10336 14958 10364 15506
rect 11532 15162 11560 22034
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11624 16590 11652 21830
rect 11716 21758 11744 22238
rect 11808 21962 11836 24142
rect 11796 21956 11848 21962
rect 11796 21898 11848 21904
rect 11704 21752 11756 21758
rect 11704 21694 11756 21700
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11900 16182 11928 28154
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10336 14482 10364 14894
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9416 13246 9536 13274
rect 9416 12850 9444 13246
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9109 12540 9417 12560
rect 9109 12538 9115 12540
rect 9171 12538 9195 12540
rect 9251 12538 9275 12540
rect 9331 12538 9355 12540
rect 9411 12538 9417 12540
rect 9171 12486 9173 12538
rect 9353 12486 9355 12538
rect 9109 12484 9115 12486
rect 9171 12484 9195 12486
rect 9251 12484 9275 12486
rect 9331 12484 9355 12486
rect 9411 12484 9417 12486
rect 9109 12464 9417 12484
rect 9508 12170 9536 13126
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11830 9444 12038
rect 9404 11824 9456 11830
rect 9404 11766 9456 11772
rect 9109 11452 9417 11472
rect 9109 11450 9115 11452
rect 9171 11450 9195 11452
rect 9251 11450 9275 11452
rect 9331 11450 9355 11452
rect 9411 11450 9417 11452
rect 9171 11398 9173 11450
rect 9353 11398 9355 11450
rect 9109 11396 9115 11398
rect 9171 11396 9195 11398
rect 9251 11396 9275 11398
rect 9331 11396 9355 11398
rect 9411 11396 9417 11398
rect 9109 11376 9417 11396
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9416 10538 9444 11154
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9109 10364 9417 10384
rect 9109 10362 9115 10364
rect 9171 10362 9195 10364
rect 9251 10362 9275 10364
rect 9331 10362 9355 10364
rect 9411 10362 9417 10364
rect 9171 10310 9173 10362
rect 9353 10310 9355 10362
rect 9109 10308 9115 10310
rect 9171 10308 9195 10310
rect 9251 10308 9275 10310
rect 9331 10308 9355 10310
rect 9411 10308 9417 10310
rect 9109 10288 9417 10308
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9232 9450 9260 10095
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9109 9276 9417 9296
rect 9109 9274 9115 9276
rect 9171 9274 9195 9276
rect 9251 9274 9275 9276
rect 9331 9274 9355 9276
rect 9411 9274 9417 9276
rect 9171 9222 9173 9274
rect 9353 9222 9355 9274
rect 9109 9220 9115 9222
rect 9171 9220 9195 9222
rect 9251 9220 9275 9222
rect 9331 9220 9355 9222
rect 9411 9220 9417 9222
rect 9109 9200 9417 9220
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9140 8673 9168 8910
rect 9126 8664 9182 8673
rect 9126 8599 9182 8608
rect 9109 8188 9417 8208
rect 9109 8186 9115 8188
rect 9171 8186 9195 8188
rect 9251 8186 9275 8188
rect 9331 8186 9355 8188
rect 9411 8186 9417 8188
rect 9171 8134 9173 8186
rect 9353 8134 9355 8186
rect 9109 8132 9115 8134
rect 9171 8132 9195 8134
rect 9251 8132 9275 8134
rect 9331 8132 9355 8134
rect 9411 8132 9417 8134
rect 9109 8112 9417 8132
rect 8956 7126 9076 7154
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8864 6458 8892 6802
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8864 5778 8892 6054
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8956 5658 8984 7126
rect 9109 7100 9417 7120
rect 9109 7098 9115 7100
rect 9171 7098 9195 7100
rect 9251 7098 9275 7100
rect 9331 7098 9355 7100
rect 9411 7098 9417 7100
rect 9171 7046 9173 7098
rect 9353 7046 9355 7098
rect 9109 7044 9115 7046
rect 9171 7044 9195 7046
rect 9251 7044 9275 7046
rect 9331 7044 9355 7046
rect 9411 7044 9417 7046
rect 9109 7024 9417 7044
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8864 5630 8984 5658
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8772 4622 8800 4966
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8864 3602 8892 5630
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 4457 8984 5170
rect 8942 4448 8998 4457
rect 8942 4383 8998 4392
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8404 3046 8524 3074
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8404 2774 8432 3046
rect 8956 2990 8984 4014
rect 9048 4010 9076 6666
rect 9109 6012 9417 6032
rect 9109 6010 9115 6012
rect 9171 6010 9195 6012
rect 9251 6010 9275 6012
rect 9331 6010 9355 6012
rect 9411 6010 9417 6012
rect 9171 5958 9173 6010
rect 9353 5958 9355 6010
rect 9109 5956 9115 5958
rect 9171 5956 9195 5958
rect 9251 5956 9275 5958
rect 9331 5956 9355 5958
rect 9411 5956 9417 5958
rect 9109 5936 9417 5956
rect 9109 4924 9417 4944
rect 9109 4922 9115 4924
rect 9171 4922 9195 4924
rect 9251 4922 9275 4924
rect 9331 4922 9355 4924
rect 9411 4922 9417 4924
rect 9171 4870 9173 4922
rect 9353 4870 9355 4922
rect 9109 4868 9115 4870
rect 9171 4868 9195 4870
rect 9251 4868 9275 4870
rect 9331 4868 9355 4870
rect 9411 4868 9417 4870
rect 9109 4848 9417 4868
rect 9508 4706 9536 10678
rect 9600 8566 9628 12922
rect 9692 12238 9720 13874
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9968 13394 9996 13806
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 10198 9720 12038
rect 9784 11286 9812 13126
rect 9968 12306 9996 13330
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9876 10810 9904 11290
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9968 10606 9996 12242
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9784 10062 9812 10406
rect 9968 10130 9996 10542
rect 10428 10169 10456 10610
rect 10414 10160 10470 10169
rect 9956 10124 10008 10130
rect 10414 10095 10470 10104
rect 9956 10066 10008 10072
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9770 9616 9826 9625
rect 9770 9551 9772 9560
rect 9824 9551 9826 9560
rect 9772 9522 9824 9528
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9876 8265 9904 8910
rect 9862 8256 9918 8265
rect 9862 8191 9918 8200
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9692 5370 9720 7346
rect 9784 6361 9812 7754
rect 9968 7342 9996 10066
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10244 7721 10272 8434
rect 10230 7712 10286 7721
rect 10230 7647 10286 7656
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9968 6866 9996 7278
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9770 6352 9826 6361
rect 9770 6287 9826 6296
rect 9968 5778 9996 6802
rect 10968 6792 11020 6798
rect 10966 6760 10968 6769
rect 11020 6760 11022 6769
rect 10966 6695 11022 6704
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 4826 9628 5102
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9232 4678 9536 4706
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9140 4049 9168 4082
rect 9232 4078 9260 4678
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9416 4214 9444 4422
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9496 4140 9548 4146
rect 9548 4100 9628 4128
rect 9496 4082 9548 4088
rect 9220 4072 9272 4078
rect 9126 4040 9182 4049
rect 9036 4004 9088 4010
rect 9220 4014 9272 4020
rect 9126 3975 9182 3984
rect 9036 3946 9088 3952
rect 9109 3836 9417 3856
rect 9109 3834 9115 3836
rect 9171 3834 9195 3836
rect 9251 3834 9275 3836
rect 9331 3834 9355 3836
rect 9411 3834 9417 3836
rect 9171 3782 9173 3834
rect 9353 3782 9355 3834
rect 9109 3780 9115 3782
rect 9171 3780 9195 3782
rect 9251 3780 9275 3782
rect 9331 3780 9355 3782
rect 9411 3780 9417 3782
rect 9109 3760 9417 3780
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8404 2746 8524 2774
rect 8496 2514 8524 2746
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8588 2446 8616 2858
rect 9109 2748 9417 2768
rect 9109 2746 9115 2748
rect 9171 2746 9195 2748
rect 9251 2746 9275 2748
rect 9331 2746 9355 2748
rect 9411 2746 9417 2748
rect 9171 2694 9173 2746
rect 9353 2694 9355 2746
rect 9109 2692 9115 2694
rect 9171 2692 9195 2694
rect 9251 2692 9275 2694
rect 9331 2692 9355 2694
rect 9411 2692 9417 2694
rect 9109 2672 9417 2692
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9324 1057 9352 2382
rect 9508 2009 9536 3470
rect 9600 2553 9628 4100
rect 9784 3738 9812 5170
rect 9968 5166 9996 5714
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 4690 9996 5102
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9968 3194 9996 4626
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9586 2544 9642 2553
rect 9586 2479 9642 2488
rect 9494 2000 9550 2009
rect 9494 1935 9550 1944
rect 9310 1048 9366 1057
rect 9310 983 9366 992
rect 8206 640 8262 649
rect 8206 575 8262 584
rect 8114 232 8170 241
rect 8114 167 8170 176
<< via2 >>
rect 3238 79600 3294 79656
rect 7562 79600 7618 79656
rect 1398 78920 1454 78976
rect 2962 78240 3018 78296
rect 2588 77818 2644 77820
rect 2668 77818 2724 77820
rect 2748 77818 2804 77820
rect 2828 77818 2884 77820
rect 2588 77766 2634 77818
rect 2634 77766 2644 77818
rect 2668 77766 2698 77818
rect 2698 77766 2710 77818
rect 2710 77766 2724 77818
rect 2748 77766 2762 77818
rect 2762 77766 2774 77818
rect 2774 77766 2804 77818
rect 2828 77766 2838 77818
rect 2838 77766 2884 77818
rect 2588 77764 2644 77766
rect 2668 77764 2724 77766
rect 2748 77764 2804 77766
rect 2828 77764 2884 77766
rect 2870 77560 2926 77616
rect 1582 76880 1638 76936
rect 2588 76730 2644 76732
rect 2668 76730 2724 76732
rect 2748 76730 2804 76732
rect 2828 76730 2884 76732
rect 2588 76678 2634 76730
rect 2634 76678 2644 76730
rect 2668 76678 2698 76730
rect 2698 76678 2710 76730
rect 2710 76678 2724 76730
rect 2748 76678 2762 76730
rect 2762 76678 2774 76730
rect 2774 76678 2804 76730
rect 2828 76678 2838 76730
rect 2838 76678 2884 76730
rect 2588 76676 2644 76678
rect 2668 76676 2724 76678
rect 2748 76676 2804 76678
rect 2828 76676 2884 76678
rect 1582 76200 1638 76256
rect 1398 75520 1454 75576
rect 1582 73616 1638 73672
rect 1582 71576 1638 71632
rect 1398 70932 1400 70952
rect 1400 70932 1452 70952
rect 1452 70932 1454 70952
rect 1398 70896 1454 70932
rect 1490 70488 1546 70544
rect 1030 63008 1086 63064
rect 1582 68312 1638 68368
rect 1398 67668 1400 67688
rect 1400 67668 1452 67688
rect 1452 67668 1454 67688
rect 1398 67632 1454 67668
rect 1490 66952 1546 67008
rect 1398 63688 1454 63744
rect 1398 62328 1454 62384
rect 1398 61104 1454 61160
rect 1582 65728 1638 65784
rect 1858 74976 1914 75032
rect 2588 75642 2644 75644
rect 2668 75642 2724 75644
rect 2748 75642 2804 75644
rect 2828 75642 2884 75644
rect 2588 75590 2634 75642
rect 2634 75590 2644 75642
rect 2668 75590 2698 75642
rect 2698 75590 2710 75642
rect 2710 75590 2724 75642
rect 2748 75590 2762 75642
rect 2762 75590 2774 75642
rect 2774 75590 2804 75642
rect 2828 75590 2838 75642
rect 2838 75590 2884 75642
rect 2588 75588 2644 75590
rect 2668 75588 2724 75590
rect 2748 75588 2804 75590
rect 2828 75588 2884 75590
rect 2226 74296 2282 74352
rect 2588 74554 2644 74556
rect 2668 74554 2724 74556
rect 2748 74554 2804 74556
rect 2828 74554 2884 74556
rect 2588 74502 2634 74554
rect 2634 74502 2644 74554
rect 2668 74502 2698 74554
rect 2698 74502 2710 74554
rect 2710 74502 2724 74554
rect 2748 74502 2762 74554
rect 2762 74502 2774 74554
rect 2774 74502 2804 74554
rect 2828 74502 2838 74554
rect 2838 74502 2884 74554
rect 2588 74500 2644 74502
rect 2668 74500 2724 74502
rect 2748 74500 2804 74502
rect 2828 74500 2884 74502
rect 2226 72256 2282 72312
rect 1858 64368 1914 64424
rect 1582 59472 1638 59528
rect 1582 58404 1638 58440
rect 1582 58384 1584 58404
rect 1584 58384 1636 58404
rect 1636 58384 1638 58404
rect 1582 57740 1584 57760
rect 1584 57740 1636 57760
rect 1636 57740 1638 57760
rect 1582 57704 1638 57740
rect 1582 57024 1638 57080
rect 1582 56480 1638 56536
rect 1582 55800 1638 55856
rect 1582 55120 1638 55176
rect 1582 54440 1638 54496
rect 1582 53780 1638 53816
rect 1582 53760 1584 53780
rect 1584 53760 1636 53780
rect 1636 53760 1638 53780
rect 1398 51176 1454 51232
rect 1582 53080 1638 53136
rect 1398 45192 1454 45248
rect 1398 42644 1400 42664
rect 1400 42644 1452 42664
rect 1452 42644 1454 42664
rect 1398 42608 1454 42644
rect 1398 41928 1454 41984
rect 1398 41248 1454 41304
rect 1398 39924 1400 39944
rect 1400 39924 1452 39944
rect 1452 39924 1454 39944
rect 1398 39888 1454 39924
rect 1858 61648 1914 61704
rect 1858 59744 1914 59800
rect 1858 59064 1914 59120
rect 2226 65048 2282 65104
rect 1858 51856 1914 51912
rect 1858 50496 1914 50552
rect 1858 49816 1914 49872
rect 1858 49172 1860 49192
rect 1860 49172 1912 49192
rect 1912 49172 1914 49192
rect 1858 49136 1914 49172
rect 1858 48456 1914 48512
rect 1858 47776 1914 47832
rect 1858 47232 1914 47288
rect 1858 46552 1914 46608
rect 1858 45908 1860 45928
rect 1860 45908 1912 45928
rect 1912 45908 1914 45928
rect 1858 45872 1914 45908
rect 1398 38528 1454 38584
rect 1398 37848 1454 37904
rect 1306 37304 1362 37360
rect 1398 36660 1400 36680
rect 1400 36660 1452 36680
rect 1452 36660 1454 36680
rect 1398 36624 1454 36660
rect 1398 33940 1400 33960
rect 1400 33940 1452 33960
rect 1452 33940 1454 33960
rect 1398 33904 1454 33940
rect 1398 33224 1454 33280
rect 1582 35944 1638 36000
rect 1582 35264 1638 35320
rect 1582 34584 1638 34640
rect 1582 32680 1638 32736
rect 1582 32000 1638 32056
rect 1582 31320 1638 31376
rect 1582 30640 1638 30696
rect 1582 29996 1584 30016
rect 1584 29996 1636 30016
rect 1636 29996 1638 30016
rect 1582 29960 1638 29996
rect 1582 29280 1638 29336
rect 1582 28600 1638 28656
rect 1582 28056 1638 28112
rect 1582 27376 1638 27432
rect 1582 26732 1584 26752
rect 1584 26732 1636 26752
rect 1636 26732 1638 26752
rect 1582 26696 1638 26732
rect 1582 26016 1638 26072
rect 1582 25336 1638 25392
rect 1582 24676 1638 24712
rect 1582 24656 1584 24676
rect 1584 24656 1636 24676
rect 1636 24656 1638 24676
rect 1582 24012 1584 24032
rect 1584 24012 1636 24032
rect 1636 24012 1638 24032
rect 1582 23976 1638 24012
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 1582 22752 1638 22808
rect 1582 22072 1638 22128
rect 1582 21412 1638 21448
rect 1582 21392 1584 21412
rect 1584 21392 1636 21412
rect 1636 21392 1638 21412
rect 1582 20748 1584 20768
rect 1584 20748 1636 20768
rect 1636 20748 1638 20768
rect 1582 20712 1638 20748
rect 1582 20032 1638 20088
rect 1582 19352 1638 19408
rect 1582 18808 1638 18864
rect 1582 18148 1638 18184
rect 1582 18128 1584 18148
rect 1584 18128 1636 18148
rect 1636 18128 1638 18148
rect 1582 17484 1584 17504
rect 1584 17484 1636 17504
rect 1636 17484 1638 17504
rect 1582 17448 1638 17484
rect 1582 16768 1638 16824
rect 1582 16088 1638 16144
rect 1582 15408 1638 15464
rect 1582 14764 1584 14784
rect 1584 14764 1636 14784
rect 1636 14764 1638 14784
rect 1582 14728 1638 14764
rect 1582 14220 1584 14240
rect 1584 14220 1636 14240
rect 1636 14220 1638 14240
rect 1582 14184 1638 14220
rect 1582 13504 1638 13560
rect 1582 12824 1638 12880
rect 1582 12144 1638 12200
rect 1582 11500 1584 11520
rect 1584 11500 1636 11520
rect 1636 11500 1638 11520
rect 1582 11464 1638 11500
rect 1582 10784 1638 10840
rect 1582 10104 1638 10160
rect 1582 9560 1638 9616
rect 1582 8880 1638 8936
rect 1582 8200 1638 8256
rect 1858 44512 1914 44568
rect 1858 43832 1914 43888
rect 1858 43152 1914 43208
rect 1858 40568 1914 40624
rect 1858 39208 1914 39264
rect 1582 7520 1638 7576
rect 1582 6840 1638 6896
rect 1582 6180 1638 6216
rect 1582 6160 1584 6180
rect 1584 6160 1636 6180
rect 1636 6160 1638 6180
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 1582 5480 1638 5516
rect 2588 73466 2644 73468
rect 2668 73466 2724 73468
rect 2748 73466 2804 73468
rect 2828 73466 2884 73468
rect 2588 73414 2634 73466
rect 2634 73414 2644 73466
rect 2668 73414 2698 73466
rect 2698 73414 2710 73466
rect 2710 73414 2724 73466
rect 2748 73414 2762 73466
rect 2762 73414 2774 73466
rect 2774 73414 2804 73466
rect 2828 73414 2838 73466
rect 2838 73414 2884 73466
rect 2588 73412 2644 73414
rect 2668 73412 2724 73414
rect 2748 73412 2804 73414
rect 2828 73412 2884 73414
rect 2870 72936 2926 72992
rect 2588 72378 2644 72380
rect 2668 72378 2724 72380
rect 2748 72378 2804 72380
rect 2828 72378 2884 72380
rect 2588 72326 2634 72378
rect 2634 72326 2644 72378
rect 2668 72326 2698 72378
rect 2698 72326 2710 72378
rect 2710 72326 2724 72378
rect 2748 72326 2762 72378
rect 2762 72326 2774 72378
rect 2774 72326 2804 72378
rect 2828 72326 2838 72378
rect 2838 72326 2884 72378
rect 2588 72324 2644 72326
rect 2668 72324 2724 72326
rect 2748 72324 2804 72326
rect 2828 72324 2884 72326
rect 2588 71290 2644 71292
rect 2668 71290 2724 71292
rect 2748 71290 2804 71292
rect 2828 71290 2884 71292
rect 2588 71238 2634 71290
rect 2634 71238 2644 71290
rect 2668 71238 2698 71290
rect 2698 71238 2710 71290
rect 2710 71238 2724 71290
rect 2748 71238 2762 71290
rect 2762 71238 2774 71290
rect 2774 71238 2804 71290
rect 2828 71238 2838 71290
rect 2838 71238 2884 71290
rect 2588 71236 2644 71238
rect 2668 71236 2724 71238
rect 2748 71236 2804 71238
rect 2828 71236 2884 71238
rect 2588 70202 2644 70204
rect 2668 70202 2724 70204
rect 2748 70202 2804 70204
rect 2828 70202 2884 70204
rect 2588 70150 2634 70202
rect 2634 70150 2644 70202
rect 2668 70150 2698 70202
rect 2698 70150 2710 70202
rect 2710 70150 2724 70202
rect 2748 70150 2762 70202
rect 2762 70150 2774 70202
rect 2774 70150 2804 70202
rect 2828 70150 2838 70202
rect 2838 70150 2884 70202
rect 2588 70148 2644 70150
rect 2668 70148 2724 70150
rect 2748 70148 2804 70150
rect 2828 70148 2884 70150
rect 2870 69264 2926 69320
rect 2588 69114 2644 69116
rect 2668 69114 2724 69116
rect 2748 69114 2804 69116
rect 2828 69114 2884 69116
rect 2588 69062 2634 69114
rect 2634 69062 2644 69114
rect 2668 69062 2698 69114
rect 2698 69062 2710 69114
rect 2710 69062 2724 69114
rect 2748 69062 2762 69114
rect 2762 69062 2774 69114
rect 2774 69062 2804 69114
rect 2828 69062 2838 69114
rect 2838 69062 2884 69114
rect 2588 69060 2644 69062
rect 2668 69060 2724 69062
rect 2748 69060 2804 69062
rect 2828 69060 2884 69062
rect 5851 77818 5907 77820
rect 5931 77818 5987 77820
rect 6011 77818 6067 77820
rect 6091 77818 6147 77820
rect 5851 77766 5897 77818
rect 5897 77766 5907 77818
rect 5931 77766 5961 77818
rect 5961 77766 5973 77818
rect 5973 77766 5987 77818
rect 6011 77766 6025 77818
rect 6025 77766 6037 77818
rect 6037 77766 6067 77818
rect 6091 77766 6101 77818
rect 6101 77766 6147 77818
rect 5851 77764 5907 77766
rect 5931 77764 5987 77766
rect 6011 77764 6067 77766
rect 6091 77764 6147 77766
rect 8574 79192 8630 79248
rect 8206 78240 8262 78296
rect 4219 77274 4275 77276
rect 4299 77274 4355 77276
rect 4379 77274 4435 77276
rect 4459 77274 4515 77276
rect 4219 77222 4265 77274
rect 4265 77222 4275 77274
rect 4299 77222 4329 77274
rect 4329 77222 4341 77274
rect 4341 77222 4355 77274
rect 4379 77222 4393 77274
rect 4393 77222 4405 77274
rect 4405 77222 4435 77274
rect 4459 77222 4469 77274
rect 4469 77222 4515 77274
rect 4219 77220 4275 77222
rect 4299 77220 4355 77222
rect 4379 77220 4435 77222
rect 4459 77220 4515 77222
rect 2588 68026 2644 68028
rect 2668 68026 2724 68028
rect 2748 68026 2804 68028
rect 2828 68026 2884 68028
rect 2588 67974 2634 68026
rect 2634 67974 2644 68026
rect 2668 67974 2698 68026
rect 2698 67974 2710 68026
rect 2710 67974 2724 68026
rect 2748 67974 2762 68026
rect 2762 67974 2774 68026
rect 2774 67974 2804 68026
rect 2828 67974 2838 68026
rect 2838 67974 2884 68026
rect 2588 67972 2644 67974
rect 2668 67972 2724 67974
rect 2748 67972 2804 67974
rect 2828 67972 2884 67974
rect 2588 66938 2644 66940
rect 2668 66938 2724 66940
rect 2748 66938 2804 66940
rect 2828 66938 2884 66940
rect 2588 66886 2634 66938
rect 2634 66886 2644 66938
rect 2668 66886 2698 66938
rect 2698 66886 2710 66938
rect 2710 66886 2724 66938
rect 2748 66886 2762 66938
rect 2762 66886 2774 66938
rect 2774 66886 2804 66938
rect 2828 66886 2838 66938
rect 2838 66886 2884 66938
rect 2588 66884 2644 66886
rect 2668 66884 2724 66886
rect 2748 66884 2804 66886
rect 2828 66884 2884 66886
rect 2962 66272 3018 66328
rect 5851 76730 5907 76732
rect 5931 76730 5987 76732
rect 6011 76730 6067 76732
rect 6091 76730 6147 76732
rect 5851 76678 5897 76730
rect 5897 76678 5907 76730
rect 5931 76678 5961 76730
rect 5961 76678 5973 76730
rect 5973 76678 5987 76730
rect 6011 76678 6025 76730
rect 6025 76678 6037 76730
rect 6037 76678 6067 76730
rect 6091 76678 6101 76730
rect 6101 76678 6147 76730
rect 5851 76676 5907 76678
rect 5931 76676 5987 76678
rect 6011 76676 6067 76678
rect 6091 76676 6147 76678
rect 4219 76186 4275 76188
rect 4299 76186 4355 76188
rect 4379 76186 4435 76188
rect 4459 76186 4515 76188
rect 4219 76134 4265 76186
rect 4265 76134 4275 76186
rect 4299 76134 4329 76186
rect 4329 76134 4341 76186
rect 4341 76134 4355 76186
rect 4379 76134 4393 76186
rect 4393 76134 4405 76186
rect 4405 76134 4435 76186
rect 4459 76134 4469 76186
rect 4469 76134 4515 76186
rect 4219 76132 4275 76134
rect 4299 76132 4355 76134
rect 4379 76132 4435 76134
rect 4459 76132 4515 76134
rect 5851 75642 5907 75644
rect 5931 75642 5987 75644
rect 6011 75642 6067 75644
rect 6091 75642 6147 75644
rect 5851 75590 5897 75642
rect 5897 75590 5907 75642
rect 5931 75590 5961 75642
rect 5961 75590 5973 75642
rect 5973 75590 5987 75642
rect 6011 75590 6025 75642
rect 6025 75590 6037 75642
rect 6037 75590 6067 75642
rect 6091 75590 6101 75642
rect 6101 75590 6147 75642
rect 5851 75588 5907 75590
rect 5931 75588 5987 75590
rect 6011 75588 6067 75590
rect 6091 75588 6147 75590
rect 4219 75098 4275 75100
rect 4299 75098 4355 75100
rect 4379 75098 4435 75100
rect 4459 75098 4515 75100
rect 4219 75046 4265 75098
rect 4265 75046 4275 75098
rect 4299 75046 4329 75098
rect 4329 75046 4341 75098
rect 4341 75046 4355 75098
rect 4379 75046 4393 75098
rect 4393 75046 4405 75098
rect 4405 75046 4435 75098
rect 4459 75046 4469 75098
rect 4469 75046 4515 75098
rect 4219 75044 4275 75046
rect 4299 75044 4355 75046
rect 4379 75044 4435 75046
rect 4459 75044 4515 75046
rect 4219 74010 4275 74012
rect 4299 74010 4355 74012
rect 4379 74010 4435 74012
rect 4459 74010 4515 74012
rect 4219 73958 4265 74010
rect 4265 73958 4275 74010
rect 4299 73958 4329 74010
rect 4329 73958 4341 74010
rect 4341 73958 4355 74010
rect 4379 73958 4393 74010
rect 4393 73958 4405 74010
rect 4405 73958 4435 74010
rect 4459 73958 4469 74010
rect 4469 73958 4515 74010
rect 4219 73956 4275 73958
rect 4299 73956 4355 73958
rect 4379 73956 4435 73958
rect 4459 73956 4515 73958
rect 4219 72922 4275 72924
rect 4299 72922 4355 72924
rect 4379 72922 4435 72924
rect 4459 72922 4515 72924
rect 4219 72870 4265 72922
rect 4265 72870 4275 72922
rect 4299 72870 4329 72922
rect 4329 72870 4341 72922
rect 4341 72870 4355 72922
rect 4379 72870 4393 72922
rect 4393 72870 4405 72922
rect 4405 72870 4435 72922
rect 4459 72870 4469 72922
rect 4469 72870 4515 72922
rect 4219 72868 4275 72870
rect 4299 72868 4355 72870
rect 4379 72868 4435 72870
rect 4459 72868 4515 72870
rect 2588 65850 2644 65852
rect 2668 65850 2724 65852
rect 2748 65850 2804 65852
rect 2828 65850 2884 65852
rect 2588 65798 2634 65850
rect 2634 65798 2644 65850
rect 2668 65798 2698 65850
rect 2698 65798 2710 65850
rect 2710 65798 2724 65850
rect 2748 65798 2762 65850
rect 2762 65798 2774 65850
rect 2774 65798 2804 65850
rect 2828 65798 2838 65850
rect 2838 65798 2884 65850
rect 2588 65796 2644 65798
rect 2668 65796 2724 65798
rect 2748 65796 2804 65798
rect 2828 65796 2884 65798
rect 2588 64762 2644 64764
rect 2668 64762 2724 64764
rect 2748 64762 2804 64764
rect 2828 64762 2884 64764
rect 2588 64710 2634 64762
rect 2634 64710 2644 64762
rect 2668 64710 2698 64762
rect 2698 64710 2710 64762
rect 2710 64710 2724 64762
rect 2748 64710 2762 64762
rect 2762 64710 2774 64762
rect 2774 64710 2804 64762
rect 2828 64710 2838 64762
rect 2838 64710 2884 64762
rect 2588 64708 2644 64710
rect 2668 64708 2724 64710
rect 2748 64708 2804 64710
rect 2828 64708 2884 64710
rect 2588 63674 2644 63676
rect 2668 63674 2724 63676
rect 2748 63674 2804 63676
rect 2828 63674 2884 63676
rect 2588 63622 2634 63674
rect 2634 63622 2644 63674
rect 2668 63622 2698 63674
rect 2698 63622 2710 63674
rect 2710 63622 2724 63674
rect 2748 63622 2762 63674
rect 2762 63622 2774 63674
rect 2774 63622 2804 63674
rect 2828 63622 2838 63674
rect 2838 63622 2884 63674
rect 2588 63620 2644 63622
rect 2668 63620 2724 63622
rect 2748 63620 2804 63622
rect 2828 63620 2884 63622
rect 2594 62736 2650 62792
rect 2588 62586 2644 62588
rect 2668 62586 2724 62588
rect 2748 62586 2804 62588
rect 2828 62586 2884 62588
rect 2588 62534 2634 62586
rect 2634 62534 2644 62586
rect 2668 62534 2698 62586
rect 2698 62534 2710 62586
rect 2710 62534 2724 62586
rect 2748 62534 2762 62586
rect 2762 62534 2774 62586
rect 2774 62534 2804 62586
rect 2828 62534 2838 62586
rect 2838 62534 2884 62586
rect 2588 62532 2644 62534
rect 2668 62532 2724 62534
rect 2748 62532 2804 62534
rect 2828 62532 2884 62534
rect 2588 61498 2644 61500
rect 2668 61498 2724 61500
rect 2748 61498 2804 61500
rect 2828 61498 2884 61500
rect 2588 61446 2634 61498
rect 2634 61446 2644 61498
rect 2668 61446 2698 61498
rect 2698 61446 2710 61498
rect 2710 61446 2724 61498
rect 2748 61446 2762 61498
rect 2762 61446 2774 61498
rect 2774 61446 2804 61498
rect 2828 61446 2838 61498
rect 2838 61446 2884 61498
rect 2588 61444 2644 61446
rect 2668 61444 2724 61446
rect 2748 61444 2804 61446
rect 2828 61444 2884 61446
rect 2778 60560 2834 60616
rect 2588 60410 2644 60412
rect 2668 60410 2724 60412
rect 2748 60410 2804 60412
rect 2828 60410 2884 60412
rect 2588 60358 2634 60410
rect 2634 60358 2644 60410
rect 2668 60358 2698 60410
rect 2698 60358 2710 60410
rect 2710 60358 2724 60410
rect 2748 60358 2762 60410
rect 2762 60358 2774 60410
rect 2774 60358 2804 60410
rect 2828 60358 2838 60410
rect 2838 60358 2884 60410
rect 2588 60356 2644 60358
rect 2668 60356 2724 60358
rect 2748 60356 2804 60358
rect 2828 60356 2884 60358
rect 2588 59322 2644 59324
rect 2668 59322 2724 59324
rect 2748 59322 2804 59324
rect 2828 59322 2884 59324
rect 2588 59270 2634 59322
rect 2634 59270 2644 59322
rect 2668 59270 2698 59322
rect 2698 59270 2710 59322
rect 2710 59270 2724 59322
rect 2748 59270 2762 59322
rect 2762 59270 2774 59322
rect 2774 59270 2804 59322
rect 2828 59270 2838 59322
rect 2838 59270 2884 59322
rect 2588 59268 2644 59270
rect 2668 59268 2724 59270
rect 2748 59268 2804 59270
rect 2828 59268 2884 59270
rect 2588 58234 2644 58236
rect 2668 58234 2724 58236
rect 2748 58234 2804 58236
rect 2828 58234 2884 58236
rect 2588 58182 2634 58234
rect 2634 58182 2644 58234
rect 2668 58182 2698 58234
rect 2698 58182 2710 58234
rect 2710 58182 2724 58234
rect 2748 58182 2762 58234
rect 2762 58182 2774 58234
rect 2774 58182 2804 58234
rect 2828 58182 2838 58234
rect 2838 58182 2884 58234
rect 2588 58180 2644 58182
rect 2668 58180 2724 58182
rect 2748 58180 2804 58182
rect 2828 58180 2884 58182
rect 2588 57146 2644 57148
rect 2668 57146 2724 57148
rect 2748 57146 2804 57148
rect 2828 57146 2884 57148
rect 2588 57094 2634 57146
rect 2634 57094 2644 57146
rect 2668 57094 2698 57146
rect 2698 57094 2710 57146
rect 2710 57094 2724 57146
rect 2748 57094 2762 57146
rect 2762 57094 2774 57146
rect 2774 57094 2804 57146
rect 2828 57094 2838 57146
rect 2838 57094 2884 57146
rect 2588 57092 2644 57094
rect 2668 57092 2724 57094
rect 2748 57092 2804 57094
rect 2828 57092 2884 57094
rect 2588 56058 2644 56060
rect 2668 56058 2724 56060
rect 2748 56058 2804 56060
rect 2828 56058 2884 56060
rect 2588 56006 2634 56058
rect 2634 56006 2644 56058
rect 2668 56006 2698 56058
rect 2698 56006 2710 56058
rect 2710 56006 2724 56058
rect 2748 56006 2762 56058
rect 2762 56006 2774 56058
rect 2774 56006 2804 56058
rect 2828 56006 2838 56058
rect 2838 56006 2884 56058
rect 2588 56004 2644 56006
rect 2668 56004 2724 56006
rect 2748 56004 2804 56006
rect 2828 56004 2884 56006
rect 2588 54970 2644 54972
rect 2668 54970 2724 54972
rect 2748 54970 2804 54972
rect 2828 54970 2884 54972
rect 2588 54918 2634 54970
rect 2634 54918 2644 54970
rect 2668 54918 2698 54970
rect 2698 54918 2710 54970
rect 2710 54918 2724 54970
rect 2748 54918 2762 54970
rect 2762 54918 2774 54970
rect 2774 54918 2804 54970
rect 2828 54918 2838 54970
rect 2838 54918 2884 54970
rect 2588 54916 2644 54918
rect 2668 54916 2724 54918
rect 2748 54916 2804 54918
rect 2828 54916 2884 54918
rect 2588 53882 2644 53884
rect 2668 53882 2724 53884
rect 2748 53882 2804 53884
rect 2828 53882 2884 53884
rect 2588 53830 2634 53882
rect 2634 53830 2644 53882
rect 2668 53830 2698 53882
rect 2698 53830 2710 53882
rect 2710 53830 2724 53882
rect 2748 53830 2762 53882
rect 2762 53830 2774 53882
rect 2774 53830 2804 53882
rect 2828 53830 2838 53882
rect 2838 53830 2884 53882
rect 2588 53828 2644 53830
rect 2668 53828 2724 53830
rect 2748 53828 2804 53830
rect 2828 53828 2884 53830
rect 2588 52794 2644 52796
rect 2668 52794 2724 52796
rect 2748 52794 2804 52796
rect 2828 52794 2884 52796
rect 2588 52742 2634 52794
rect 2634 52742 2644 52794
rect 2668 52742 2698 52794
rect 2698 52742 2710 52794
rect 2710 52742 2724 52794
rect 2748 52742 2762 52794
rect 2762 52742 2774 52794
rect 2774 52742 2804 52794
rect 2828 52742 2838 52794
rect 2838 52742 2884 52794
rect 2588 52740 2644 52742
rect 2668 52740 2724 52742
rect 2748 52740 2804 52742
rect 2828 52740 2884 52742
rect 2778 52400 2834 52456
rect 2588 51706 2644 51708
rect 2668 51706 2724 51708
rect 2748 51706 2804 51708
rect 2828 51706 2884 51708
rect 2588 51654 2634 51706
rect 2634 51654 2644 51706
rect 2668 51654 2698 51706
rect 2698 51654 2710 51706
rect 2710 51654 2724 51706
rect 2748 51654 2762 51706
rect 2762 51654 2774 51706
rect 2774 51654 2804 51706
rect 2828 51654 2838 51706
rect 2838 51654 2884 51706
rect 2588 51652 2644 51654
rect 2668 51652 2724 51654
rect 2748 51652 2804 51654
rect 2828 51652 2884 51654
rect 3054 51176 3110 51232
rect 3146 50904 3202 50960
rect 2226 39480 2282 39536
rect 2588 50618 2644 50620
rect 2668 50618 2724 50620
rect 2748 50618 2804 50620
rect 2828 50618 2884 50620
rect 2588 50566 2634 50618
rect 2634 50566 2644 50618
rect 2668 50566 2698 50618
rect 2698 50566 2710 50618
rect 2710 50566 2724 50618
rect 2748 50566 2762 50618
rect 2762 50566 2774 50618
rect 2774 50566 2804 50618
rect 2828 50566 2838 50618
rect 2838 50566 2884 50618
rect 2588 50564 2644 50566
rect 2668 50564 2724 50566
rect 2748 50564 2804 50566
rect 2828 50564 2884 50566
rect 2588 49530 2644 49532
rect 2668 49530 2724 49532
rect 2748 49530 2804 49532
rect 2828 49530 2884 49532
rect 2588 49478 2634 49530
rect 2634 49478 2644 49530
rect 2668 49478 2698 49530
rect 2698 49478 2710 49530
rect 2710 49478 2724 49530
rect 2748 49478 2762 49530
rect 2762 49478 2774 49530
rect 2774 49478 2804 49530
rect 2828 49478 2838 49530
rect 2838 49478 2884 49530
rect 2588 49476 2644 49478
rect 2668 49476 2724 49478
rect 2748 49476 2804 49478
rect 2828 49476 2884 49478
rect 2588 48442 2644 48444
rect 2668 48442 2724 48444
rect 2748 48442 2804 48444
rect 2828 48442 2884 48444
rect 2588 48390 2634 48442
rect 2634 48390 2644 48442
rect 2668 48390 2698 48442
rect 2698 48390 2710 48442
rect 2710 48390 2724 48442
rect 2748 48390 2762 48442
rect 2762 48390 2774 48442
rect 2774 48390 2804 48442
rect 2828 48390 2838 48442
rect 2838 48390 2884 48442
rect 2588 48388 2644 48390
rect 2668 48388 2724 48390
rect 2748 48388 2804 48390
rect 2828 48388 2884 48390
rect 2502 47504 2558 47560
rect 2588 47354 2644 47356
rect 2668 47354 2724 47356
rect 2748 47354 2804 47356
rect 2828 47354 2884 47356
rect 2588 47302 2634 47354
rect 2634 47302 2644 47354
rect 2668 47302 2698 47354
rect 2698 47302 2710 47354
rect 2710 47302 2724 47354
rect 2748 47302 2762 47354
rect 2762 47302 2774 47354
rect 2774 47302 2804 47354
rect 2828 47302 2838 47354
rect 2838 47302 2884 47354
rect 2588 47300 2644 47302
rect 2668 47300 2724 47302
rect 2748 47300 2804 47302
rect 2828 47300 2884 47302
rect 2588 46266 2644 46268
rect 2668 46266 2724 46268
rect 2748 46266 2804 46268
rect 2828 46266 2884 46268
rect 2588 46214 2634 46266
rect 2634 46214 2644 46266
rect 2668 46214 2698 46266
rect 2698 46214 2710 46266
rect 2710 46214 2724 46266
rect 2748 46214 2762 46266
rect 2762 46214 2774 46266
rect 2774 46214 2804 46266
rect 2828 46214 2838 46266
rect 2838 46214 2884 46266
rect 2588 46212 2644 46214
rect 2668 46212 2724 46214
rect 2748 46212 2804 46214
rect 2828 46212 2884 46214
rect 2588 45178 2644 45180
rect 2668 45178 2724 45180
rect 2748 45178 2804 45180
rect 2828 45178 2884 45180
rect 2588 45126 2634 45178
rect 2634 45126 2644 45178
rect 2668 45126 2698 45178
rect 2698 45126 2710 45178
rect 2710 45126 2724 45178
rect 2748 45126 2762 45178
rect 2762 45126 2774 45178
rect 2774 45126 2804 45178
rect 2828 45126 2838 45178
rect 2838 45126 2884 45178
rect 2588 45124 2644 45126
rect 2668 45124 2724 45126
rect 2748 45124 2804 45126
rect 2828 45124 2884 45126
rect 2588 44090 2644 44092
rect 2668 44090 2724 44092
rect 2748 44090 2804 44092
rect 2828 44090 2884 44092
rect 2588 44038 2634 44090
rect 2634 44038 2644 44090
rect 2668 44038 2698 44090
rect 2698 44038 2710 44090
rect 2710 44038 2724 44090
rect 2748 44038 2762 44090
rect 2762 44038 2774 44090
rect 2774 44038 2804 44090
rect 2828 44038 2838 44090
rect 2838 44038 2884 44090
rect 2588 44036 2644 44038
rect 2668 44036 2724 44038
rect 2748 44036 2804 44038
rect 2828 44036 2884 44038
rect 2588 43002 2644 43004
rect 2668 43002 2724 43004
rect 2748 43002 2804 43004
rect 2828 43002 2884 43004
rect 2588 42950 2634 43002
rect 2634 42950 2644 43002
rect 2668 42950 2698 43002
rect 2698 42950 2710 43002
rect 2710 42950 2724 43002
rect 2748 42950 2762 43002
rect 2762 42950 2774 43002
rect 2774 42950 2804 43002
rect 2828 42950 2838 43002
rect 2838 42950 2884 43002
rect 2588 42948 2644 42950
rect 2668 42948 2724 42950
rect 2748 42948 2804 42950
rect 2828 42948 2884 42950
rect 2588 41914 2644 41916
rect 2668 41914 2724 41916
rect 2748 41914 2804 41916
rect 2828 41914 2884 41916
rect 2588 41862 2634 41914
rect 2634 41862 2644 41914
rect 2668 41862 2698 41914
rect 2698 41862 2710 41914
rect 2710 41862 2724 41914
rect 2748 41862 2762 41914
rect 2762 41862 2774 41914
rect 2774 41862 2804 41914
rect 2828 41862 2838 41914
rect 2838 41862 2884 41914
rect 2588 41860 2644 41862
rect 2668 41860 2724 41862
rect 2748 41860 2804 41862
rect 2828 41860 2884 41862
rect 2588 40826 2644 40828
rect 2668 40826 2724 40828
rect 2748 40826 2804 40828
rect 2828 40826 2884 40828
rect 2588 40774 2634 40826
rect 2634 40774 2644 40826
rect 2668 40774 2698 40826
rect 2698 40774 2710 40826
rect 2710 40774 2724 40826
rect 2748 40774 2762 40826
rect 2762 40774 2774 40826
rect 2774 40774 2804 40826
rect 2828 40774 2838 40826
rect 2838 40774 2884 40826
rect 2588 40772 2644 40774
rect 2668 40772 2724 40774
rect 2748 40772 2804 40774
rect 2828 40772 2884 40774
rect 2588 39738 2644 39740
rect 2668 39738 2724 39740
rect 2748 39738 2804 39740
rect 2828 39738 2884 39740
rect 2588 39686 2634 39738
rect 2634 39686 2644 39738
rect 2668 39686 2698 39738
rect 2698 39686 2710 39738
rect 2710 39686 2724 39738
rect 2748 39686 2762 39738
rect 2762 39686 2774 39738
rect 2774 39686 2804 39738
rect 2828 39686 2838 39738
rect 2838 39686 2884 39738
rect 2588 39684 2644 39686
rect 2668 39684 2724 39686
rect 2748 39684 2804 39686
rect 2828 39684 2884 39686
rect 2588 38650 2644 38652
rect 2668 38650 2724 38652
rect 2748 38650 2804 38652
rect 2828 38650 2884 38652
rect 2588 38598 2634 38650
rect 2634 38598 2644 38650
rect 2668 38598 2698 38650
rect 2698 38598 2710 38650
rect 2710 38598 2724 38650
rect 2748 38598 2762 38650
rect 2762 38598 2774 38650
rect 2774 38598 2804 38650
rect 2828 38598 2838 38650
rect 2838 38598 2884 38650
rect 2588 38596 2644 38598
rect 2668 38596 2724 38598
rect 2748 38596 2804 38598
rect 2828 38596 2884 38598
rect 2686 37732 2742 37768
rect 2686 37712 2688 37732
rect 2688 37712 2740 37732
rect 2740 37712 2742 37732
rect 2588 37562 2644 37564
rect 2668 37562 2724 37564
rect 2748 37562 2804 37564
rect 2828 37562 2884 37564
rect 2588 37510 2634 37562
rect 2634 37510 2644 37562
rect 2668 37510 2698 37562
rect 2698 37510 2710 37562
rect 2710 37510 2724 37562
rect 2748 37510 2762 37562
rect 2762 37510 2774 37562
rect 2774 37510 2804 37562
rect 2828 37510 2838 37562
rect 2838 37510 2884 37562
rect 2588 37508 2644 37510
rect 2668 37508 2724 37510
rect 2748 37508 2804 37510
rect 2828 37508 2884 37510
rect 2588 36474 2644 36476
rect 2668 36474 2724 36476
rect 2748 36474 2804 36476
rect 2828 36474 2884 36476
rect 2588 36422 2634 36474
rect 2634 36422 2644 36474
rect 2668 36422 2698 36474
rect 2698 36422 2710 36474
rect 2710 36422 2724 36474
rect 2748 36422 2762 36474
rect 2762 36422 2774 36474
rect 2774 36422 2804 36474
rect 2828 36422 2838 36474
rect 2838 36422 2884 36474
rect 2588 36420 2644 36422
rect 2668 36420 2724 36422
rect 2748 36420 2804 36422
rect 2828 36420 2884 36422
rect 2588 35386 2644 35388
rect 2668 35386 2724 35388
rect 2748 35386 2804 35388
rect 2828 35386 2884 35388
rect 2588 35334 2634 35386
rect 2634 35334 2644 35386
rect 2668 35334 2698 35386
rect 2698 35334 2710 35386
rect 2710 35334 2724 35386
rect 2748 35334 2762 35386
rect 2762 35334 2774 35386
rect 2774 35334 2804 35386
rect 2828 35334 2838 35386
rect 2838 35334 2884 35386
rect 2588 35332 2644 35334
rect 2668 35332 2724 35334
rect 2748 35332 2804 35334
rect 2828 35332 2884 35334
rect 2588 34298 2644 34300
rect 2668 34298 2724 34300
rect 2748 34298 2804 34300
rect 2828 34298 2884 34300
rect 2588 34246 2634 34298
rect 2634 34246 2644 34298
rect 2668 34246 2698 34298
rect 2698 34246 2710 34298
rect 2710 34246 2724 34298
rect 2748 34246 2762 34298
rect 2762 34246 2774 34298
rect 2774 34246 2804 34298
rect 2828 34246 2838 34298
rect 2838 34246 2884 34298
rect 2588 34244 2644 34246
rect 2668 34244 2724 34246
rect 2748 34244 2804 34246
rect 2828 34244 2884 34246
rect 2588 33210 2644 33212
rect 2668 33210 2724 33212
rect 2748 33210 2804 33212
rect 2828 33210 2884 33212
rect 2588 33158 2634 33210
rect 2634 33158 2644 33210
rect 2668 33158 2698 33210
rect 2698 33158 2710 33210
rect 2710 33158 2724 33210
rect 2748 33158 2762 33210
rect 2762 33158 2774 33210
rect 2774 33158 2804 33210
rect 2828 33158 2838 33210
rect 2838 33158 2884 33210
rect 2588 33156 2644 33158
rect 2668 33156 2724 33158
rect 2748 33156 2804 33158
rect 2828 33156 2884 33158
rect 2588 32122 2644 32124
rect 2668 32122 2724 32124
rect 2748 32122 2804 32124
rect 2828 32122 2884 32124
rect 2588 32070 2634 32122
rect 2634 32070 2644 32122
rect 2668 32070 2698 32122
rect 2698 32070 2710 32122
rect 2710 32070 2724 32122
rect 2748 32070 2762 32122
rect 2762 32070 2774 32122
rect 2774 32070 2804 32122
rect 2828 32070 2838 32122
rect 2838 32070 2884 32122
rect 2588 32068 2644 32070
rect 2668 32068 2724 32070
rect 2748 32068 2804 32070
rect 2828 32068 2884 32070
rect 2588 31034 2644 31036
rect 2668 31034 2724 31036
rect 2748 31034 2804 31036
rect 2828 31034 2884 31036
rect 2588 30982 2634 31034
rect 2634 30982 2644 31034
rect 2668 30982 2698 31034
rect 2698 30982 2710 31034
rect 2710 30982 2724 31034
rect 2748 30982 2762 31034
rect 2762 30982 2774 31034
rect 2774 30982 2804 31034
rect 2828 30982 2838 31034
rect 2838 30982 2884 31034
rect 2588 30980 2644 30982
rect 2668 30980 2724 30982
rect 2748 30980 2804 30982
rect 2828 30980 2884 30982
rect 2588 29946 2644 29948
rect 2668 29946 2724 29948
rect 2748 29946 2804 29948
rect 2828 29946 2884 29948
rect 2588 29894 2634 29946
rect 2634 29894 2644 29946
rect 2668 29894 2698 29946
rect 2698 29894 2710 29946
rect 2710 29894 2724 29946
rect 2748 29894 2762 29946
rect 2762 29894 2774 29946
rect 2774 29894 2804 29946
rect 2828 29894 2838 29946
rect 2838 29894 2884 29946
rect 2588 29892 2644 29894
rect 2668 29892 2724 29894
rect 2748 29892 2804 29894
rect 2828 29892 2884 29894
rect 2588 28858 2644 28860
rect 2668 28858 2724 28860
rect 2748 28858 2804 28860
rect 2828 28858 2884 28860
rect 2588 28806 2634 28858
rect 2634 28806 2644 28858
rect 2668 28806 2698 28858
rect 2698 28806 2710 28858
rect 2710 28806 2724 28858
rect 2748 28806 2762 28858
rect 2762 28806 2774 28858
rect 2774 28806 2804 28858
rect 2828 28806 2838 28858
rect 2838 28806 2884 28858
rect 2588 28804 2644 28806
rect 2668 28804 2724 28806
rect 2748 28804 2804 28806
rect 2828 28804 2884 28806
rect 2588 27770 2644 27772
rect 2668 27770 2724 27772
rect 2748 27770 2804 27772
rect 2828 27770 2884 27772
rect 2588 27718 2634 27770
rect 2634 27718 2644 27770
rect 2668 27718 2698 27770
rect 2698 27718 2710 27770
rect 2710 27718 2724 27770
rect 2748 27718 2762 27770
rect 2762 27718 2774 27770
rect 2774 27718 2804 27770
rect 2828 27718 2838 27770
rect 2838 27718 2884 27770
rect 2588 27716 2644 27718
rect 2668 27716 2724 27718
rect 2748 27716 2804 27718
rect 2828 27716 2884 27718
rect 2588 26682 2644 26684
rect 2668 26682 2724 26684
rect 2748 26682 2804 26684
rect 2828 26682 2884 26684
rect 2588 26630 2634 26682
rect 2634 26630 2644 26682
rect 2668 26630 2698 26682
rect 2698 26630 2710 26682
rect 2710 26630 2724 26682
rect 2748 26630 2762 26682
rect 2762 26630 2774 26682
rect 2774 26630 2804 26682
rect 2828 26630 2838 26682
rect 2838 26630 2884 26682
rect 2588 26628 2644 26630
rect 2668 26628 2724 26630
rect 2748 26628 2804 26630
rect 2828 26628 2884 26630
rect 2588 25594 2644 25596
rect 2668 25594 2724 25596
rect 2748 25594 2804 25596
rect 2828 25594 2884 25596
rect 2588 25542 2634 25594
rect 2634 25542 2644 25594
rect 2668 25542 2698 25594
rect 2698 25542 2710 25594
rect 2710 25542 2724 25594
rect 2748 25542 2762 25594
rect 2762 25542 2774 25594
rect 2774 25542 2804 25594
rect 2828 25542 2838 25594
rect 2838 25542 2884 25594
rect 2588 25540 2644 25542
rect 2668 25540 2724 25542
rect 2748 25540 2804 25542
rect 2828 25540 2884 25542
rect 2588 24506 2644 24508
rect 2668 24506 2724 24508
rect 2748 24506 2804 24508
rect 2828 24506 2884 24508
rect 2588 24454 2634 24506
rect 2634 24454 2644 24506
rect 2668 24454 2698 24506
rect 2698 24454 2710 24506
rect 2710 24454 2724 24506
rect 2748 24454 2762 24506
rect 2762 24454 2774 24506
rect 2774 24454 2804 24506
rect 2828 24454 2838 24506
rect 2838 24454 2884 24506
rect 2588 24452 2644 24454
rect 2668 24452 2724 24454
rect 2748 24452 2804 24454
rect 2828 24452 2884 24454
rect 2588 23418 2644 23420
rect 2668 23418 2724 23420
rect 2748 23418 2804 23420
rect 2828 23418 2884 23420
rect 2588 23366 2634 23418
rect 2634 23366 2644 23418
rect 2668 23366 2698 23418
rect 2698 23366 2710 23418
rect 2710 23366 2724 23418
rect 2748 23366 2762 23418
rect 2762 23366 2774 23418
rect 2774 23366 2804 23418
rect 2828 23366 2838 23418
rect 2838 23366 2884 23418
rect 2588 23364 2644 23366
rect 2668 23364 2724 23366
rect 2748 23364 2804 23366
rect 2828 23364 2884 23366
rect 2588 22330 2644 22332
rect 2668 22330 2724 22332
rect 2748 22330 2804 22332
rect 2828 22330 2884 22332
rect 2588 22278 2634 22330
rect 2634 22278 2644 22330
rect 2668 22278 2698 22330
rect 2698 22278 2710 22330
rect 2710 22278 2724 22330
rect 2748 22278 2762 22330
rect 2762 22278 2774 22330
rect 2774 22278 2804 22330
rect 2828 22278 2838 22330
rect 2838 22278 2884 22330
rect 2588 22276 2644 22278
rect 2668 22276 2724 22278
rect 2748 22276 2804 22278
rect 2828 22276 2884 22278
rect 2588 21242 2644 21244
rect 2668 21242 2724 21244
rect 2748 21242 2804 21244
rect 2828 21242 2884 21244
rect 2588 21190 2634 21242
rect 2634 21190 2644 21242
rect 2668 21190 2698 21242
rect 2698 21190 2710 21242
rect 2710 21190 2724 21242
rect 2748 21190 2762 21242
rect 2762 21190 2774 21242
rect 2774 21190 2804 21242
rect 2828 21190 2838 21242
rect 2838 21190 2884 21242
rect 2588 21188 2644 21190
rect 2668 21188 2724 21190
rect 2748 21188 2804 21190
rect 2828 21188 2884 21190
rect 2588 20154 2644 20156
rect 2668 20154 2724 20156
rect 2748 20154 2804 20156
rect 2828 20154 2884 20156
rect 2588 20102 2634 20154
rect 2634 20102 2644 20154
rect 2668 20102 2698 20154
rect 2698 20102 2710 20154
rect 2710 20102 2724 20154
rect 2748 20102 2762 20154
rect 2762 20102 2774 20154
rect 2774 20102 2804 20154
rect 2828 20102 2838 20154
rect 2838 20102 2884 20154
rect 2588 20100 2644 20102
rect 2668 20100 2724 20102
rect 2748 20100 2804 20102
rect 2828 20100 2884 20102
rect 2588 19066 2644 19068
rect 2668 19066 2724 19068
rect 2748 19066 2804 19068
rect 2828 19066 2884 19068
rect 2588 19014 2634 19066
rect 2634 19014 2644 19066
rect 2668 19014 2698 19066
rect 2698 19014 2710 19066
rect 2710 19014 2724 19066
rect 2748 19014 2762 19066
rect 2762 19014 2774 19066
rect 2774 19014 2804 19066
rect 2828 19014 2838 19066
rect 2838 19014 2884 19066
rect 2588 19012 2644 19014
rect 2668 19012 2724 19014
rect 2748 19012 2804 19014
rect 2828 19012 2884 19014
rect 2588 17978 2644 17980
rect 2668 17978 2724 17980
rect 2748 17978 2804 17980
rect 2828 17978 2884 17980
rect 2588 17926 2634 17978
rect 2634 17926 2644 17978
rect 2668 17926 2698 17978
rect 2698 17926 2710 17978
rect 2710 17926 2724 17978
rect 2748 17926 2762 17978
rect 2762 17926 2774 17978
rect 2774 17926 2804 17978
rect 2828 17926 2838 17978
rect 2838 17926 2884 17978
rect 2588 17924 2644 17926
rect 2668 17924 2724 17926
rect 2748 17924 2804 17926
rect 2828 17924 2884 17926
rect 3974 69672 4030 69728
rect 3606 50904 3662 50960
rect 3698 49680 3754 49736
rect 3606 49544 3662 49600
rect 3790 49544 3846 49600
rect 3698 49408 3754 49464
rect 3790 45328 3846 45384
rect 4219 71834 4275 71836
rect 4299 71834 4355 71836
rect 4379 71834 4435 71836
rect 4459 71834 4515 71836
rect 4219 71782 4265 71834
rect 4265 71782 4275 71834
rect 4299 71782 4329 71834
rect 4329 71782 4341 71834
rect 4341 71782 4355 71834
rect 4379 71782 4393 71834
rect 4393 71782 4405 71834
rect 4405 71782 4435 71834
rect 4459 71782 4469 71834
rect 4469 71782 4515 71834
rect 4219 71780 4275 71782
rect 4299 71780 4355 71782
rect 4379 71780 4435 71782
rect 4459 71780 4515 71782
rect 5851 74554 5907 74556
rect 5931 74554 5987 74556
rect 6011 74554 6067 74556
rect 6091 74554 6147 74556
rect 5851 74502 5897 74554
rect 5897 74502 5907 74554
rect 5931 74502 5961 74554
rect 5961 74502 5973 74554
rect 5973 74502 5987 74554
rect 6011 74502 6025 74554
rect 6025 74502 6037 74554
rect 6037 74502 6067 74554
rect 6091 74502 6101 74554
rect 6101 74502 6147 74554
rect 5851 74500 5907 74502
rect 5931 74500 5987 74502
rect 6011 74500 6067 74502
rect 6091 74500 6147 74502
rect 7483 77274 7539 77276
rect 7563 77274 7619 77276
rect 7643 77274 7699 77276
rect 7723 77274 7779 77276
rect 7483 77222 7529 77274
rect 7529 77222 7539 77274
rect 7563 77222 7593 77274
rect 7593 77222 7605 77274
rect 7605 77222 7619 77274
rect 7643 77222 7657 77274
rect 7657 77222 7669 77274
rect 7669 77222 7699 77274
rect 7723 77222 7733 77274
rect 7733 77222 7779 77274
rect 7483 77220 7539 77222
rect 7563 77220 7619 77222
rect 7643 77220 7699 77222
rect 7723 77220 7779 77222
rect 9494 78648 9550 78704
rect 9115 77818 9171 77820
rect 9195 77818 9251 77820
rect 9275 77818 9331 77820
rect 9355 77818 9411 77820
rect 9115 77766 9161 77818
rect 9161 77766 9171 77818
rect 9195 77766 9225 77818
rect 9225 77766 9237 77818
rect 9237 77766 9251 77818
rect 9275 77766 9289 77818
rect 9289 77766 9301 77818
rect 9301 77766 9331 77818
rect 9355 77766 9365 77818
rect 9365 77766 9411 77818
rect 9115 77764 9171 77766
rect 9195 77764 9251 77766
rect 9275 77764 9331 77766
rect 9355 77764 9411 77766
rect 7483 76186 7539 76188
rect 7563 76186 7619 76188
rect 7643 76186 7699 76188
rect 7723 76186 7779 76188
rect 7483 76134 7529 76186
rect 7529 76134 7539 76186
rect 7563 76134 7593 76186
rect 7593 76134 7605 76186
rect 7605 76134 7619 76186
rect 7643 76134 7657 76186
rect 7657 76134 7669 76186
rect 7669 76134 7699 76186
rect 7723 76134 7733 76186
rect 7733 76134 7779 76186
rect 7483 76132 7539 76134
rect 7563 76132 7619 76134
rect 7643 76132 7699 76134
rect 7723 76132 7779 76134
rect 7483 75098 7539 75100
rect 7563 75098 7619 75100
rect 7643 75098 7699 75100
rect 7723 75098 7779 75100
rect 7483 75046 7529 75098
rect 7529 75046 7539 75098
rect 7563 75046 7593 75098
rect 7593 75046 7605 75098
rect 7605 75046 7619 75098
rect 7643 75046 7657 75098
rect 7657 75046 7669 75098
rect 7669 75046 7699 75098
rect 7723 75046 7733 75098
rect 7733 75046 7779 75098
rect 7483 75044 7539 75046
rect 7563 75044 7619 75046
rect 7643 75044 7699 75046
rect 7723 75044 7779 75046
rect 5851 73466 5907 73468
rect 5931 73466 5987 73468
rect 6011 73466 6067 73468
rect 6091 73466 6147 73468
rect 5851 73414 5897 73466
rect 5897 73414 5907 73466
rect 5931 73414 5961 73466
rect 5961 73414 5973 73466
rect 5973 73414 5987 73466
rect 6011 73414 6025 73466
rect 6025 73414 6037 73466
rect 6037 73414 6067 73466
rect 6091 73414 6101 73466
rect 6101 73414 6147 73466
rect 5851 73412 5907 73414
rect 5931 73412 5987 73414
rect 6011 73412 6067 73414
rect 6091 73412 6147 73414
rect 5851 72378 5907 72380
rect 5931 72378 5987 72380
rect 6011 72378 6067 72380
rect 6091 72378 6147 72380
rect 5851 72326 5897 72378
rect 5897 72326 5907 72378
rect 5931 72326 5961 72378
rect 5961 72326 5973 72378
rect 5973 72326 5987 72378
rect 6011 72326 6025 72378
rect 6025 72326 6037 72378
rect 6037 72326 6067 72378
rect 6091 72326 6101 72378
rect 6101 72326 6147 72378
rect 5851 72324 5907 72326
rect 5931 72324 5987 72326
rect 6011 72324 6067 72326
rect 6091 72324 6147 72326
rect 4219 70746 4275 70748
rect 4299 70746 4355 70748
rect 4379 70746 4435 70748
rect 4459 70746 4515 70748
rect 4219 70694 4265 70746
rect 4265 70694 4275 70746
rect 4299 70694 4329 70746
rect 4329 70694 4341 70746
rect 4341 70694 4355 70746
rect 4379 70694 4393 70746
rect 4393 70694 4405 70746
rect 4405 70694 4435 70746
rect 4459 70694 4469 70746
rect 4469 70694 4515 70746
rect 4219 70692 4275 70694
rect 4299 70692 4355 70694
rect 4379 70692 4435 70694
rect 4459 70692 4515 70694
rect 4219 69658 4275 69660
rect 4299 69658 4355 69660
rect 4379 69658 4435 69660
rect 4459 69658 4515 69660
rect 4219 69606 4265 69658
rect 4265 69606 4275 69658
rect 4299 69606 4329 69658
rect 4329 69606 4341 69658
rect 4341 69606 4355 69658
rect 4379 69606 4393 69658
rect 4393 69606 4405 69658
rect 4405 69606 4435 69658
rect 4459 69606 4469 69658
rect 4469 69606 4515 69658
rect 4219 69604 4275 69606
rect 4299 69604 4355 69606
rect 4379 69604 4435 69606
rect 4459 69604 4515 69606
rect 4219 68570 4275 68572
rect 4299 68570 4355 68572
rect 4379 68570 4435 68572
rect 4459 68570 4515 68572
rect 4219 68518 4265 68570
rect 4265 68518 4275 68570
rect 4299 68518 4329 68570
rect 4329 68518 4341 68570
rect 4341 68518 4355 68570
rect 4379 68518 4393 68570
rect 4393 68518 4405 68570
rect 4405 68518 4435 68570
rect 4459 68518 4469 68570
rect 4469 68518 4515 68570
rect 4219 68516 4275 68518
rect 4299 68516 4355 68518
rect 4379 68516 4435 68518
rect 4459 68516 4515 68518
rect 4219 67482 4275 67484
rect 4299 67482 4355 67484
rect 4379 67482 4435 67484
rect 4459 67482 4515 67484
rect 4219 67430 4265 67482
rect 4265 67430 4275 67482
rect 4299 67430 4329 67482
rect 4329 67430 4341 67482
rect 4341 67430 4355 67482
rect 4379 67430 4393 67482
rect 4393 67430 4405 67482
rect 4405 67430 4435 67482
rect 4459 67430 4469 67482
rect 4469 67430 4515 67482
rect 4219 67428 4275 67430
rect 4299 67428 4355 67430
rect 4379 67428 4435 67430
rect 4459 67428 4515 67430
rect 4219 66394 4275 66396
rect 4299 66394 4355 66396
rect 4379 66394 4435 66396
rect 4459 66394 4515 66396
rect 4219 66342 4265 66394
rect 4265 66342 4275 66394
rect 4299 66342 4329 66394
rect 4329 66342 4341 66394
rect 4341 66342 4355 66394
rect 4379 66342 4393 66394
rect 4393 66342 4405 66394
rect 4405 66342 4435 66394
rect 4459 66342 4469 66394
rect 4469 66342 4515 66394
rect 4219 66340 4275 66342
rect 4299 66340 4355 66342
rect 4379 66340 4435 66342
rect 4459 66340 4515 66342
rect 4219 65306 4275 65308
rect 4299 65306 4355 65308
rect 4379 65306 4435 65308
rect 4459 65306 4515 65308
rect 4219 65254 4265 65306
rect 4265 65254 4275 65306
rect 4299 65254 4329 65306
rect 4329 65254 4341 65306
rect 4341 65254 4355 65306
rect 4379 65254 4393 65306
rect 4393 65254 4405 65306
rect 4405 65254 4435 65306
rect 4459 65254 4469 65306
rect 4469 65254 4515 65306
rect 4219 65252 4275 65254
rect 4299 65252 4355 65254
rect 4379 65252 4435 65254
rect 4459 65252 4515 65254
rect 4219 64218 4275 64220
rect 4299 64218 4355 64220
rect 4379 64218 4435 64220
rect 4459 64218 4515 64220
rect 4219 64166 4265 64218
rect 4265 64166 4275 64218
rect 4299 64166 4329 64218
rect 4329 64166 4341 64218
rect 4341 64166 4355 64218
rect 4379 64166 4393 64218
rect 4393 64166 4405 64218
rect 4405 64166 4435 64218
rect 4459 64166 4469 64218
rect 4469 64166 4515 64218
rect 4219 64164 4275 64166
rect 4299 64164 4355 64166
rect 4379 64164 4435 64166
rect 4459 64164 4515 64166
rect 4219 63130 4275 63132
rect 4299 63130 4355 63132
rect 4379 63130 4435 63132
rect 4459 63130 4515 63132
rect 4219 63078 4265 63130
rect 4265 63078 4275 63130
rect 4299 63078 4329 63130
rect 4329 63078 4341 63130
rect 4341 63078 4355 63130
rect 4379 63078 4393 63130
rect 4393 63078 4405 63130
rect 4405 63078 4435 63130
rect 4459 63078 4469 63130
rect 4469 63078 4515 63130
rect 4219 63076 4275 63078
rect 4299 63076 4355 63078
rect 4379 63076 4435 63078
rect 4459 63076 4515 63078
rect 4219 62042 4275 62044
rect 4299 62042 4355 62044
rect 4379 62042 4435 62044
rect 4459 62042 4515 62044
rect 4219 61990 4265 62042
rect 4265 61990 4275 62042
rect 4299 61990 4329 62042
rect 4329 61990 4341 62042
rect 4341 61990 4355 62042
rect 4379 61990 4393 62042
rect 4393 61990 4405 62042
rect 4405 61990 4435 62042
rect 4459 61990 4469 62042
rect 4469 61990 4515 62042
rect 4219 61988 4275 61990
rect 4299 61988 4355 61990
rect 4379 61988 4435 61990
rect 4459 61988 4515 61990
rect 4219 60954 4275 60956
rect 4299 60954 4355 60956
rect 4379 60954 4435 60956
rect 4459 60954 4515 60956
rect 4219 60902 4265 60954
rect 4265 60902 4275 60954
rect 4299 60902 4329 60954
rect 4329 60902 4341 60954
rect 4341 60902 4355 60954
rect 4379 60902 4393 60954
rect 4393 60902 4405 60954
rect 4405 60902 4435 60954
rect 4459 60902 4469 60954
rect 4469 60902 4515 60954
rect 4219 60900 4275 60902
rect 4299 60900 4355 60902
rect 4379 60900 4435 60902
rect 4459 60900 4515 60902
rect 4219 59866 4275 59868
rect 4299 59866 4355 59868
rect 4379 59866 4435 59868
rect 4459 59866 4515 59868
rect 4219 59814 4265 59866
rect 4265 59814 4275 59866
rect 4299 59814 4329 59866
rect 4329 59814 4341 59866
rect 4341 59814 4355 59866
rect 4379 59814 4393 59866
rect 4393 59814 4405 59866
rect 4405 59814 4435 59866
rect 4459 59814 4469 59866
rect 4469 59814 4515 59866
rect 4219 59812 4275 59814
rect 4299 59812 4355 59814
rect 4379 59812 4435 59814
rect 4459 59812 4515 59814
rect 4219 58778 4275 58780
rect 4299 58778 4355 58780
rect 4379 58778 4435 58780
rect 4459 58778 4515 58780
rect 4219 58726 4265 58778
rect 4265 58726 4275 58778
rect 4299 58726 4329 58778
rect 4329 58726 4341 58778
rect 4341 58726 4355 58778
rect 4379 58726 4393 58778
rect 4393 58726 4405 58778
rect 4405 58726 4435 58778
rect 4459 58726 4469 58778
rect 4469 58726 4515 58778
rect 4219 58724 4275 58726
rect 4299 58724 4355 58726
rect 4379 58724 4435 58726
rect 4459 58724 4515 58726
rect 4219 57690 4275 57692
rect 4299 57690 4355 57692
rect 4379 57690 4435 57692
rect 4459 57690 4515 57692
rect 4219 57638 4265 57690
rect 4265 57638 4275 57690
rect 4299 57638 4329 57690
rect 4329 57638 4341 57690
rect 4341 57638 4355 57690
rect 4379 57638 4393 57690
rect 4393 57638 4405 57690
rect 4405 57638 4435 57690
rect 4459 57638 4469 57690
rect 4469 57638 4515 57690
rect 4219 57636 4275 57638
rect 4299 57636 4355 57638
rect 4379 57636 4435 57638
rect 4459 57636 4515 57638
rect 4219 56602 4275 56604
rect 4299 56602 4355 56604
rect 4379 56602 4435 56604
rect 4459 56602 4515 56604
rect 4219 56550 4265 56602
rect 4265 56550 4275 56602
rect 4299 56550 4329 56602
rect 4329 56550 4341 56602
rect 4341 56550 4355 56602
rect 4379 56550 4393 56602
rect 4393 56550 4405 56602
rect 4405 56550 4435 56602
rect 4459 56550 4469 56602
rect 4469 56550 4515 56602
rect 4219 56548 4275 56550
rect 4299 56548 4355 56550
rect 4379 56548 4435 56550
rect 4459 56548 4515 56550
rect 4219 55514 4275 55516
rect 4299 55514 4355 55516
rect 4379 55514 4435 55516
rect 4459 55514 4515 55516
rect 4219 55462 4265 55514
rect 4265 55462 4275 55514
rect 4299 55462 4329 55514
rect 4329 55462 4341 55514
rect 4341 55462 4355 55514
rect 4379 55462 4393 55514
rect 4393 55462 4405 55514
rect 4405 55462 4435 55514
rect 4459 55462 4469 55514
rect 4469 55462 4515 55514
rect 4219 55460 4275 55462
rect 4299 55460 4355 55462
rect 4379 55460 4435 55462
rect 4459 55460 4515 55462
rect 4219 54426 4275 54428
rect 4299 54426 4355 54428
rect 4379 54426 4435 54428
rect 4459 54426 4515 54428
rect 4219 54374 4265 54426
rect 4265 54374 4275 54426
rect 4299 54374 4329 54426
rect 4329 54374 4341 54426
rect 4341 54374 4355 54426
rect 4379 54374 4393 54426
rect 4393 54374 4405 54426
rect 4405 54374 4435 54426
rect 4459 54374 4469 54426
rect 4469 54374 4515 54426
rect 4219 54372 4275 54374
rect 4299 54372 4355 54374
rect 4379 54372 4435 54374
rect 4459 54372 4515 54374
rect 4219 53338 4275 53340
rect 4299 53338 4355 53340
rect 4379 53338 4435 53340
rect 4459 53338 4515 53340
rect 4219 53286 4265 53338
rect 4265 53286 4275 53338
rect 4299 53286 4329 53338
rect 4329 53286 4341 53338
rect 4341 53286 4355 53338
rect 4379 53286 4393 53338
rect 4393 53286 4405 53338
rect 4405 53286 4435 53338
rect 4459 53286 4469 53338
rect 4469 53286 4515 53338
rect 4219 53284 4275 53286
rect 4299 53284 4355 53286
rect 4379 53284 4435 53286
rect 4459 53284 4515 53286
rect 4219 52250 4275 52252
rect 4299 52250 4355 52252
rect 4379 52250 4435 52252
rect 4459 52250 4515 52252
rect 4219 52198 4265 52250
rect 4265 52198 4275 52250
rect 4299 52198 4329 52250
rect 4329 52198 4341 52250
rect 4341 52198 4355 52250
rect 4379 52198 4393 52250
rect 4393 52198 4405 52250
rect 4405 52198 4435 52250
rect 4459 52198 4469 52250
rect 4469 52198 4515 52250
rect 4219 52196 4275 52198
rect 4299 52196 4355 52198
rect 4379 52196 4435 52198
rect 4459 52196 4515 52198
rect 4219 51162 4275 51164
rect 4299 51162 4355 51164
rect 4379 51162 4435 51164
rect 4459 51162 4515 51164
rect 4219 51110 4265 51162
rect 4265 51110 4275 51162
rect 4299 51110 4329 51162
rect 4329 51110 4341 51162
rect 4341 51110 4355 51162
rect 4379 51110 4393 51162
rect 4393 51110 4405 51162
rect 4405 51110 4435 51162
rect 4459 51110 4469 51162
rect 4469 51110 4515 51162
rect 4219 51108 4275 51110
rect 4299 51108 4355 51110
rect 4379 51108 4435 51110
rect 4459 51108 4515 51110
rect 4219 50074 4275 50076
rect 4299 50074 4355 50076
rect 4379 50074 4435 50076
rect 4459 50074 4515 50076
rect 4219 50022 4265 50074
rect 4265 50022 4275 50074
rect 4299 50022 4329 50074
rect 4329 50022 4341 50074
rect 4341 50022 4355 50074
rect 4379 50022 4393 50074
rect 4393 50022 4405 50074
rect 4405 50022 4435 50074
rect 4459 50022 4469 50074
rect 4469 50022 4515 50074
rect 4219 50020 4275 50022
rect 4299 50020 4355 50022
rect 4379 50020 4435 50022
rect 4459 50020 4515 50022
rect 4219 48986 4275 48988
rect 4299 48986 4355 48988
rect 4379 48986 4435 48988
rect 4459 48986 4515 48988
rect 4219 48934 4265 48986
rect 4265 48934 4275 48986
rect 4299 48934 4329 48986
rect 4329 48934 4341 48986
rect 4341 48934 4355 48986
rect 4379 48934 4393 48986
rect 4393 48934 4405 48986
rect 4405 48934 4435 48986
rect 4459 48934 4469 48986
rect 4469 48934 4515 48986
rect 4219 48932 4275 48934
rect 4299 48932 4355 48934
rect 4379 48932 4435 48934
rect 4459 48932 4515 48934
rect 4219 47898 4275 47900
rect 4299 47898 4355 47900
rect 4379 47898 4435 47900
rect 4459 47898 4515 47900
rect 4219 47846 4265 47898
rect 4265 47846 4275 47898
rect 4299 47846 4329 47898
rect 4329 47846 4341 47898
rect 4341 47846 4355 47898
rect 4379 47846 4393 47898
rect 4393 47846 4405 47898
rect 4405 47846 4435 47898
rect 4459 47846 4469 47898
rect 4469 47846 4515 47898
rect 4219 47844 4275 47846
rect 4299 47844 4355 47846
rect 4379 47844 4435 47846
rect 4459 47844 4515 47846
rect 4219 46810 4275 46812
rect 4299 46810 4355 46812
rect 4379 46810 4435 46812
rect 4459 46810 4515 46812
rect 4219 46758 4265 46810
rect 4265 46758 4275 46810
rect 4299 46758 4329 46810
rect 4329 46758 4341 46810
rect 4341 46758 4355 46810
rect 4379 46758 4393 46810
rect 4393 46758 4405 46810
rect 4405 46758 4435 46810
rect 4459 46758 4469 46810
rect 4469 46758 4515 46810
rect 4219 46756 4275 46758
rect 4299 46756 4355 46758
rect 4379 46756 4435 46758
rect 4459 46756 4515 46758
rect 4219 45722 4275 45724
rect 4299 45722 4355 45724
rect 4379 45722 4435 45724
rect 4459 45722 4515 45724
rect 4219 45670 4265 45722
rect 4265 45670 4275 45722
rect 4299 45670 4329 45722
rect 4329 45670 4341 45722
rect 4341 45670 4355 45722
rect 4379 45670 4393 45722
rect 4393 45670 4405 45722
rect 4405 45670 4435 45722
rect 4459 45670 4469 45722
rect 4469 45670 4515 45722
rect 4219 45668 4275 45670
rect 4299 45668 4355 45670
rect 4379 45668 4435 45670
rect 4459 45668 4515 45670
rect 4219 44634 4275 44636
rect 4299 44634 4355 44636
rect 4379 44634 4435 44636
rect 4459 44634 4515 44636
rect 4219 44582 4265 44634
rect 4265 44582 4275 44634
rect 4299 44582 4329 44634
rect 4329 44582 4341 44634
rect 4341 44582 4355 44634
rect 4379 44582 4393 44634
rect 4393 44582 4405 44634
rect 4405 44582 4435 44634
rect 4459 44582 4469 44634
rect 4469 44582 4515 44634
rect 4219 44580 4275 44582
rect 4299 44580 4355 44582
rect 4379 44580 4435 44582
rect 4459 44580 4515 44582
rect 4219 43546 4275 43548
rect 4299 43546 4355 43548
rect 4379 43546 4435 43548
rect 4459 43546 4515 43548
rect 4219 43494 4265 43546
rect 4265 43494 4275 43546
rect 4299 43494 4329 43546
rect 4329 43494 4341 43546
rect 4341 43494 4355 43546
rect 4379 43494 4393 43546
rect 4393 43494 4405 43546
rect 4405 43494 4435 43546
rect 4459 43494 4469 43546
rect 4469 43494 4515 43546
rect 4219 43492 4275 43494
rect 4299 43492 4355 43494
rect 4379 43492 4435 43494
rect 4459 43492 4515 43494
rect 4219 42458 4275 42460
rect 4299 42458 4355 42460
rect 4379 42458 4435 42460
rect 4459 42458 4515 42460
rect 4219 42406 4265 42458
rect 4265 42406 4275 42458
rect 4299 42406 4329 42458
rect 4329 42406 4341 42458
rect 4341 42406 4355 42458
rect 4379 42406 4393 42458
rect 4393 42406 4405 42458
rect 4405 42406 4435 42458
rect 4459 42406 4469 42458
rect 4469 42406 4515 42458
rect 4219 42404 4275 42406
rect 4299 42404 4355 42406
rect 4379 42404 4435 42406
rect 4459 42404 4515 42406
rect 4219 41370 4275 41372
rect 4299 41370 4355 41372
rect 4379 41370 4435 41372
rect 4459 41370 4515 41372
rect 4219 41318 4265 41370
rect 4265 41318 4275 41370
rect 4299 41318 4329 41370
rect 4329 41318 4341 41370
rect 4341 41318 4355 41370
rect 4379 41318 4393 41370
rect 4393 41318 4405 41370
rect 4405 41318 4435 41370
rect 4459 41318 4469 41370
rect 4469 41318 4515 41370
rect 4219 41316 4275 41318
rect 4299 41316 4355 41318
rect 4379 41316 4435 41318
rect 4459 41316 4515 41318
rect 4219 40282 4275 40284
rect 4299 40282 4355 40284
rect 4379 40282 4435 40284
rect 4459 40282 4515 40284
rect 4219 40230 4265 40282
rect 4265 40230 4275 40282
rect 4299 40230 4329 40282
rect 4329 40230 4341 40282
rect 4341 40230 4355 40282
rect 4379 40230 4393 40282
rect 4393 40230 4405 40282
rect 4405 40230 4435 40282
rect 4459 40230 4469 40282
rect 4469 40230 4515 40282
rect 4219 40228 4275 40230
rect 4299 40228 4355 40230
rect 4379 40228 4435 40230
rect 4459 40228 4515 40230
rect 4219 39194 4275 39196
rect 4299 39194 4355 39196
rect 4379 39194 4435 39196
rect 4459 39194 4515 39196
rect 4219 39142 4265 39194
rect 4265 39142 4275 39194
rect 4299 39142 4329 39194
rect 4329 39142 4341 39194
rect 4341 39142 4355 39194
rect 4379 39142 4393 39194
rect 4393 39142 4405 39194
rect 4405 39142 4435 39194
rect 4459 39142 4469 39194
rect 4469 39142 4515 39194
rect 4219 39140 4275 39142
rect 4299 39140 4355 39142
rect 4379 39140 4435 39142
rect 4459 39140 4515 39142
rect 4219 38106 4275 38108
rect 4299 38106 4355 38108
rect 4379 38106 4435 38108
rect 4459 38106 4515 38108
rect 4219 38054 4265 38106
rect 4265 38054 4275 38106
rect 4299 38054 4329 38106
rect 4329 38054 4341 38106
rect 4341 38054 4355 38106
rect 4379 38054 4393 38106
rect 4393 38054 4405 38106
rect 4405 38054 4435 38106
rect 4459 38054 4469 38106
rect 4469 38054 4515 38106
rect 4219 38052 4275 38054
rect 4299 38052 4355 38054
rect 4379 38052 4435 38054
rect 4459 38052 4515 38054
rect 4219 37018 4275 37020
rect 4299 37018 4355 37020
rect 4379 37018 4435 37020
rect 4459 37018 4515 37020
rect 4219 36966 4265 37018
rect 4265 36966 4275 37018
rect 4299 36966 4329 37018
rect 4329 36966 4341 37018
rect 4341 36966 4355 37018
rect 4379 36966 4393 37018
rect 4393 36966 4405 37018
rect 4405 36966 4435 37018
rect 4459 36966 4469 37018
rect 4469 36966 4515 37018
rect 4219 36964 4275 36966
rect 4299 36964 4355 36966
rect 4379 36964 4435 36966
rect 4459 36964 4515 36966
rect 4219 35930 4275 35932
rect 4299 35930 4355 35932
rect 4379 35930 4435 35932
rect 4459 35930 4515 35932
rect 4219 35878 4265 35930
rect 4265 35878 4275 35930
rect 4299 35878 4329 35930
rect 4329 35878 4341 35930
rect 4341 35878 4355 35930
rect 4379 35878 4393 35930
rect 4393 35878 4405 35930
rect 4405 35878 4435 35930
rect 4459 35878 4469 35930
rect 4469 35878 4515 35930
rect 4219 35876 4275 35878
rect 4299 35876 4355 35878
rect 4379 35876 4435 35878
rect 4459 35876 4515 35878
rect 4219 34842 4275 34844
rect 4299 34842 4355 34844
rect 4379 34842 4435 34844
rect 4459 34842 4515 34844
rect 4219 34790 4265 34842
rect 4265 34790 4275 34842
rect 4299 34790 4329 34842
rect 4329 34790 4341 34842
rect 4341 34790 4355 34842
rect 4379 34790 4393 34842
rect 4393 34790 4405 34842
rect 4405 34790 4435 34842
rect 4459 34790 4469 34842
rect 4469 34790 4515 34842
rect 4219 34788 4275 34790
rect 4299 34788 4355 34790
rect 4379 34788 4435 34790
rect 4459 34788 4515 34790
rect 4219 33754 4275 33756
rect 4299 33754 4355 33756
rect 4379 33754 4435 33756
rect 4459 33754 4515 33756
rect 4219 33702 4265 33754
rect 4265 33702 4275 33754
rect 4299 33702 4329 33754
rect 4329 33702 4341 33754
rect 4341 33702 4355 33754
rect 4379 33702 4393 33754
rect 4393 33702 4405 33754
rect 4405 33702 4435 33754
rect 4459 33702 4469 33754
rect 4469 33702 4515 33754
rect 4219 33700 4275 33702
rect 4299 33700 4355 33702
rect 4379 33700 4435 33702
rect 4459 33700 4515 33702
rect 4219 32666 4275 32668
rect 4299 32666 4355 32668
rect 4379 32666 4435 32668
rect 4459 32666 4515 32668
rect 4219 32614 4265 32666
rect 4265 32614 4275 32666
rect 4299 32614 4329 32666
rect 4329 32614 4341 32666
rect 4341 32614 4355 32666
rect 4379 32614 4393 32666
rect 4393 32614 4405 32666
rect 4405 32614 4435 32666
rect 4459 32614 4469 32666
rect 4469 32614 4515 32666
rect 4219 32612 4275 32614
rect 4299 32612 4355 32614
rect 4379 32612 4435 32614
rect 4459 32612 4515 32614
rect 4219 31578 4275 31580
rect 4299 31578 4355 31580
rect 4379 31578 4435 31580
rect 4459 31578 4515 31580
rect 4219 31526 4265 31578
rect 4265 31526 4275 31578
rect 4299 31526 4329 31578
rect 4329 31526 4341 31578
rect 4341 31526 4355 31578
rect 4379 31526 4393 31578
rect 4393 31526 4405 31578
rect 4405 31526 4435 31578
rect 4459 31526 4469 31578
rect 4469 31526 4515 31578
rect 4219 31524 4275 31526
rect 4299 31524 4355 31526
rect 4379 31524 4435 31526
rect 4459 31524 4515 31526
rect 4219 30490 4275 30492
rect 4299 30490 4355 30492
rect 4379 30490 4435 30492
rect 4459 30490 4515 30492
rect 4219 30438 4265 30490
rect 4265 30438 4275 30490
rect 4299 30438 4329 30490
rect 4329 30438 4341 30490
rect 4341 30438 4355 30490
rect 4379 30438 4393 30490
rect 4393 30438 4405 30490
rect 4405 30438 4435 30490
rect 4459 30438 4469 30490
rect 4469 30438 4515 30490
rect 4219 30436 4275 30438
rect 4299 30436 4355 30438
rect 4379 30436 4435 30438
rect 4459 30436 4515 30438
rect 4219 29402 4275 29404
rect 4299 29402 4355 29404
rect 4379 29402 4435 29404
rect 4459 29402 4515 29404
rect 4219 29350 4265 29402
rect 4265 29350 4275 29402
rect 4299 29350 4329 29402
rect 4329 29350 4341 29402
rect 4341 29350 4355 29402
rect 4379 29350 4393 29402
rect 4393 29350 4405 29402
rect 4405 29350 4435 29402
rect 4459 29350 4469 29402
rect 4469 29350 4515 29402
rect 4219 29348 4275 29350
rect 4299 29348 4355 29350
rect 4379 29348 4435 29350
rect 4459 29348 4515 29350
rect 4219 28314 4275 28316
rect 4299 28314 4355 28316
rect 4379 28314 4435 28316
rect 4459 28314 4515 28316
rect 4219 28262 4265 28314
rect 4265 28262 4275 28314
rect 4299 28262 4329 28314
rect 4329 28262 4341 28314
rect 4341 28262 4355 28314
rect 4379 28262 4393 28314
rect 4393 28262 4405 28314
rect 4405 28262 4435 28314
rect 4459 28262 4469 28314
rect 4469 28262 4515 28314
rect 4219 28260 4275 28262
rect 4299 28260 4355 28262
rect 4379 28260 4435 28262
rect 4459 28260 4515 28262
rect 4219 27226 4275 27228
rect 4299 27226 4355 27228
rect 4379 27226 4435 27228
rect 4459 27226 4515 27228
rect 4219 27174 4265 27226
rect 4265 27174 4275 27226
rect 4299 27174 4329 27226
rect 4329 27174 4341 27226
rect 4341 27174 4355 27226
rect 4379 27174 4393 27226
rect 4393 27174 4405 27226
rect 4405 27174 4435 27226
rect 4459 27174 4469 27226
rect 4469 27174 4515 27226
rect 4219 27172 4275 27174
rect 4299 27172 4355 27174
rect 4379 27172 4435 27174
rect 4459 27172 4515 27174
rect 4219 26138 4275 26140
rect 4299 26138 4355 26140
rect 4379 26138 4435 26140
rect 4459 26138 4515 26140
rect 4219 26086 4265 26138
rect 4265 26086 4275 26138
rect 4299 26086 4329 26138
rect 4329 26086 4341 26138
rect 4341 26086 4355 26138
rect 4379 26086 4393 26138
rect 4393 26086 4405 26138
rect 4405 26086 4435 26138
rect 4459 26086 4469 26138
rect 4469 26086 4515 26138
rect 4219 26084 4275 26086
rect 4299 26084 4355 26086
rect 4379 26084 4435 26086
rect 4459 26084 4515 26086
rect 4219 25050 4275 25052
rect 4299 25050 4355 25052
rect 4379 25050 4435 25052
rect 4459 25050 4515 25052
rect 4219 24998 4265 25050
rect 4265 24998 4275 25050
rect 4299 24998 4329 25050
rect 4329 24998 4341 25050
rect 4341 24998 4355 25050
rect 4379 24998 4393 25050
rect 4393 24998 4405 25050
rect 4405 24998 4435 25050
rect 4459 24998 4469 25050
rect 4469 24998 4515 25050
rect 4219 24996 4275 24998
rect 4299 24996 4355 24998
rect 4379 24996 4435 24998
rect 4459 24996 4515 24998
rect 4219 23962 4275 23964
rect 4299 23962 4355 23964
rect 4379 23962 4435 23964
rect 4459 23962 4515 23964
rect 4219 23910 4265 23962
rect 4265 23910 4275 23962
rect 4299 23910 4329 23962
rect 4329 23910 4341 23962
rect 4341 23910 4355 23962
rect 4379 23910 4393 23962
rect 4393 23910 4405 23962
rect 4405 23910 4435 23962
rect 4459 23910 4469 23962
rect 4469 23910 4515 23962
rect 4219 23908 4275 23910
rect 4299 23908 4355 23910
rect 4379 23908 4435 23910
rect 4459 23908 4515 23910
rect 4219 22874 4275 22876
rect 4299 22874 4355 22876
rect 4379 22874 4435 22876
rect 4459 22874 4515 22876
rect 4219 22822 4265 22874
rect 4265 22822 4275 22874
rect 4299 22822 4329 22874
rect 4329 22822 4341 22874
rect 4341 22822 4355 22874
rect 4379 22822 4393 22874
rect 4393 22822 4405 22874
rect 4405 22822 4435 22874
rect 4459 22822 4469 22874
rect 4469 22822 4515 22874
rect 4219 22820 4275 22822
rect 4299 22820 4355 22822
rect 4379 22820 4435 22822
rect 4459 22820 4515 22822
rect 4219 21786 4275 21788
rect 4299 21786 4355 21788
rect 4379 21786 4435 21788
rect 4459 21786 4515 21788
rect 4219 21734 4265 21786
rect 4265 21734 4275 21786
rect 4299 21734 4329 21786
rect 4329 21734 4341 21786
rect 4341 21734 4355 21786
rect 4379 21734 4393 21786
rect 4393 21734 4405 21786
rect 4405 21734 4435 21786
rect 4459 21734 4469 21786
rect 4469 21734 4515 21786
rect 4219 21732 4275 21734
rect 4299 21732 4355 21734
rect 4379 21732 4435 21734
rect 4459 21732 4515 21734
rect 4219 20698 4275 20700
rect 4299 20698 4355 20700
rect 4379 20698 4435 20700
rect 4459 20698 4515 20700
rect 4219 20646 4265 20698
rect 4265 20646 4275 20698
rect 4299 20646 4329 20698
rect 4329 20646 4341 20698
rect 4341 20646 4355 20698
rect 4379 20646 4393 20698
rect 4393 20646 4405 20698
rect 4405 20646 4435 20698
rect 4459 20646 4469 20698
rect 4469 20646 4515 20698
rect 4219 20644 4275 20646
rect 4299 20644 4355 20646
rect 4379 20644 4435 20646
rect 4459 20644 4515 20646
rect 4219 19610 4275 19612
rect 4299 19610 4355 19612
rect 4379 19610 4435 19612
rect 4459 19610 4515 19612
rect 4219 19558 4265 19610
rect 4265 19558 4275 19610
rect 4299 19558 4329 19610
rect 4329 19558 4341 19610
rect 4341 19558 4355 19610
rect 4379 19558 4393 19610
rect 4393 19558 4405 19610
rect 4405 19558 4435 19610
rect 4459 19558 4469 19610
rect 4469 19558 4515 19610
rect 4219 19556 4275 19558
rect 4299 19556 4355 19558
rect 4379 19556 4435 19558
rect 4459 19556 4515 19558
rect 4219 18522 4275 18524
rect 4299 18522 4355 18524
rect 4379 18522 4435 18524
rect 4459 18522 4515 18524
rect 4219 18470 4265 18522
rect 4265 18470 4275 18522
rect 4299 18470 4329 18522
rect 4329 18470 4341 18522
rect 4341 18470 4355 18522
rect 4379 18470 4393 18522
rect 4393 18470 4405 18522
rect 4405 18470 4435 18522
rect 4459 18470 4469 18522
rect 4469 18470 4515 18522
rect 4219 18468 4275 18470
rect 4299 18468 4355 18470
rect 4379 18468 4435 18470
rect 4459 18468 4515 18470
rect 4219 17434 4275 17436
rect 4299 17434 4355 17436
rect 4379 17434 4435 17436
rect 4459 17434 4515 17436
rect 4219 17382 4265 17434
rect 4265 17382 4275 17434
rect 4299 17382 4329 17434
rect 4329 17382 4341 17434
rect 4341 17382 4355 17434
rect 4379 17382 4393 17434
rect 4393 17382 4405 17434
rect 4405 17382 4435 17434
rect 4459 17382 4469 17434
rect 4469 17382 4515 17434
rect 4219 17380 4275 17382
rect 4299 17380 4355 17382
rect 4379 17380 4435 17382
rect 4459 17380 4515 17382
rect 2588 16890 2644 16892
rect 2668 16890 2724 16892
rect 2748 16890 2804 16892
rect 2828 16890 2884 16892
rect 2588 16838 2634 16890
rect 2634 16838 2644 16890
rect 2668 16838 2698 16890
rect 2698 16838 2710 16890
rect 2710 16838 2724 16890
rect 2748 16838 2762 16890
rect 2762 16838 2774 16890
rect 2774 16838 2804 16890
rect 2828 16838 2838 16890
rect 2838 16838 2884 16890
rect 2588 16836 2644 16838
rect 2668 16836 2724 16838
rect 2748 16836 2804 16838
rect 2828 16836 2884 16838
rect 4219 16346 4275 16348
rect 4299 16346 4355 16348
rect 4379 16346 4435 16348
rect 4459 16346 4515 16348
rect 4219 16294 4265 16346
rect 4265 16294 4275 16346
rect 4299 16294 4329 16346
rect 4329 16294 4341 16346
rect 4341 16294 4355 16346
rect 4379 16294 4393 16346
rect 4393 16294 4405 16346
rect 4405 16294 4435 16346
rect 4459 16294 4469 16346
rect 4469 16294 4515 16346
rect 4219 16292 4275 16294
rect 4299 16292 4355 16294
rect 4379 16292 4435 16294
rect 4459 16292 4515 16294
rect 2588 15802 2644 15804
rect 2668 15802 2724 15804
rect 2748 15802 2804 15804
rect 2828 15802 2884 15804
rect 2588 15750 2634 15802
rect 2634 15750 2644 15802
rect 2668 15750 2698 15802
rect 2698 15750 2710 15802
rect 2710 15750 2724 15802
rect 2748 15750 2762 15802
rect 2762 15750 2774 15802
rect 2774 15750 2804 15802
rect 2828 15750 2838 15802
rect 2838 15750 2884 15802
rect 2588 15748 2644 15750
rect 2668 15748 2724 15750
rect 2748 15748 2804 15750
rect 2828 15748 2884 15750
rect 4219 15258 4275 15260
rect 4299 15258 4355 15260
rect 4379 15258 4435 15260
rect 4459 15258 4515 15260
rect 4219 15206 4265 15258
rect 4265 15206 4275 15258
rect 4299 15206 4329 15258
rect 4329 15206 4341 15258
rect 4341 15206 4355 15258
rect 4379 15206 4393 15258
rect 4393 15206 4405 15258
rect 4405 15206 4435 15258
rect 4459 15206 4469 15258
rect 4469 15206 4515 15258
rect 4219 15204 4275 15206
rect 4299 15204 4355 15206
rect 4379 15204 4435 15206
rect 4459 15204 4515 15206
rect 2588 14714 2644 14716
rect 2668 14714 2724 14716
rect 2748 14714 2804 14716
rect 2828 14714 2884 14716
rect 2588 14662 2634 14714
rect 2634 14662 2644 14714
rect 2668 14662 2698 14714
rect 2698 14662 2710 14714
rect 2710 14662 2724 14714
rect 2748 14662 2762 14714
rect 2762 14662 2774 14714
rect 2774 14662 2804 14714
rect 2828 14662 2838 14714
rect 2838 14662 2884 14714
rect 2588 14660 2644 14662
rect 2668 14660 2724 14662
rect 2748 14660 2804 14662
rect 2828 14660 2884 14662
rect 4219 14170 4275 14172
rect 4299 14170 4355 14172
rect 4379 14170 4435 14172
rect 4459 14170 4515 14172
rect 4219 14118 4265 14170
rect 4265 14118 4275 14170
rect 4299 14118 4329 14170
rect 4329 14118 4341 14170
rect 4341 14118 4355 14170
rect 4379 14118 4393 14170
rect 4393 14118 4405 14170
rect 4405 14118 4435 14170
rect 4459 14118 4469 14170
rect 4469 14118 4515 14170
rect 4219 14116 4275 14118
rect 4299 14116 4355 14118
rect 4379 14116 4435 14118
rect 4459 14116 4515 14118
rect 2588 13626 2644 13628
rect 2668 13626 2724 13628
rect 2748 13626 2804 13628
rect 2828 13626 2884 13628
rect 2588 13574 2634 13626
rect 2634 13574 2644 13626
rect 2668 13574 2698 13626
rect 2698 13574 2710 13626
rect 2710 13574 2724 13626
rect 2748 13574 2762 13626
rect 2762 13574 2774 13626
rect 2774 13574 2804 13626
rect 2828 13574 2838 13626
rect 2838 13574 2884 13626
rect 2588 13572 2644 13574
rect 2668 13572 2724 13574
rect 2748 13572 2804 13574
rect 2828 13572 2884 13574
rect 4219 13082 4275 13084
rect 4299 13082 4355 13084
rect 4379 13082 4435 13084
rect 4459 13082 4515 13084
rect 4219 13030 4265 13082
rect 4265 13030 4275 13082
rect 4299 13030 4329 13082
rect 4329 13030 4341 13082
rect 4341 13030 4355 13082
rect 4379 13030 4393 13082
rect 4393 13030 4405 13082
rect 4405 13030 4435 13082
rect 4459 13030 4469 13082
rect 4469 13030 4515 13082
rect 4219 13028 4275 13030
rect 4299 13028 4355 13030
rect 4379 13028 4435 13030
rect 4459 13028 4515 13030
rect 2588 12538 2644 12540
rect 2668 12538 2724 12540
rect 2748 12538 2804 12540
rect 2828 12538 2884 12540
rect 2588 12486 2634 12538
rect 2634 12486 2644 12538
rect 2668 12486 2698 12538
rect 2698 12486 2710 12538
rect 2710 12486 2724 12538
rect 2748 12486 2762 12538
rect 2762 12486 2774 12538
rect 2774 12486 2804 12538
rect 2828 12486 2838 12538
rect 2838 12486 2884 12538
rect 2588 12484 2644 12486
rect 2668 12484 2724 12486
rect 2748 12484 2804 12486
rect 2828 12484 2884 12486
rect 4219 11994 4275 11996
rect 4299 11994 4355 11996
rect 4379 11994 4435 11996
rect 4459 11994 4515 11996
rect 4219 11942 4265 11994
rect 4265 11942 4275 11994
rect 4299 11942 4329 11994
rect 4329 11942 4341 11994
rect 4341 11942 4355 11994
rect 4379 11942 4393 11994
rect 4393 11942 4405 11994
rect 4405 11942 4435 11994
rect 4459 11942 4469 11994
rect 4469 11942 4515 11994
rect 4219 11940 4275 11942
rect 4299 11940 4355 11942
rect 4379 11940 4435 11942
rect 4459 11940 4515 11942
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 4219 10906 4275 10908
rect 4299 10906 4355 10908
rect 4379 10906 4435 10908
rect 4459 10906 4515 10908
rect 4219 10854 4265 10906
rect 4265 10854 4275 10906
rect 4299 10854 4329 10906
rect 4329 10854 4341 10906
rect 4341 10854 4355 10906
rect 4379 10854 4393 10906
rect 4393 10854 4405 10906
rect 4405 10854 4435 10906
rect 4459 10854 4469 10906
rect 4469 10854 4515 10906
rect 4219 10852 4275 10854
rect 4299 10852 4355 10854
rect 4379 10852 4435 10854
rect 4459 10852 4515 10854
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 5078 42608 5134 42664
rect 5078 40432 5134 40488
rect 4219 9818 4275 9820
rect 4299 9818 4355 9820
rect 4379 9818 4435 9820
rect 4459 9818 4515 9820
rect 4219 9766 4265 9818
rect 4265 9766 4275 9818
rect 4299 9766 4329 9818
rect 4329 9766 4341 9818
rect 4341 9766 4355 9818
rect 4379 9766 4393 9818
rect 4393 9766 4405 9818
rect 4405 9766 4435 9818
rect 4459 9766 4469 9818
rect 4469 9766 4515 9818
rect 4219 9764 4275 9766
rect 4299 9764 4355 9766
rect 4379 9764 4435 9766
rect 4459 9764 4515 9766
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 4219 8730 4275 8732
rect 4299 8730 4355 8732
rect 4379 8730 4435 8732
rect 4459 8730 4515 8732
rect 4219 8678 4265 8730
rect 4265 8678 4275 8730
rect 4299 8678 4329 8730
rect 4329 8678 4341 8730
rect 4341 8678 4355 8730
rect 4379 8678 4393 8730
rect 4393 8678 4405 8730
rect 4405 8678 4435 8730
rect 4459 8678 4469 8730
rect 4469 8678 4515 8730
rect 4219 8676 4275 8678
rect 4299 8676 4355 8678
rect 4379 8676 4435 8678
rect 4459 8676 4515 8678
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 4219 7642 4275 7644
rect 4299 7642 4355 7644
rect 4379 7642 4435 7644
rect 4459 7642 4515 7644
rect 4219 7590 4265 7642
rect 4265 7590 4275 7642
rect 4299 7590 4329 7642
rect 4329 7590 4341 7642
rect 4341 7590 4355 7642
rect 4379 7590 4393 7642
rect 4393 7590 4405 7642
rect 4405 7590 4435 7642
rect 4459 7590 4469 7642
rect 4469 7590 4515 7642
rect 4219 7588 4275 7590
rect 4299 7588 4355 7590
rect 4379 7588 4435 7590
rect 4459 7588 4515 7590
rect 5851 71290 5907 71292
rect 5931 71290 5987 71292
rect 6011 71290 6067 71292
rect 6091 71290 6147 71292
rect 5851 71238 5897 71290
rect 5897 71238 5907 71290
rect 5931 71238 5961 71290
rect 5961 71238 5973 71290
rect 5973 71238 5987 71290
rect 6011 71238 6025 71290
rect 6025 71238 6037 71290
rect 6037 71238 6067 71290
rect 6091 71238 6101 71290
rect 6101 71238 6147 71290
rect 5851 71236 5907 71238
rect 5931 71236 5987 71238
rect 6011 71236 6067 71238
rect 6091 71236 6147 71238
rect 7483 74010 7539 74012
rect 7563 74010 7619 74012
rect 7643 74010 7699 74012
rect 7723 74010 7779 74012
rect 7483 73958 7529 74010
rect 7529 73958 7539 74010
rect 7563 73958 7593 74010
rect 7593 73958 7605 74010
rect 7605 73958 7619 74010
rect 7643 73958 7657 74010
rect 7657 73958 7669 74010
rect 7669 73958 7699 74010
rect 7723 73958 7733 74010
rect 7733 73958 7779 74010
rect 7483 73956 7539 73958
rect 7563 73956 7619 73958
rect 7643 73956 7699 73958
rect 7723 73956 7779 73958
rect 5851 70202 5907 70204
rect 5931 70202 5987 70204
rect 6011 70202 6067 70204
rect 6091 70202 6147 70204
rect 5851 70150 5897 70202
rect 5897 70150 5907 70202
rect 5931 70150 5961 70202
rect 5961 70150 5973 70202
rect 5973 70150 5987 70202
rect 6011 70150 6025 70202
rect 6025 70150 6037 70202
rect 6037 70150 6067 70202
rect 6091 70150 6101 70202
rect 6101 70150 6147 70202
rect 5851 70148 5907 70150
rect 5931 70148 5987 70150
rect 6011 70148 6067 70150
rect 6091 70148 6147 70150
rect 5851 69114 5907 69116
rect 5931 69114 5987 69116
rect 6011 69114 6067 69116
rect 6091 69114 6147 69116
rect 5851 69062 5897 69114
rect 5897 69062 5907 69114
rect 5931 69062 5961 69114
rect 5961 69062 5973 69114
rect 5973 69062 5987 69114
rect 6011 69062 6025 69114
rect 6025 69062 6037 69114
rect 6037 69062 6067 69114
rect 6091 69062 6101 69114
rect 6101 69062 6147 69114
rect 5851 69060 5907 69062
rect 5931 69060 5987 69062
rect 6011 69060 6067 69062
rect 6091 69060 6147 69062
rect 5851 68026 5907 68028
rect 5931 68026 5987 68028
rect 6011 68026 6067 68028
rect 6091 68026 6147 68028
rect 5851 67974 5897 68026
rect 5897 67974 5907 68026
rect 5931 67974 5961 68026
rect 5961 67974 5973 68026
rect 5973 67974 5987 68026
rect 6011 67974 6025 68026
rect 6025 67974 6037 68026
rect 6037 67974 6067 68026
rect 6091 67974 6101 68026
rect 6101 67974 6147 68026
rect 5851 67972 5907 67974
rect 5931 67972 5987 67974
rect 6011 67972 6067 67974
rect 6091 67972 6147 67974
rect 5851 66938 5907 66940
rect 5931 66938 5987 66940
rect 6011 66938 6067 66940
rect 6091 66938 6147 66940
rect 5851 66886 5897 66938
rect 5897 66886 5907 66938
rect 5931 66886 5961 66938
rect 5961 66886 5973 66938
rect 5973 66886 5987 66938
rect 6011 66886 6025 66938
rect 6025 66886 6037 66938
rect 6037 66886 6067 66938
rect 6091 66886 6101 66938
rect 6101 66886 6147 66938
rect 5851 66884 5907 66886
rect 5931 66884 5987 66886
rect 6011 66884 6067 66886
rect 6091 66884 6147 66886
rect 5851 65850 5907 65852
rect 5931 65850 5987 65852
rect 6011 65850 6067 65852
rect 6091 65850 6147 65852
rect 5851 65798 5897 65850
rect 5897 65798 5907 65850
rect 5931 65798 5961 65850
rect 5961 65798 5973 65850
rect 5973 65798 5987 65850
rect 6011 65798 6025 65850
rect 6025 65798 6037 65850
rect 6037 65798 6067 65850
rect 6091 65798 6101 65850
rect 6101 65798 6147 65850
rect 5851 65796 5907 65798
rect 5931 65796 5987 65798
rect 6011 65796 6067 65798
rect 6091 65796 6147 65798
rect 5851 64762 5907 64764
rect 5931 64762 5987 64764
rect 6011 64762 6067 64764
rect 6091 64762 6147 64764
rect 5851 64710 5897 64762
rect 5897 64710 5907 64762
rect 5931 64710 5961 64762
rect 5961 64710 5973 64762
rect 5973 64710 5987 64762
rect 6011 64710 6025 64762
rect 6025 64710 6037 64762
rect 6037 64710 6067 64762
rect 6091 64710 6101 64762
rect 6101 64710 6147 64762
rect 5851 64708 5907 64710
rect 5931 64708 5987 64710
rect 6011 64708 6067 64710
rect 6091 64708 6147 64710
rect 5851 63674 5907 63676
rect 5931 63674 5987 63676
rect 6011 63674 6067 63676
rect 6091 63674 6147 63676
rect 5851 63622 5897 63674
rect 5897 63622 5907 63674
rect 5931 63622 5961 63674
rect 5961 63622 5973 63674
rect 5973 63622 5987 63674
rect 6011 63622 6025 63674
rect 6025 63622 6037 63674
rect 6037 63622 6067 63674
rect 6091 63622 6101 63674
rect 6101 63622 6147 63674
rect 5851 63620 5907 63622
rect 5931 63620 5987 63622
rect 6011 63620 6067 63622
rect 6091 63620 6147 63622
rect 5851 62586 5907 62588
rect 5931 62586 5987 62588
rect 6011 62586 6067 62588
rect 6091 62586 6147 62588
rect 5851 62534 5897 62586
rect 5897 62534 5907 62586
rect 5931 62534 5961 62586
rect 5961 62534 5973 62586
rect 5973 62534 5987 62586
rect 6011 62534 6025 62586
rect 6025 62534 6037 62586
rect 6037 62534 6067 62586
rect 6091 62534 6101 62586
rect 6101 62534 6147 62586
rect 5851 62532 5907 62534
rect 5931 62532 5987 62534
rect 6011 62532 6067 62534
rect 6091 62532 6147 62534
rect 5851 61498 5907 61500
rect 5931 61498 5987 61500
rect 6011 61498 6067 61500
rect 6091 61498 6147 61500
rect 5851 61446 5897 61498
rect 5897 61446 5907 61498
rect 5931 61446 5961 61498
rect 5961 61446 5973 61498
rect 5973 61446 5987 61498
rect 6011 61446 6025 61498
rect 6025 61446 6037 61498
rect 6037 61446 6067 61498
rect 6091 61446 6101 61498
rect 6101 61446 6147 61498
rect 5851 61444 5907 61446
rect 5931 61444 5987 61446
rect 6011 61444 6067 61446
rect 6091 61444 6147 61446
rect 5851 60410 5907 60412
rect 5931 60410 5987 60412
rect 6011 60410 6067 60412
rect 6091 60410 6147 60412
rect 5851 60358 5897 60410
rect 5897 60358 5907 60410
rect 5931 60358 5961 60410
rect 5961 60358 5973 60410
rect 5973 60358 5987 60410
rect 6011 60358 6025 60410
rect 6025 60358 6037 60410
rect 6037 60358 6067 60410
rect 6091 60358 6101 60410
rect 6101 60358 6147 60410
rect 5851 60356 5907 60358
rect 5931 60356 5987 60358
rect 6011 60356 6067 60358
rect 6091 60356 6147 60358
rect 5851 59322 5907 59324
rect 5931 59322 5987 59324
rect 6011 59322 6067 59324
rect 6091 59322 6147 59324
rect 5851 59270 5897 59322
rect 5897 59270 5907 59322
rect 5931 59270 5961 59322
rect 5961 59270 5973 59322
rect 5973 59270 5987 59322
rect 6011 59270 6025 59322
rect 6025 59270 6037 59322
rect 6037 59270 6067 59322
rect 6091 59270 6101 59322
rect 6101 59270 6147 59322
rect 5851 59268 5907 59270
rect 5931 59268 5987 59270
rect 6011 59268 6067 59270
rect 6091 59268 6147 59270
rect 5851 58234 5907 58236
rect 5931 58234 5987 58236
rect 6011 58234 6067 58236
rect 6091 58234 6147 58236
rect 5851 58182 5897 58234
rect 5897 58182 5907 58234
rect 5931 58182 5961 58234
rect 5961 58182 5973 58234
rect 5973 58182 5987 58234
rect 6011 58182 6025 58234
rect 6025 58182 6037 58234
rect 6037 58182 6067 58234
rect 6091 58182 6101 58234
rect 6101 58182 6147 58234
rect 5851 58180 5907 58182
rect 5931 58180 5987 58182
rect 6011 58180 6067 58182
rect 6091 58180 6147 58182
rect 5851 57146 5907 57148
rect 5931 57146 5987 57148
rect 6011 57146 6067 57148
rect 6091 57146 6147 57148
rect 5851 57094 5897 57146
rect 5897 57094 5907 57146
rect 5931 57094 5961 57146
rect 5961 57094 5973 57146
rect 5973 57094 5987 57146
rect 6011 57094 6025 57146
rect 6025 57094 6037 57146
rect 6037 57094 6067 57146
rect 6091 57094 6101 57146
rect 6101 57094 6147 57146
rect 5851 57092 5907 57094
rect 5931 57092 5987 57094
rect 6011 57092 6067 57094
rect 6091 57092 6147 57094
rect 5851 56058 5907 56060
rect 5931 56058 5987 56060
rect 6011 56058 6067 56060
rect 6091 56058 6147 56060
rect 5851 56006 5897 56058
rect 5897 56006 5907 56058
rect 5931 56006 5961 56058
rect 5961 56006 5973 56058
rect 5973 56006 5987 56058
rect 6011 56006 6025 56058
rect 6025 56006 6037 56058
rect 6037 56006 6067 56058
rect 6091 56006 6101 56058
rect 6101 56006 6147 56058
rect 5851 56004 5907 56006
rect 5931 56004 5987 56006
rect 6011 56004 6067 56006
rect 6091 56004 6147 56006
rect 5851 54970 5907 54972
rect 5931 54970 5987 54972
rect 6011 54970 6067 54972
rect 6091 54970 6147 54972
rect 5851 54918 5897 54970
rect 5897 54918 5907 54970
rect 5931 54918 5961 54970
rect 5961 54918 5973 54970
rect 5973 54918 5987 54970
rect 6011 54918 6025 54970
rect 6025 54918 6037 54970
rect 6037 54918 6067 54970
rect 6091 54918 6101 54970
rect 6101 54918 6147 54970
rect 5851 54916 5907 54918
rect 5931 54916 5987 54918
rect 6011 54916 6067 54918
rect 6091 54916 6147 54918
rect 5851 53882 5907 53884
rect 5931 53882 5987 53884
rect 6011 53882 6067 53884
rect 6091 53882 6147 53884
rect 5851 53830 5897 53882
rect 5897 53830 5907 53882
rect 5931 53830 5961 53882
rect 5961 53830 5973 53882
rect 5973 53830 5987 53882
rect 6011 53830 6025 53882
rect 6025 53830 6037 53882
rect 6037 53830 6067 53882
rect 6091 53830 6101 53882
rect 6101 53830 6147 53882
rect 5851 53828 5907 53830
rect 5931 53828 5987 53830
rect 6011 53828 6067 53830
rect 6091 53828 6147 53830
rect 5851 52794 5907 52796
rect 5931 52794 5987 52796
rect 6011 52794 6067 52796
rect 6091 52794 6147 52796
rect 5851 52742 5897 52794
rect 5897 52742 5907 52794
rect 5931 52742 5961 52794
rect 5961 52742 5973 52794
rect 5973 52742 5987 52794
rect 6011 52742 6025 52794
rect 6025 52742 6037 52794
rect 6037 52742 6067 52794
rect 6091 52742 6101 52794
rect 6101 52742 6147 52794
rect 5851 52740 5907 52742
rect 5931 52740 5987 52742
rect 6011 52740 6067 52742
rect 6091 52740 6147 52742
rect 5851 51706 5907 51708
rect 5931 51706 5987 51708
rect 6011 51706 6067 51708
rect 6091 51706 6147 51708
rect 5851 51654 5897 51706
rect 5897 51654 5907 51706
rect 5931 51654 5961 51706
rect 5961 51654 5973 51706
rect 5973 51654 5987 51706
rect 6011 51654 6025 51706
rect 6025 51654 6037 51706
rect 6037 51654 6067 51706
rect 6091 51654 6101 51706
rect 6101 51654 6147 51706
rect 5851 51652 5907 51654
rect 5931 51652 5987 51654
rect 6011 51652 6067 51654
rect 6091 51652 6147 51654
rect 5851 50618 5907 50620
rect 5931 50618 5987 50620
rect 6011 50618 6067 50620
rect 6091 50618 6147 50620
rect 5851 50566 5897 50618
rect 5897 50566 5907 50618
rect 5931 50566 5961 50618
rect 5961 50566 5973 50618
rect 5973 50566 5987 50618
rect 6011 50566 6025 50618
rect 6025 50566 6037 50618
rect 6037 50566 6067 50618
rect 6091 50566 6101 50618
rect 6101 50566 6147 50618
rect 5851 50564 5907 50566
rect 5931 50564 5987 50566
rect 6011 50564 6067 50566
rect 6091 50564 6147 50566
rect 5851 49530 5907 49532
rect 5931 49530 5987 49532
rect 6011 49530 6067 49532
rect 6091 49530 6147 49532
rect 5851 49478 5897 49530
rect 5897 49478 5907 49530
rect 5931 49478 5961 49530
rect 5961 49478 5973 49530
rect 5973 49478 5987 49530
rect 6011 49478 6025 49530
rect 6025 49478 6037 49530
rect 6037 49478 6067 49530
rect 6091 49478 6101 49530
rect 6101 49478 6147 49530
rect 5851 49476 5907 49478
rect 5931 49476 5987 49478
rect 6011 49476 6067 49478
rect 6091 49476 6147 49478
rect 5851 48442 5907 48444
rect 5931 48442 5987 48444
rect 6011 48442 6067 48444
rect 6091 48442 6147 48444
rect 5851 48390 5897 48442
rect 5897 48390 5907 48442
rect 5931 48390 5961 48442
rect 5961 48390 5973 48442
rect 5973 48390 5987 48442
rect 6011 48390 6025 48442
rect 6025 48390 6037 48442
rect 6037 48390 6067 48442
rect 6091 48390 6101 48442
rect 6101 48390 6147 48442
rect 5851 48388 5907 48390
rect 5931 48388 5987 48390
rect 6011 48388 6067 48390
rect 6091 48388 6147 48390
rect 5851 47354 5907 47356
rect 5931 47354 5987 47356
rect 6011 47354 6067 47356
rect 6091 47354 6147 47356
rect 5851 47302 5897 47354
rect 5897 47302 5907 47354
rect 5931 47302 5961 47354
rect 5961 47302 5973 47354
rect 5973 47302 5987 47354
rect 6011 47302 6025 47354
rect 6025 47302 6037 47354
rect 6037 47302 6067 47354
rect 6091 47302 6101 47354
rect 6101 47302 6147 47354
rect 5851 47300 5907 47302
rect 5931 47300 5987 47302
rect 6011 47300 6067 47302
rect 6091 47300 6147 47302
rect 5354 13388 5410 13424
rect 5354 13368 5356 13388
rect 5356 13368 5408 13388
rect 5408 13368 5410 13388
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 4219 6554 4275 6556
rect 4299 6554 4355 6556
rect 4379 6554 4435 6556
rect 4459 6554 4515 6556
rect 4219 6502 4265 6554
rect 4265 6502 4275 6554
rect 4299 6502 4329 6554
rect 4329 6502 4341 6554
rect 4341 6502 4355 6554
rect 4379 6502 4393 6554
rect 4393 6502 4405 6554
rect 4405 6502 4435 6554
rect 4459 6502 4469 6554
rect 4469 6502 4515 6554
rect 4219 6500 4275 6502
rect 4299 6500 4355 6502
rect 4379 6500 4435 6502
rect 4459 6500 4515 6502
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 5851 46266 5907 46268
rect 5931 46266 5987 46268
rect 6011 46266 6067 46268
rect 6091 46266 6147 46268
rect 5851 46214 5897 46266
rect 5897 46214 5907 46266
rect 5931 46214 5961 46266
rect 5961 46214 5973 46266
rect 5973 46214 5987 46266
rect 6011 46214 6025 46266
rect 6025 46214 6037 46266
rect 6037 46214 6067 46266
rect 6091 46214 6101 46266
rect 6101 46214 6147 46266
rect 5851 46212 5907 46214
rect 5931 46212 5987 46214
rect 6011 46212 6067 46214
rect 6091 46212 6147 46214
rect 5851 45178 5907 45180
rect 5931 45178 5987 45180
rect 6011 45178 6067 45180
rect 6091 45178 6147 45180
rect 5851 45126 5897 45178
rect 5897 45126 5907 45178
rect 5931 45126 5961 45178
rect 5961 45126 5973 45178
rect 5973 45126 5987 45178
rect 6011 45126 6025 45178
rect 6025 45126 6037 45178
rect 6037 45126 6067 45178
rect 6091 45126 6101 45178
rect 6101 45126 6147 45178
rect 5851 45124 5907 45126
rect 5931 45124 5987 45126
rect 6011 45124 6067 45126
rect 6091 45124 6147 45126
rect 5851 44090 5907 44092
rect 5931 44090 5987 44092
rect 6011 44090 6067 44092
rect 6091 44090 6147 44092
rect 5851 44038 5897 44090
rect 5897 44038 5907 44090
rect 5931 44038 5961 44090
rect 5961 44038 5973 44090
rect 5973 44038 5987 44090
rect 6011 44038 6025 44090
rect 6025 44038 6037 44090
rect 6037 44038 6067 44090
rect 6091 44038 6101 44090
rect 6101 44038 6147 44090
rect 5851 44036 5907 44038
rect 5931 44036 5987 44038
rect 6011 44036 6067 44038
rect 6091 44036 6147 44038
rect 5851 43002 5907 43004
rect 5931 43002 5987 43004
rect 6011 43002 6067 43004
rect 6091 43002 6147 43004
rect 5851 42950 5897 43002
rect 5897 42950 5907 43002
rect 5931 42950 5961 43002
rect 5961 42950 5973 43002
rect 5973 42950 5987 43002
rect 6011 42950 6025 43002
rect 6025 42950 6037 43002
rect 6037 42950 6067 43002
rect 6091 42950 6101 43002
rect 6101 42950 6147 43002
rect 5851 42948 5907 42950
rect 5931 42948 5987 42950
rect 6011 42948 6067 42950
rect 6091 42948 6147 42950
rect 6090 42608 6146 42664
rect 5851 41914 5907 41916
rect 5931 41914 5987 41916
rect 6011 41914 6067 41916
rect 6091 41914 6147 41916
rect 5851 41862 5897 41914
rect 5897 41862 5907 41914
rect 5931 41862 5961 41914
rect 5961 41862 5973 41914
rect 5973 41862 5987 41914
rect 6011 41862 6025 41914
rect 6025 41862 6037 41914
rect 6037 41862 6067 41914
rect 6091 41862 6101 41914
rect 6101 41862 6147 41914
rect 5851 41860 5907 41862
rect 5931 41860 5987 41862
rect 6011 41860 6067 41862
rect 6091 41860 6147 41862
rect 5851 40826 5907 40828
rect 5931 40826 5987 40828
rect 6011 40826 6067 40828
rect 6091 40826 6147 40828
rect 5851 40774 5897 40826
rect 5897 40774 5907 40826
rect 5931 40774 5961 40826
rect 5961 40774 5973 40826
rect 5973 40774 5987 40826
rect 6011 40774 6025 40826
rect 6025 40774 6037 40826
rect 6037 40774 6067 40826
rect 6091 40774 6101 40826
rect 6101 40774 6147 40826
rect 5851 40772 5907 40774
rect 5931 40772 5987 40774
rect 6011 40772 6067 40774
rect 6091 40772 6147 40774
rect 5851 39738 5907 39740
rect 5931 39738 5987 39740
rect 6011 39738 6067 39740
rect 6091 39738 6147 39740
rect 5851 39686 5897 39738
rect 5897 39686 5907 39738
rect 5931 39686 5961 39738
rect 5961 39686 5973 39738
rect 5973 39686 5987 39738
rect 6011 39686 6025 39738
rect 6025 39686 6037 39738
rect 6037 39686 6067 39738
rect 6091 39686 6101 39738
rect 6101 39686 6147 39738
rect 5851 39684 5907 39686
rect 5931 39684 5987 39686
rect 6011 39684 6067 39686
rect 6091 39684 6147 39686
rect 5851 38650 5907 38652
rect 5931 38650 5987 38652
rect 6011 38650 6067 38652
rect 6091 38650 6147 38652
rect 5851 38598 5897 38650
rect 5897 38598 5907 38650
rect 5931 38598 5961 38650
rect 5961 38598 5973 38650
rect 5973 38598 5987 38650
rect 6011 38598 6025 38650
rect 6025 38598 6037 38650
rect 6037 38598 6067 38650
rect 6091 38598 6101 38650
rect 6101 38598 6147 38650
rect 5851 38596 5907 38598
rect 5931 38596 5987 38598
rect 6011 38596 6067 38598
rect 6091 38596 6147 38598
rect 5851 37562 5907 37564
rect 5931 37562 5987 37564
rect 6011 37562 6067 37564
rect 6091 37562 6147 37564
rect 5851 37510 5897 37562
rect 5897 37510 5907 37562
rect 5931 37510 5961 37562
rect 5961 37510 5973 37562
rect 5973 37510 5987 37562
rect 6011 37510 6025 37562
rect 6025 37510 6037 37562
rect 6037 37510 6067 37562
rect 6091 37510 6101 37562
rect 6101 37510 6147 37562
rect 5851 37508 5907 37510
rect 5931 37508 5987 37510
rect 6011 37508 6067 37510
rect 6091 37508 6147 37510
rect 5851 36474 5907 36476
rect 5931 36474 5987 36476
rect 6011 36474 6067 36476
rect 6091 36474 6147 36476
rect 5851 36422 5897 36474
rect 5897 36422 5907 36474
rect 5931 36422 5961 36474
rect 5961 36422 5973 36474
rect 5973 36422 5987 36474
rect 6011 36422 6025 36474
rect 6025 36422 6037 36474
rect 6037 36422 6067 36474
rect 6091 36422 6101 36474
rect 6101 36422 6147 36474
rect 5851 36420 5907 36422
rect 5931 36420 5987 36422
rect 6011 36420 6067 36422
rect 6091 36420 6147 36422
rect 5851 35386 5907 35388
rect 5931 35386 5987 35388
rect 6011 35386 6067 35388
rect 6091 35386 6147 35388
rect 5851 35334 5897 35386
rect 5897 35334 5907 35386
rect 5931 35334 5961 35386
rect 5961 35334 5973 35386
rect 5973 35334 5987 35386
rect 6011 35334 6025 35386
rect 6025 35334 6037 35386
rect 6037 35334 6067 35386
rect 6091 35334 6101 35386
rect 6101 35334 6147 35386
rect 5851 35332 5907 35334
rect 5931 35332 5987 35334
rect 6011 35332 6067 35334
rect 6091 35332 6147 35334
rect 5851 34298 5907 34300
rect 5931 34298 5987 34300
rect 6011 34298 6067 34300
rect 6091 34298 6147 34300
rect 5851 34246 5897 34298
rect 5897 34246 5907 34298
rect 5931 34246 5961 34298
rect 5961 34246 5973 34298
rect 5973 34246 5987 34298
rect 6011 34246 6025 34298
rect 6025 34246 6037 34298
rect 6037 34246 6067 34298
rect 6091 34246 6101 34298
rect 6101 34246 6147 34298
rect 5851 34244 5907 34246
rect 5931 34244 5987 34246
rect 6011 34244 6067 34246
rect 6091 34244 6147 34246
rect 5851 33210 5907 33212
rect 5931 33210 5987 33212
rect 6011 33210 6067 33212
rect 6091 33210 6147 33212
rect 5851 33158 5897 33210
rect 5897 33158 5907 33210
rect 5931 33158 5961 33210
rect 5961 33158 5973 33210
rect 5973 33158 5987 33210
rect 6011 33158 6025 33210
rect 6025 33158 6037 33210
rect 6037 33158 6067 33210
rect 6091 33158 6101 33210
rect 6101 33158 6147 33210
rect 5851 33156 5907 33158
rect 5931 33156 5987 33158
rect 6011 33156 6067 33158
rect 6091 33156 6147 33158
rect 5851 32122 5907 32124
rect 5931 32122 5987 32124
rect 6011 32122 6067 32124
rect 6091 32122 6147 32124
rect 5851 32070 5897 32122
rect 5897 32070 5907 32122
rect 5931 32070 5961 32122
rect 5961 32070 5973 32122
rect 5973 32070 5987 32122
rect 6011 32070 6025 32122
rect 6025 32070 6037 32122
rect 6037 32070 6067 32122
rect 6091 32070 6101 32122
rect 6101 32070 6147 32122
rect 5851 32068 5907 32070
rect 5931 32068 5987 32070
rect 6011 32068 6067 32070
rect 6091 32068 6147 32070
rect 6642 43016 6698 43072
rect 6550 39072 6606 39128
rect 5851 31034 5907 31036
rect 5931 31034 5987 31036
rect 6011 31034 6067 31036
rect 6091 31034 6147 31036
rect 5851 30982 5897 31034
rect 5897 30982 5907 31034
rect 5931 30982 5961 31034
rect 5961 30982 5973 31034
rect 5973 30982 5987 31034
rect 6011 30982 6025 31034
rect 6025 30982 6037 31034
rect 6037 30982 6067 31034
rect 6091 30982 6101 31034
rect 6101 30982 6147 31034
rect 5851 30980 5907 30982
rect 5931 30980 5987 30982
rect 6011 30980 6067 30982
rect 6091 30980 6147 30982
rect 5851 29946 5907 29948
rect 5931 29946 5987 29948
rect 6011 29946 6067 29948
rect 6091 29946 6147 29948
rect 5851 29894 5897 29946
rect 5897 29894 5907 29946
rect 5931 29894 5961 29946
rect 5961 29894 5973 29946
rect 5973 29894 5987 29946
rect 6011 29894 6025 29946
rect 6025 29894 6037 29946
rect 6037 29894 6067 29946
rect 6091 29894 6101 29946
rect 6101 29894 6147 29946
rect 5851 29892 5907 29894
rect 5931 29892 5987 29894
rect 6011 29892 6067 29894
rect 6091 29892 6147 29894
rect 5851 28858 5907 28860
rect 5931 28858 5987 28860
rect 6011 28858 6067 28860
rect 6091 28858 6147 28860
rect 5851 28806 5897 28858
rect 5897 28806 5907 28858
rect 5931 28806 5961 28858
rect 5961 28806 5973 28858
rect 5973 28806 5987 28858
rect 6011 28806 6025 28858
rect 6025 28806 6037 28858
rect 6037 28806 6067 28858
rect 6091 28806 6101 28858
rect 6101 28806 6147 28858
rect 5851 28804 5907 28806
rect 5931 28804 5987 28806
rect 6011 28804 6067 28806
rect 6091 28804 6147 28806
rect 5851 27770 5907 27772
rect 5931 27770 5987 27772
rect 6011 27770 6067 27772
rect 6091 27770 6147 27772
rect 5851 27718 5897 27770
rect 5897 27718 5907 27770
rect 5931 27718 5961 27770
rect 5961 27718 5973 27770
rect 5973 27718 5987 27770
rect 6011 27718 6025 27770
rect 6025 27718 6037 27770
rect 6037 27718 6067 27770
rect 6091 27718 6101 27770
rect 6101 27718 6147 27770
rect 5851 27716 5907 27718
rect 5931 27716 5987 27718
rect 6011 27716 6067 27718
rect 6091 27716 6147 27718
rect 5851 26682 5907 26684
rect 5931 26682 5987 26684
rect 6011 26682 6067 26684
rect 6091 26682 6147 26684
rect 5851 26630 5897 26682
rect 5897 26630 5907 26682
rect 5931 26630 5961 26682
rect 5961 26630 5973 26682
rect 5973 26630 5987 26682
rect 6011 26630 6025 26682
rect 6025 26630 6037 26682
rect 6037 26630 6067 26682
rect 6091 26630 6101 26682
rect 6101 26630 6147 26682
rect 5851 26628 5907 26630
rect 5931 26628 5987 26630
rect 6011 26628 6067 26630
rect 6091 26628 6147 26630
rect 5851 25594 5907 25596
rect 5931 25594 5987 25596
rect 6011 25594 6067 25596
rect 6091 25594 6147 25596
rect 5851 25542 5897 25594
rect 5897 25542 5907 25594
rect 5931 25542 5961 25594
rect 5961 25542 5973 25594
rect 5973 25542 5987 25594
rect 6011 25542 6025 25594
rect 6025 25542 6037 25594
rect 6037 25542 6067 25594
rect 6091 25542 6101 25594
rect 6101 25542 6147 25594
rect 5851 25540 5907 25542
rect 5931 25540 5987 25542
rect 6011 25540 6067 25542
rect 6091 25540 6147 25542
rect 5851 24506 5907 24508
rect 5931 24506 5987 24508
rect 6011 24506 6067 24508
rect 6091 24506 6147 24508
rect 5851 24454 5897 24506
rect 5897 24454 5907 24506
rect 5931 24454 5961 24506
rect 5961 24454 5973 24506
rect 5973 24454 5987 24506
rect 6011 24454 6025 24506
rect 6025 24454 6037 24506
rect 6037 24454 6067 24506
rect 6091 24454 6101 24506
rect 6101 24454 6147 24506
rect 5851 24452 5907 24454
rect 5931 24452 5987 24454
rect 6011 24452 6067 24454
rect 6091 24452 6147 24454
rect 5851 23418 5907 23420
rect 5931 23418 5987 23420
rect 6011 23418 6067 23420
rect 6091 23418 6147 23420
rect 5851 23366 5897 23418
rect 5897 23366 5907 23418
rect 5931 23366 5961 23418
rect 5961 23366 5973 23418
rect 5973 23366 5987 23418
rect 6011 23366 6025 23418
rect 6025 23366 6037 23418
rect 6037 23366 6067 23418
rect 6091 23366 6101 23418
rect 6101 23366 6147 23418
rect 5851 23364 5907 23366
rect 5931 23364 5987 23366
rect 6011 23364 6067 23366
rect 6091 23364 6147 23366
rect 5851 22330 5907 22332
rect 5931 22330 5987 22332
rect 6011 22330 6067 22332
rect 6091 22330 6147 22332
rect 5851 22278 5897 22330
rect 5897 22278 5907 22330
rect 5931 22278 5961 22330
rect 5961 22278 5973 22330
rect 5973 22278 5987 22330
rect 6011 22278 6025 22330
rect 6025 22278 6037 22330
rect 6037 22278 6067 22330
rect 6091 22278 6101 22330
rect 6101 22278 6147 22330
rect 5851 22276 5907 22278
rect 5931 22276 5987 22278
rect 6011 22276 6067 22278
rect 6091 22276 6147 22278
rect 5851 21242 5907 21244
rect 5931 21242 5987 21244
rect 6011 21242 6067 21244
rect 6091 21242 6147 21244
rect 5851 21190 5897 21242
rect 5897 21190 5907 21242
rect 5931 21190 5961 21242
rect 5961 21190 5973 21242
rect 5973 21190 5987 21242
rect 6011 21190 6025 21242
rect 6025 21190 6037 21242
rect 6037 21190 6067 21242
rect 6091 21190 6101 21242
rect 6101 21190 6147 21242
rect 5851 21188 5907 21190
rect 5931 21188 5987 21190
rect 6011 21188 6067 21190
rect 6091 21188 6147 21190
rect 5851 20154 5907 20156
rect 5931 20154 5987 20156
rect 6011 20154 6067 20156
rect 6091 20154 6147 20156
rect 5851 20102 5897 20154
rect 5897 20102 5907 20154
rect 5931 20102 5961 20154
rect 5961 20102 5973 20154
rect 5973 20102 5987 20154
rect 6011 20102 6025 20154
rect 6025 20102 6037 20154
rect 6037 20102 6067 20154
rect 6091 20102 6101 20154
rect 6101 20102 6147 20154
rect 5851 20100 5907 20102
rect 5931 20100 5987 20102
rect 6011 20100 6067 20102
rect 6091 20100 6147 20102
rect 5851 19066 5907 19068
rect 5931 19066 5987 19068
rect 6011 19066 6067 19068
rect 6091 19066 6147 19068
rect 5851 19014 5897 19066
rect 5897 19014 5907 19066
rect 5931 19014 5961 19066
rect 5961 19014 5973 19066
rect 5973 19014 5987 19066
rect 6011 19014 6025 19066
rect 6025 19014 6037 19066
rect 6037 19014 6067 19066
rect 6091 19014 6101 19066
rect 6101 19014 6147 19066
rect 5851 19012 5907 19014
rect 5931 19012 5987 19014
rect 6011 19012 6067 19014
rect 6091 19012 6147 19014
rect 5851 17978 5907 17980
rect 5931 17978 5987 17980
rect 6011 17978 6067 17980
rect 6091 17978 6147 17980
rect 5851 17926 5897 17978
rect 5897 17926 5907 17978
rect 5931 17926 5961 17978
rect 5961 17926 5973 17978
rect 5973 17926 5987 17978
rect 6011 17926 6025 17978
rect 6025 17926 6037 17978
rect 6037 17926 6067 17978
rect 6091 17926 6101 17978
rect 6101 17926 6147 17978
rect 5851 17924 5907 17926
rect 5931 17924 5987 17926
rect 6011 17924 6067 17926
rect 6091 17924 6147 17926
rect 7483 72922 7539 72924
rect 7563 72922 7619 72924
rect 7643 72922 7699 72924
rect 7723 72922 7779 72924
rect 7483 72870 7529 72922
rect 7529 72870 7539 72922
rect 7563 72870 7593 72922
rect 7593 72870 7605 72922
rect 7605 72870 7619 72922
rect 7643 72870 7657 72922
rect 7657 72870 7669 72922
rect 7669 72870 7699 72922
rect 7723 72870 7733 72922
rect 7733 72870 7779 72922
rect 7483 72868 7539 72870
rect 7563 72868 7619 72870
rect 7643 72868 7699 72870
rect 7723 72868 7779 72870
rect 9310 77324 9312 77344
rect 9312 77324 9364 77344
rect 9364 77324 9366 77344
rect 9310 77288 9366 77324
rect 9115 76730 9171 76732
rect 9195 76730 9251 76732
rect 9275 76730 9331 76732
rect 9355 76730 9411 76732
rect 9115 76678 9161 76730
rect 9161 76678 9171 76730
rect 9195 76678 9225 76730
rect 9225 76678 9237 76730
rect 9237 76678 9251 76730
rect 9275 76678 9289 76730
rect 9289 76678 9301 76730
rect 9301 76678 9331 76730
rect 9355 76678 9365 76730
rect 9365 76678 9411 76730
rect 9115 76676 9171 76678
rect 9195 76676 9251 76678
rect 9275 76676 9331 76678
rect 9355 76676 9411 76678
rect 9586 77696 9642 77752
rect 10138 76744 10194 76800
rect 10046 76336 10102 76392
rect 9310 75792 9366 75848
rect 9115 75642 9171 75644
rect 9195 75642 9251 75644
rect 9275 75642 9331 75644
rect 9355 75642 9411 75644
rect 9115 75590 9161 75642
rect 9161 75590 9171 75642
rect 9195 75590 9225 75642
rect 9225 75590 9237 75642
rect 9237 75590 9251 75642
rect 9275 75590 9289 75642
rect 9289 75590 9301 75642
rect 9301 75590 9331 75642
rect 9355 75590 9365 75642
rect 9365 75590 9411 75642
rect 9115 75588 9171 75590
rect 9195 75588 9251 75590
rect 9275 75588 9331 75590
rect 9355 75588 9411 75590
rect 9115 74554 9171 74556
rect 9195 74554 9251 74556
rect 9275 74554 9331 74556
rect 9355 74554 9411 74556
rect 9115 74502 9161 74554
rect 9161 74502 9171 74554
rect 9195 74502 9225 74554
rect 9225 74502 9237 74554
rect 9237 74502 9251 74554
rect 9275 74502 9289 74554
rect 9289 74502 9301 74554
rect 9301 74502 9331 74554
rect 9355 74502 9365 74554
rect 9365 74502 9411 74554
rect 9115 74500 9171 74502
rect 9195 74500 9251 74502
rect 9275 74500 9331 74502
rect 9355 74500 9411 74502
rect 8574 71848 8630 71904
rect 7483 71834 7539 71836
rect 7563 71834 7619 71836
rect 7643 71834 7699 71836
rect 7723 71834 7779 71836
rect 7483 71782 7529 71834
rect 7529 71782 7539 71834
rect 7563 71782 7593 71834
rect 7593 71782 7605 71834
rect 7605 71782 7619 71834
rect 7643 71782 7657 71834
rect 7657 71782 7669 71834
rect 7669 71782 7699 71834
rect 7723 71782 7733 71834
rect 7733 71782 7779 71834
rect 7483 71780 7539 71782
rect 7563 71780 7619 71782
rect 7643 71780 7699 71782
rect 7723 71780 7779 71782
rect 7483 70746 7539 70748
rect 7563 70746 7619 70748
rect 7643 70746 7699 70748
rect 7723 70746 7779 70748
rect 7483 70694 7529 70746
rect 7529 70694 7539 70746
rect 7563 70694 7593 70746
rect 7593 70694 7605 70746
rect 7605 70694 7619 70746
rect 7643 70694 7657 70746
rect 7657 70694 7669 70746
rect 7669 70694 7699 70746
rect 7723 70694 7733 70746
rect 7733 70694 7779 70746
rect 7483 70692 7539 70694
rect 7563 70692 7619 70694
rect 7643 70692 7699 70694
rect 7723 70692 7779 70694
rect 7010 51176 7066 51232
rect 7010 51060 7066 51096
rect 7010 51040 7012 51060
rect 7012 51040 7064 51060
rect 7064 51040 7066 51060
rect 7010 50904 7066 50960
rect 7010 49544 7066 49600
rect 7194 51448 7250 51504
rect 7483 69658 7539 69660
rect 7563 69658 7619 69660
rect 7643 69658 7699 69660
rect 7723 69658 7779 69660
rect 7483 69606 7529 69658
rect 7529 69606 7539 69658
rect 7563 69606 7593 69658
rect 7593 69606 7605 69658
rect 7605 69606 7619 69658
rect 7643 69606 7657 69658
rect 7657 69606 7669 69658
rect 7669 69606 7699 69658
rect 7723 69606 7733 69658
rect 7733 69606 7779 69658
rect 7483 69604 7539 69606
rect 7563 69604 7619 69606
rect 7643 69604 7699 69606
rect 7723 69604 7779 69606
rect 7483 68570 7539 68572
rect 7563 68570 7619 68572
rect 7643 68570 7699 68572
rect 7723 68570 7779 68572
rect 7483 68518 7529 68570
rect 7529 68518 7539 68570
rect 7563 68518 7593 68570
rect 7593 68518 7605 68570
rect 7605 68518 7619 68570
rect 7643 68518 7657 68570
rect 7657 68518 7669 68570
rect 7669 68518 7699 68570
rect 7723 68518 7733 68570
rect 7733 68518 7779 68570
rect 7483 68516 7539 68518
rect 7563 68516 7619 68518
rect 7643 68516 7699 68518
rect 7723 68516 7779 68518
rect 7483 67482 7539 67484
rect 7563 67482 7619 67484
rect 7643 67482 7699 67484
rect 7723 67482 7779 67484
rect 7483 67430 7529 67482
rect 7529 67430 7539 67482
rect 7563 67430 7593 67482
rect 7593 67430 7605 67482
rect 7605 67430 7619 67482
rect 7643 67430 7657 67482
rect 7657 67430 7669 67482
rect 7669 67430 7699 67482
rect 7723 67430 7733 67482
rect 7733 67430 7779 67482
rect 7483 67428 7539 67430
rect 7563 67428 7619 67430
rect 7643 67428 7699 67430
rect 7723 67428 7779 67430
rect 7483 66394 7539 66396
rect 7563 66394 7619 66396
rect 7643 66394 7699 66396
rect 7723 66394 7779 66396
rect 7483 66342 7529 66394
rect 7529 66342 7539 66394
rect 7563 66342 7593 66394
rect 7593 66342 7605 66394
rect 7605 66342 7619 66394
rect 7643 66342 7657 66394
rect 7657 66342 7669 66394
rect 7669 66342 7699 66394
rect 7723 66342 7733 66394
rect 7733 66342 7779 66394
rect 7483 66340 7539 66342
rect 7563 66340 7619 66342
rect 7643 66340 7699 66342
rect 7723 66340 7779 66342
rect 7483 65306 7539 65308
rect 7563 65306 7619 65308
rect 7643 65306 7699 65308
rect 7723 65306 7779 65308
rect 7483 65254 7529 65306
rect 7529 65254 7539 65306
rect 7563 65254 7593 65306
rect 7593 65254 7605 65306
rect 7605 65254 7619 65306
rect 7643 65254 7657 65306
rect 7657 65254 7669 65306
rect 7669 65254 7699 65306
rect 7723 65254 7733 65306
rect 7733 65254 7779 65306
rect 7483 65252 7539 65254
rect 7563 65252 7619 65254
rect 7643 65252 7699 65254
rect 7723 65252 7779 65254
rect 7483 64218 7539 64220
rect 7563 64218 7619 64220
rect 7643 64218 7699 64220
rect 7723 64218 7779 64220
rect 7483 64166 7529 64218
rect 7529 64166 7539 64218
rect 7563 64166 7593 64218
rect 7593 64166 7605 64218
rect 7605 64166 7619 64218
rect 7643 64166 7657 64218
rect 7657 64166 7669 64218
rect 7669 64166 7699 64218
rect 7723 64166 7733 64218
rect 7733 64166 7779 64218
rect 7483 64164 7539 64166
rect 7563 64164 7619 64166
rect 7643 64164 7699 64166
rect 7723 64164 7779 64166
rect 7483 63130 7539 63132
rect 7563 63130 7619 63132
rect 7643 63130 7699 63132
rect 7723 63130 7779 63132
rect 7483 63078 7529 63130
rect 7529 63078 7539 63130
rect 7563 63078 7593 63130
rect 7593 63078 7605 63130
rect 7605 63078 7619 63130
rect 7643 63078 7657 63130
rect 7657 63078 7669 63130
rect 7669 63078 7699 63130
rect 7723 63078 7733 63130
rect 7733 63078 7779 63130
rect 7483 63076 7539 63078
rect 7563 63076 7619 63078
rect 7643 63076 7699 63078
rect 7723 63076 7779 63078
rect 7483 62042 7539 62044
rect 7563 62042 7619 62044
rect 7643 62042 7699 62044
rect 7723 62042 7779 62044
rect 7483 61990 7529 62042
rect 7529 61990 7539 62042
rect 7563 61990 7593 62042
rect 7593 61990 7605 62042
rect 7605 61990 7619 62042
rect 7643 61990 7657 62042
rect 7657 61990 7669 62042
rect 7669 61990 7699 62042
rect 7723 61990 7733 62042
rect 7733 61990 7779 62042
rect 7483 61988 7539 61990
rect 7563 61988 7619 61990
rect 7643 61988 7699 61990
rect 7723 61988 7779 61990
rect 7483 60954 7539 60956
rect 7563 60954 7619 60956
rect 7643 60954 7699 60956
rect 7723 60954 7779 60956
rect 7483 60902 7529 60954
rect 7529 60902 7539 60954
rect 7563 60902 7593 60954
rect 7593 60902 7605 60954
rect 7605 60902 7619 60954
rect 7643 60902 7657 60954
rect 7657 60902 7669 60954
rect 7669 60902 7699 60954
rect 7723 60902 7733 60954
rect 7733 60902 7779 60954
rect 7483 60900 7539 60902
rect 7563 60900 7619 60902
rect 7643 60900 7699 60902
rect 7723 60900 7779 60902
rect 7483 59866 7539 59868
rect 7563 59866 7619 59868
rect 7643 59866 7699 59868
rect 7723 59866 7779 59868
rect 7483 59814 7529 59866
rect 7529 59814 7539 59866
rect 7563 59814 7593 59866
rect 7593 59814 7605 59866
rect 7605 59814 7619 59866
rect 7643 59814 7657 59866
rect 7657 59814 7669 59866
rect 7669 59814 7699 59866
rect 7723 59814 7733 59866
rect 7733 59814 7779 59866
rect 7483 59812 7539 59814
rect 7563 59812 7619 59814
rect 7643 59812 7699 59814
rect 7723 59812 7779 59814
rect 7483 58778 7539 58780
rect 7563 58778 7619 58780
rect 7643 58778 7699 58780
rect 7723 58778 7779 58780
rect 7483 58726 7529 58778
rect 7529 58726 7539 58778
rect 7563 58726 7593 58778
rect 7593 58726 7605 58778
rect 7605 58726 7619 58778
rect 7643 58726 7657 58778
rect 7657 58726 7669 58778
rect 7669 58726 7699 58778
rect 7723 58726 7733 58778
rect 7733 58726 7779 58778
rect 7483 58724 7539 58726
rect 7563 58724 7619 58726
rect 7643 58724 7699 58726
rect 7723 58724 7779 58726
rect 7483 57690 7539 57692
rect 7563 57690 7619 57692
rect 7643 57690 7699 57692
rect 7723 57690 7779 57692
rect 7483 57638 7529 57690
rect 7529 57638 7539 57690
rect 7563 57638 7593 57690
rect 7593 57638 7605 57690
rect 7605 57638 7619 57690
rect 7643 57638 7657 57690
rect 7657 57638 7669 57690
rect 7669 57638 7699 57690
rect 7723 57638 7733 57690
rect 7733 57638 7779 57690
rect 7483 57636 7539 57638
rect 7563 57636 7619 57638
rect 7643 57636 7699 57638
rect 7723 57636 7779 57638
rect 7483 56602 7539 56604
rect 7563 56602 7619 56604
rect 7643 56602 7699 56604
rect 7723 56602 7779 56604
rect 7483 56550 7529 56602
rect 7529 56550 7539 56602
rect 7563 56550 7593 56602
rect 7593 56550 7605 56602
rect 7605 56550 7619 56602
rect 7643 56550 7657 56602
rect 7657 56550 7669 56602
rect 7669 56550 7699 56602
rect 7723 56550 7733 56602
rect 7733 56550 7779 56602
rect 7483 56548 7539 56550
rect 7563 56548 7619 56550
rect 7643 56548 7699 56550
rect 7723 56548 7779 56550
rect 8206 68720 8262 68776
rect 8298 67360 8354 67416
rect 8298 66272 8354 66328
rect 8114 60696 8170 60752
rect 7483 55514 7539 55516
rect 7563 55514 7619 55516
rect 7643 55514 7699 55516
rect 7723 55514 7779 55516
rect 7483 55462 7529 55514
rect 7529 55462 7539 55514
rect 7563 55462 7593 55514
rect 7593 55462 7605 55514
rect 7605 55462 7619 55514
rect 7643 55462 7657 55514
rect 7657 55462 7669 55514
rect 7669 55462 7699 55514
rect 7723 55462 7733 55514
rect 7733 55462 7779 55514
rect 7483 55460 7539 55462
rect 7563 55460 7619 55462
rect 7643 55460 7699 55462
rect 7723 55460 7779 55462
rect 7483 54426 7539 54428
rect 7563 54426 7619 54428
rect 7643 54426 7699 54428
rect 7723 54426 7779 54428
rect 7483 54374 7529 54426
rect 7529 54374 7539 54426
rect 7563 54374 7593 54426
rect 7593 54374 7605 54426
rect 7605 54374 7619 54426
rect 7643 54374 7657 54426
rect 7657 54374 7669 54426
rect 7669 54374 7699 54426
rect 7723 54374 7733 54426
rect 7733 54374 7779 54426
rect 7483 54372 7539 54374
rect 7563 54372 7619 54374
rect 7643 54372 7699 54374
rect 7723 54372 7779 54374
rect 7483 53338 7539 53340
rect 7563 53338 7619 53340
rect 7643 53338 7699 53340
rect 7723 53338 7779 53340
rect 7483 53286 7529 53338
rect 7529 53286 7539 53338
rect 7563 53286 7593 53338
rect 7593 53286 7605 53338
rect 7605 53286 7619 53338
rect 7643 53286 7657 53338
rect 7657 53286 7669 53338
rect 7669 53286 7699 53338
rect 7723 53286 7733 53338
rect 7733 53286 7779 53338
rect 7483 53284 7539 53286
rect 7563 53284 7619 53286
rect 7643 53284 7699 53286
rect 7723 53284 7779 53286
rect 7483 52250 7539 52252
rect 7563 52250 7619 52252
rect 7643 52250 7699 52252
rect 7723 52250 7779 52252
rect 7483 52198 7529 52250
rect 7529 52198 7539 52250
rect 7563 52198 7593 52250
rect 7593 52198 7605 52250
rect 7605 52198 7619 52250
rect 7643 52198 7657 52250
rect 7657 52198 7669 52250
rect 7669 52198 7699 52250
rect 7723 52198 7733 52250
rect 7733 52198 7779 52250
rect 7483 52196 7539 52198
rect 7563 52196 7619 52198
rect 7643 52196 7699 52198
rect 7723 52196 7779 52198
rect 7483 51162 7539 51164
rect 7563 51162 7619 51164
rect 7643 51162 7699 51164
rect 7723 51162 7779 51164
rect 7483 51110 7529 51162
rect 7529 51110 7539 51162
rect 7563 51110 7593 51162
rect 7593 51110 7605 51162
rect 7605 51110 7619 51162
rect 7643 51110 7657 51162
rect 7657 51110 7669 51162
rect 7669 51110 7699 51162
rect 7723 51110 7733 51162
rect 7733 51110 7779 51162
rect 7483 51108 7539 51110
rect 7563 51108 7619 51110
rect 7643 51108 7699 51110
rect 7723 51108 7779 51110
rect 7194 46280 7250 46336
rect 6826 42764 6882 42800
rect 6826 42744 6828 42764
rect 6828 42744 6880 42764
rect 6880 42744 6882 42764
rect 6918 42608 6974 42664
rect 7286 43832 7342 43888
rect 7010 38392 7066 38448
rect 7010 38120 7066 38176
rect 7483 50074 7539 50076
rect 7563 50074 7619 50076
rect 7643 50074 7699 50076
rect 7723 50074 7779 50076
rect 7483 50022 7529 50074
rect 7529 50022 7539 50074
rect 7563 50022 7593 50074
rect 7593 50022 7605 50074
rect 7605 50022 7619 50074
rect 7643 50022 7657 50074
rect 7657 50022 7669 50074
rect 7669 50022 7699 50074
rect 7723 50022 7733 50074
rect 7733 50022 7779 50074
rect 7483 50020 7539 50022
rect 7563 50020 7619 50022
rect 7643 50020 7699 50022
rect 7723 50020 7779 50022
rect 7483 48986 7539 48988
rect 7563 48986 7619 48988
rect 7643 48986 7699 48988
rect 7723 48986 7779 48988
rect 7483 48934 7529 48986
rect 7529 48934 7539 48986
rect 7563 48934 7593 48986
rect 7593 48934 7605 48986
rect 7605 48934 7619 48986
rect 7643 48934 7657 48986
rect 7657 48934 7669 48986
rect 7669 48934 7699 48986
rect 7723 48934 7733 48986
rect 7733 48934 7779 48986
rect 7483 48932 7539 48934
rect 7563 48932 7619 48934
rect 7643 48932 7699 48934
rect 7723 48932 7779 48934
rect 7746 48728 7802 48784
rect 7746 48048 7802 48104
rect 7483 47898 7539 47900
rect 7563 47898 7619 47900
rect 7643 47898 7699 47900
rect 7723 47898 7779 47900
rect 7483 47846 7529 47898
rect 7529 47846 7539 47898
rect 7563 47846 7593 47898
rect 7593 47846 7605 47898
rect 7605 47846 7619 47898
rect 7643 47846 7657 47898
rect 7657 47846 7669 47898
rect 7669 47846 7699 47898
rect 7723 47846 7733 47898
rect 7733 47846 7779 47898
rect 7483 47844 7539 47846
rect 7563 47844 7619 47846
rect 7643 47844 7699 47846
rect 7723 47844 7779 47846
rect 7483 46810 7539 46812
rect 7563 46810 7619 46812
rect 7643 46810 7699 46812
rect 7723 46810 7779 46812
rect 7483 46758 7529 46810
rect 7529 46758 7539 46810
rect 7563 46758 7593 46810
rect 7593 46758 7605 46810
rect 7605 46758 7619 46810
rect 7643 46758 7657 46810
rect 7657 46758 7669 46810
rect 7669 46758 7699 46810
rect 7723 46758 7733 46810
rect 7733 46758 7779 46810
rect 7483 46756 7539 46758
rect 7563 46756 7619 46758
rect 7643 46756 7699 46758
rect 7723 46756 7779 46758
rect 7483 45722 7539 45724
rect 7563 45722 7619 45724
rect 7643 45722 7699 45724
rect 7723 45722 7779 45724
rect 7483 45670 7529 45722
rect 7529 45670 7539 45722
rect 7563 45670 7593 45722
rect 7593 45670 7605 45722
rect 7605 45670 7619 45722
rect 7643 45670 7657 45722
rect 7657 45670 7669 45722
rect 7669 45670 7699 45722
rect 7723 45670 7733 45722
rect 7733 45670 7779 45722
rect 7483 45668 7539 45670
rect 7563 45668 7619 45670
rect 7643 45668 7699 45670
rect 7723 45668 7779 45670
rect 7483 44634 7539 44636
rect 7563 44634 7619 44636
rect 7643 44634 7699 44636
rect 7723 44634 7779 44636
rect 7483 44582 7529 44634
rect 7529 44582 7539 44634
rect 7563 44582 7593 44634
rect 7593 44582 7605 44634
rect 7605 44582 7619 44634
rect 7643 44582 7657 44634
rect 7657 44582 7669 44634
rect 7669 44582 7699 44634
rect 7723 44582 7733 44634
rect 7733 44582 7779 44634
rect 7483 44580 7539 44582
rect 7563 44580 7619 44582
rect 7643 44580 7699 44582
rect 7723 44580 7779 44582
rect 7562 44240 7618 44296
rect 7483 43546 7539 43548
rect 7563 43546 7619 43548
rect 7643 43546 7699 43548
rect 7723 43546 7779 43548
rect 7483 43494 7529 43546
rect 7529 43494 7539 43546
rect 7563 43494 7593 43546
rect 7593 43494 7605 43546
rect 7605 43494 7619 43546
rect 7643 43494 7657 43546
rect 7657 43494 7669 43546
rect 7669 43494 7699 43546
rect 7723 43494 7733 43546
rect 7733 43494 7779 43546
rect 7483 43492 7539 43494
rect 7563 43492 7619 43494
rect 7643 43492 7699 43494
rect 7723 43492 7779 43494
rect 7483 42458 7539 42460
rect 7563 42458 7619 42460
rect 7643 42458 7699 42460
rect 7723 42458 7779 42460
rect 7483 42406 7529 42458
rect 7529 42406 7539 42458
rect 7563 42406 7593 42458
rect 7593 42406 7605 42458
rect 7605 42406 7619 42458
rect 7643 42406 7657 42458
rect 7657 42406 7669 42458
rect 7669 42406 7699 42458
rect 7723 42406 7733 42458
rect 7733 42406 7779 42458
rect 7483 42404 7539 42406
rect 7563 42404 7619 42406
rect 7643 42404 7699 42406
rect 7723 42404 7779 42406
rect 7483 41370 7539 41372
rect 7563 41370 7619 41372
rect 7643 41370 7699 41372
rect 7723 41370 7779 41372
rect 7483 41318 7529 41370
rect 7529 41318 7539 41370
rect 7563 41318 7593 41370
rect 7593 41318 7605 41370
rect 7605 41318 7619 41370
rect 7643 41318 7657 41370
rect 7657 41318 7669 41370
rect 7669 41318 7699 41370
rect 7723 41318 7733 41370
rect 7733 41318 7779 41370
rect 7483 41316 7539 41318
rect 7563 41316 7619 41318
rect 7643 41316 7699 41318
rect 7723 41316 7779 41318
rect 8298 60968 8354 61024
rect 8298 51312 8354 51368
rect 8298 51176 8354 51232
rect 8114 50260 8116 50280
rect 8116 50260 8168 50280
rect 8168 50260 8170 50280
rect 8114 50224 8170 50260
rect 8206 48864 8262 48920
rect 8206 48592 8262 48648
rect 8206 47912 8262 47968
rect 8206 46996 8208 47016
rect 8208 46996 8260 47016
rect 8260 46996 8262 47016
rect 8206 46960 8262 46996
rect 8022 46280 8078 46336
rect 8206 44648 8262 44704
rect 7483 40282 7539 40284
rect 7563 40282 7619 40284
rect 7643 40282 7699 40284
rect 7723 40282 7779 40284
rect 7483 40230 7529 40282
rect 7529 40230 7539 40282
rect 7563 40230 7593 40282
rect 7593 40230 7605 40282
rect 7605 40230 7619 40282
rect 7643 40230 7657 40282
rect 7657 40230 7669 40282
rect 7669 40230 7699 40282
rect 7723 40230 7733 40282
rect 7733 40230 7779 40282
rect 7483 40228 7539 40230
rect 7563 40228 7619 40230
rect 7643 40228 7699 40230
rect 7723 40228 7779 40230
rect 7470 39344 7526 39400
rect 7483 39194 7539 39196
rect 7563 39194 7619 39196
rect 7643 39194 7699 39196
rect 7723 39194 7779 39196
rect 7483 39142 7529 39194
rect 7529 39142 7539 39194
rect 7563 39142 7593 39194
rect 7593 39142 7605 39194
rect 7605 39142 7619 39194
rect 7643 39142 7657 39194
rect 7657 39142 7669 39194
rect 7669 39142 7699 39194
rect 7723 39142 7733 39194
rect 7733 39142 7779 39194
rect 7483 39140 7539 39142
rect 7563 39140 7619 39142
rect 7643 39140 7699 39142
rect 7723 39140 7779 39142
rect 7746 38256 7802 38312
rect 7483 38106 7539 38108
rect 7563 38106 7619 38108
rect 7643 38106 7699 38108
rect 7723 38106 7779 38108
rect 7483 38054 7529 38106
rect 7529 38054 7539 38106
rect 7563 38054 7593 38106
rect 7593 38054 7605 38106
rect 7605 38054 7619 38106
rect 7643 38054 7657 38106
rect 7657 38054 7669 38106
rect 7669 38054 7699 38106
rect 7723 38054 7733 38106
rect 7733 38054 7779 38106
rect 7483 38052 7539 38054
rect 7563 38052 7619 38054
rect 7643 38052 7699 38054
rect 7723 38052 7779 38054
rect 7483 37018 7539 37020
rect 7563 37018 7619 37020
rect 7643 37018 7699 37020
rect 7723 37018 7779 37020
rect 7483 36966 7529 37018
rect 7529 36966 7539 37018
rect 7563 36966 7593 37018
rect 7593 36966 7605 37018
rect 7605 36966 7619 37018
rect 7643 36966 7657 37018
rect 7657 36966 7669 37018
rect 7669 36966 7699 37018
rect 7723 36966 7733 37018
rect 7733 36966 7779 37018
rect 7483 36964 7539 36966
rect 7563 36964 7619 36966
rect 7643 36964 7699 36966
rect 7723 36964 7779 36966
rect 7483 35930 7539 35932
rect 7563 35930 7619 35932
rect 7643 35930 7699 35932
rect 7723 35930 7779 35932
rect 7483 35878 7529 35930
rect 7529 35878 7539 35930
rect 7563 35878 7593 35930
rect 7593 35878 7605 35930
rect 7605 35878 7619 35930
rect 7643 35878 7657 35930
rect 7657 35878 7669 35930
rect 7669 35878 7699 35930
rect 7723 35878 7733 35930
rect 7733 35878 7779 35930
rect 7483 35876 7539 35878
rect 7563 35876 7619 35878
rect 7643 35876 7699 35878
rect 7723 35876 7779 35878
rect 7483 34842 7539 34844
rect 7563 34842 7619 34844
rect 7643 34842 7699 34844
rect 7723 34842 7779 34844
rect 7483 34790 7529 34842
rect 7529 34790 7539 34842
rect 7563 34790 7593 34842
rect 7593 34790 7605 34842
rect 7605 34790 7619 34842
rect 7643 34790 7657 34842
rect 7657 34790 7669 34842
rect 7669 34790 7699 34842
rect 7723 34790 7733 34842
rect 7733 34790 7779 34842
rect 7483 34788 7539 34790
rect 7563 34788 7619 34790
rect 7643 34788 7699 34790
rect 7723 34788 7779 34790
rect 7483 33754 7539 33756
rect 7563 33754 7619 33756
rect 7643 33754 7699 33756
rect 7723 33754 7779 33756
rect 7483 33702 7529 33754
rect 7529 33702 7539 33754
rect 7563 33702 7593 33754
rect 7593 33702 7605 33754
rect 7605 33702 7619 33754
rect 7643 33702 7657 33754
rect 7657 33702 7669 33754
rect 7669 33702 7699 33754
rect 7723 33702 7733 33754
rect 7733 33702 7779 33754
rect 7483 33700 7539 33702
rect 7563 33700 7619 33702
rect 7643 33700 7699 33702
rect 7723 33700 7779 33702
rect 7483 32666 7539 32668
rect 7563 32666 7619 32668
rect 7643 32666 7699 32668
rect 7723 32666 7779 32668
rect 7483 32614 7529 32666
rect 7529 32614 7539 32666
rect 7563 32614 7593 32666
rect 7593 32614 7605 32666
rect 7605 32614 7619 32666
rect 7643 32614 7657 32666
rect 7657 32614 7669 32666
rect 7669 32614 7699 32666
rect 7723 32614 7733 32666
rect 7733 32614 7779 32666
rect 7483 32612 7539 32614
rect 7563 32612 7619 32614
rect 7643 32612 7699 32614
rect 7723 32612 7779 32614
rect 7483 31578 7539 31580
rect 7563 31578 7619 31580
rect 7643 31578 7699 31580
rect 7723 31578 7779 31580
rect 7483 31526 7529 31578
rect 7529 31526 7539 31578
rect 7563 31526 7593 31578
rect 7593 31526 7605 31578
rect 7605 31526 7619 31578
rect 7643 31526 7657 31578
rect 7657 31526 7669 31578
rect 7669 31526 7699 31578
rect 7723 31526 7733 31578
rect 7733 31526 7779 31578
rect 7483 31524 7539 31526
rect 7563 31524 7619 31526
rect 7643 31524 7699 31526
rect 7723 31524 7779 31526
rect 7483 30490 7539 30492
rect 7563 30490 7619 30492
rect 7643 30490 7699 30492
rect 7723 30490 7779 30492
rect 7483 30438 7529 30490
rect 7529 30438 7539 30490
rect 7563 30438 7593 30490
rect 7593 30438 7605 30490
rect 7605 30438 7619 30490
rect 7643 30438 7657 30490
rect 7657 30438 7669 30490
rect 7669 30438 7699 30490
rect 7723 30438 7733 30490
rect 7733 30438 7779 30490
rect 7483 30436 7539 30438
rect 7563 30436 7619 30438
rect 7643 30436 7699 30438
rect 7723 30436 7779 30438
rect 7483 29402 7539 29404
rect 7563 29402 7619 29404
rect 7643 29402 7699 29404
rect 7723 29402 7779 29404
rect 7483 29350 7529 29402
rect 7529 29350 7539 29402
rect 7563 29350 7593 29402
rect 7593 29350 7605 29402
rect 7605 29350 7619 29402
rect 7643 29350 7657 29402
rect 7657 29350 7669 29402
rect 7669 29350 7699 29402
rect 7723 29350 7733 29402
rect 7733 29350 7779 29402
rect 7483 29348 7539 29350
rect 7563 29348 7619 29350
rect 7643 29348 7699 29350
rect 7723 29348 7779 29350
rect 5851 16890 5907 16892
rect 5931 16890 5987 16892
rect 6011 16890 6067 16892
rect 6091 16890 6147 16892
rect 5851 16838 5897 16890
rect 5897 16838 5907 16890
rect 5931 16838 5961 16890
rect 5961 16838 5973 16890
rect 5973 16838 5987 16890
rect 6011 16838 6025 16890
rect 6025 16838 6037 16890
rect 6037 16838 6067 16890
rect 6091 16838 6101 16890
rect 6101 16838 6147 16890
rect 5851 16836 5907 16838
rect 5931 16836 5987 16838
rect 6011 16836 6067 16838
rect 6091 16836 6147 16838
rect 5851 15802 5907 15804
rect 5931 15802 5987 15804
rect 6011 15802 6067 15804
rect 6091 15802 6147 15804
rect 5851 15750 5897 15802
rect 5897 15750 5907 15802
rect 5931 15750 5961 15802
rect 5961 15750 5973 15802
rect 5973 15750 5987 15802
rect 6011 15750 6025 15802
rect 6025 15750 6037 15802
rect 6037 15750 6067 15802
rect 6091 15750 6101 15802
rect 6101 15750 6147 15802
rect 5851 15748 5907 15750
rect 5931 15748 5987 15750
rect 6011 15748 6067 15750
rect 6091 15748 6147 15750
rect 5851 14714 5907 14716
rect 5931 14714 5987 14716
rect 6011 14714 6067 14716
rect 6091 14714 6147 14716
rect 5851 14662 5897 14714
rect 5897 14662 5907 14714
rect 5931 14662 5961 14714
rect 5961 14662 5973 14714
rect 5973 14662 5987 14714
rect 6011 14662 6025 14714
rect 6025 14662 6037 14714
rect 6037 14662 6067 14714
rect 6091 14662 6101 14714
rect 6101 14662 6147 14714
rect 5851 14660 5907 14662
rect 5931 14660 5987 14662
rect 6011 14660 6067 14662
rect 6091 14660 6147 14662
rect 6182 14456 6238 14512
rect 5851 13626 5907 13628
rect 5931 13626 5987 13628
rect 6011 13626 6067 13628
rect 6091 13626 6147 13628
rect 5851 13574 5897 13626
rect 5897 13574 5907 13626
rect 5931 13574 5961 13626
rect 5961 13574 5973 13626
rect 5973 13574 5987 13626
rect 6011 13574 6025 13626
rect 6025 13574 6037 13626
rect 6037 13574 6067 13626
rect 6091 13574 6101 13626
rect 6101 13574 6147 13626
rect 5851 13572 5907 13574
rect 5931 13572 5987 13574
rect 6011 13572 6067 13574
rect 6091 13572 6147 13574
rect 6366 14728 6422 14784
rect 7483 28314 7539 28316
rect 7563 28314 7619 28316
rect 7643 28314 7699 28316
rect 7723 28314 7779 28316
rect 7483 28262 7529 28314
rect 7529 28262 7539 28314
rect 7563 28262 7593 28314
rect 7593 28262 7605 28314
rect 7605 28262 7619 28314
rect 7643 28262 7657 28314
rect 7657 28262 7669 28314
rect 7669 28262 7699 28314
rect 7723 28262 7733 28314
rect 7733 28262 7779 28314
rect 7483 28260 7539 28262
rect 7563 28260 7619 28262
rect 7643 28260 7699 28262
rect 7723 28260 7779 28262
rect 7483 27226 7539 27228
rect 7563 27226 7619 27228
rect 7643 27226 7699 27228
rect 7723 27226 7779 27228
rect 7483 27174 7529 27226
rect 7529 27174 7539 27226
rect 7563 27174 7593 27226
rect 7593 27174 7605 27226
rect 7605 27174 7619 27226
rect 7643 27174 7657 27226
rect 7657 27174 7669 27226
rect 7669 27174 7699 27226
rect 7723 27174 7733 27226
rect 7733 27174 7779 27226
rect 7483 27172 7539 27174
rect 7563 27172 7619 27174
rect 7643 27172 7699 27174
rect 7723 27172 7779 27174
rect 8390 50360 8446 50416
rect 8206 40296 8262 40352
rect 8114 38392 8170 38448
rect 8114 37984 8170 38040
rect 8114 37204 8116 37224
rect 8116 37204 8168 37224
rect 8168 37204 8170 37224
rect 8114 37168 8170 37204
rect 8114 37068 8116 37088
rect 8116 37068 8168 37088
rect 8168 37068 8170 37088
rect 8114 37032 8170 37068
rect 8114 36644 8170 36680
rect 8114 36624 8116 36644
rect 8116 36624 8168 36644
rect 8168 36624 8170 36644
rect 8114 35128 8170 35184
rect 7483 26138 7539 26140
rect 7563 26138 7619 26140
rect 7643 26138 7699 26140
rect 7723 26138 7779 26140
rect 7483 26086 7529 26138
rect 7529 26086 7539 26138
rect 7563 26086 7593 26138
rect 7593 26086 7605 26138
rect 7605 26086 7619 26138
rect 7643 26086 7657 26138
rect 7657 26086 7669 26138
rect 7669 26086 7699 26138
rect 7723 26086 7733 26138
rect 7733 26086 7779 26138
rect 7483 26084 7539 26086
rect 7563 26084 7619 26086
rect 7643 26084 7699 26086
rect 7723 26084 7779 26086
rect 7483 25050 7539 25052
rect 7563 25050 7619 25052
rect 7643 25050 7699 25052
rect 7723 25050 7779 25052
rect 7483 24998 7529 25050
rect 7529 24998 7539 25050
rect 7563 24998 7593 25050
rect 7593 24998 7605 25050
rect 7605 24998 7619 25050
rect 7643 24998 7657 25050
rect 7657 24998 7669 25050
rect 7669 24998 7699 25050
rect 7723 24998 7733 25050
rect 7733 24998 7779 25050
rect 7483 24996 7539 24998
rect 7563 24996 7619 24998
rect 7643 24996 7699 24998
rect 7723 24996 7779 24998
rect 7483 23962 7539 23964
rect 7563 23962 7619 23964
rect 7643 23962 7699 23964
rect 7723 23962 7779 23964
rect 7483 23910 7529 23962
rect 7529 23910 7539 23962
rect 7563 23910 7593 23962
rect 7593 23910 7605 23962
rect 7605 23910 7619 23962
rect 7643 23910 7657 23962
rect 7657 23910 7669 23962
rect 7669 23910 7699 23962
rect 7723 23910 7733 23962
rect 7733 23910 7779 23962
rect 7483 23908 7539 23910
rect 7563 23908 7619 23910
rect 7643 23908 7699 23910
rect 7723 23908 7779 23910
rect 7483 22874 7539 22876
rect 7563 22874 7619 22876
rect 7643 22874 7699 22876
rect 7723 22874 7779 22876
rect 7483 22822 7529 22874
rect 7529 22822 7539 22874
rect 7563 22822 7593 22874
rect 7593 22822 7605 22874
rect 7605 22822 7619 22874
rect 7643 22822 7657 22874
rect 7657 22822 7669 22874
rect 7669 22822 7699 22874
rect 7723 22822 7733 22874
rect 7733 22822 7779 22874
rect 7483 22820 7539 22822
rect 7563 22820 7619 22822
rect 7643 22820 7699 22822
rect 7723 22820 7779 22822
rect 7483 21786 7539 21788
rect 7563 21786 7619 21788
rect 7643 21786 7699 21788
rect 7723 21786 7779 21788
rect 7483 21734 7529 21786
rect 7529 21734 7539 21786
rect 7563 21734 7593 21786
rect 7593 21734 7605 21786
rect 7605 21734 7619 21786
rect 7643 21734 7657 21786
rect 7657 21734 7669 21786
rect 7669 21734 7699 21786
rect 7723 21734 7733 21786
rect 7733 21734 7779 21786
rect 7483 21732 7539 21734
rect 7563 21732 7619 21734
rect 7643 21732 7699 21734
rect 7723 21732 7779 21734
rect 7483 20698 7539 20700
rect 7563 20698 7619 20700
rect 7643 20698 7699 20700
rect 7723 20698 7779 20700
rect 7483 20646 7529 20698
rect 7529 20646 7539 20698
rect 7563 20646 7593 20698
rect 7593 20646 7605 20698
rect 7605 20646 7619 20698
rect 7643 20646 7657 20698
rect 7657 20646 7669 20698
rect 7669 20646 7699 20698
rect 7723 20646 7733 20698
rect 7733 20646 7779 20698
rect 7483 20644 7539 20646
rect 7563 20644 7619 20646
rect 7643 20644 7699 20646
rect 7723 20644 7779 20646
rect 8114 21956 8170 21992
rect 8114 21936 8116 21956
rect 8116 21936 8168 21956
rect 8168 21936 8170 21956
rect 8114 20304 8170 20360
rect 7483 19610 7539 19612
rect 7563 19610 7619 19612
rect 7643 19610 7699 19612
rect 7723 19610 7779 19612
rect 7483 19558 7529 19610
rect 7529 19558 7539 19610
rect 7563 19558 7593 19610
rect 7593 19558 7605 19610
rect 7605 19558 7619 19610
rect 7643 19558 7657 19610
rect 7657 19558 7669 19610
rect 7669 19558 7699 19610
rect 7723 19558 7733 19610
rect 7733 19558 7779 19610
rect 7483 19556 7539 19558
rect 7563 19556 7619 19558
rect 7643 19556 7699 19558
rect 7723 19556 7779 19558
rect 8114 19488 8170 19544
rect 7483 18522 7539 18524
rect 7563 18522 7619 18524
rect 7643 18522 7699 18524
rect 7723 18522 7779 18524
rect 7483 18470 7529 18522
rect 7529 18470 7539 18522
rect 7563 18470 7593 18522
rect 7593 18470 7605 18522
rect 7605 18470 7619 18522
rect 7643 18470 7657 18522
rect 7657 18470 7669 18522
rect 7669 18470 7699 18522
rect 7723 18470 7733 18522
rect 7733 18470 7779 18522
rect 7483 18468 7539 18470
rect 7563 18468 7619 18470
rect 7643 18468 7699 18470
rect 7723 18468 7779 18470
rect 5851 12538 5907 12540
rect 5931 12538 5987 12540
rect 6011 12538 6067 12540
rect 6091 12538 6147 12540
rect 5851 12486 5897 12538
rect 5897 12486 5907 12538
rect 5931 12486 5961 12538
rect 5961 12486 5973 12538
rect 5973 12486 5987 12538
rect 6011 12486 6025 12538
rect 6025 12486 6037 12538
rect 6037 12486 6067 12538
rect 6091 12486 6101 12538
rect 6101 12486 6147 12538
rect 5851 12484 5907 12486
rect 5931 12484 5987 12486
rect 6011 12484 6067 12486
rect 6091 12484 6147 12486
rect 6274 12960 6330 13016
rect 5906 12180 5908 12200
rect 5908 12180 5960 12200
rect 5960 12180 5962 12200
rect 5906 12144 5962 12180
rect 5851 11450 5907 11452
rect 5931 11450 5987 11452
rect 6011 11450 6067 11452
rect 6091 11450 6147 11452
rect 5851 11398 5897 11450
rect 5897 11398 5907 11450
rect 5931 11398 5961 11450
rect 5961 11398 5973 11450
rect 5973 11398 5987 11450
rect 6011 11398 6025 11450
rect 6025 11398 6037 11450
rect 6037 11398 6067 11450
rect 6091 11398 6101 11450
rect 6101 11398 6147 11450
rect 5851 11396 5907 11398
rect 5931 11396 5987 11398
rect 6011 11396 6067 11398
rect 6091 11396 6147 11398
rect 5851 10362 5907 10364
rect 5931 10362 5987 10364
rect 6011 10362 6067 10364
rect 6091 10362 6147 10364
rect 5851 10310 5897 10362
rect 5897 10310 5907 10362
rect 5931 10310 5961 10362
rect 5961 10310 5973 10362
rect 5973 10310 5987 10362
rect 6011 10310 6025 10362
rect 6025 10310 6037 10362
rect 6037 10310 6067 10362
rect 6091 10310 6101 10362
rect 6101 10310 6147 10362
rect 5851 10308 5907 10310
rect 5931 10308 5987 10310
rect 6011 10308 6067 10310
rect 6091 10308 6147 10310
rect 5851 9274 5907 9276
rect 5931 9274 5987 9276
rect 6011 9274 6067 9276
rect 6091 9274 6147 9276
rect 5851 9222 5897 9274
rect 5897 9222 5907 9274
rect 5931 9222 5961 9274
rect 5961 9222 5973 9274
rect 5973 9222 5987 9274
rect 6011 9222 6025 9274
rect 6025 9222 6037 9274
rect 6037 9222 6067 9274
rect 6091 9222 6101 9274
rect 6101 9222 6147 9274
rect 5851 9220 5907 9222
rect 5931 9220 5987 9222
rect 6011 9220 6067 9222
rect 6091 9220 6147 9222
rect 5851 8186 5907 8188
rect 5931 8186 5987 8188
rect 6011 8186 6067 8188
rect 6091 8186 6147 8188
rect 5851 8134 5897 8186
rect 5897 8134 5907 8186
rect 5931 8134 5961 8186
rect 5961 8134 5973 8186
rect 5973 8134 5987 8186
rect 6011 8134 6025 8186
rect 6025 8134 6037 8186
rect 6037 8134 6067 8186
rect 6091 8134 6101 8186
rect 6101 8134 6147 8186
rect 5851 8132 5907 8134
rect 5931 8132 5987 8134
rect 6011 8132 6067 8134
rect 6091 8132 6147 8134
rect 5851 7098 5907 7100
rect 5931 7098 5987 7100
rect 6011 7098 6067 7100
rect 6091 7098 6147 7100
rect 5851 7046 5897 7098
rect 5897 7046 5907 7098
rect 5931 7046 5961 7098
rect 5961 7046 5973 7098
rect 5973 7046 5987 7098
rect 6011 7046 6025 7098
rect 6025 7046 6037 7098
rect 6037 7046 6067 7098
rect 6091 7046 6101 7098
rect 6101 7046 6147 7098
rect 5851 7044 5907 7046
rect 5931 7044 5987 7046
rect 6011 7044 6067 7046
rect 6091 7044 6147 7046
rect 6918 15952 6974 16008
rect 6918 14864 6974 14920
rect 6918 13776 6974 13832
rect 7838 18128 7894 18184
rect 7286 16632 7342 16688
rect 7483 17434 7539 17436
rect 7563 17434 7619 17436
rect 7643 17434 7699 17436
rect 7723 17434 7779 17436
rect 7483 17382 7529 17434
rect 7529 17382 7539 17434
rect 7563 17382 7593 17434
rect 7593 17382 7605 17434
rect 7605 17382 7619 17434
rect 7643 17382 7657 17434
rect 7657 17382 7669 17434
rect 7669 17382 7699 17434
rect 7723 17382 7733 17434
rect 7733 17382 7779 17434
rect 7483 17380 7539 17382
rect 7563 17380 7619 17382
rect 7643 17380 7699 17382
rect 7723 17380 7779 17382
rect 7102 15408 7158 15464
rect 7483 16346 7539 16348
rect 7563 16346 7619 16348
rect 7643 16346 7699 16348
rect 7723 16346 7779 16348
rect 7483 16294 7529 16346
rect 7529 16294 7539 16346
rect 7563 16294 7593 16346
rect 7593 16294 7605 16346
rect 7605 16294 7619 16346
rect 7643 16294 7657 16346
rect 7657 16294 7669 16346
rect 7669 16294 7699 16346
rect 7723 16294 7733 16346
rect 7733 16294 7779 16346
rect 7483 16292 7539 16294
rect 7563 16292 7619 16294
rect 7643 16292 7699 16294
rect 7723 16292 7779 16294
rect 7930 17176 7986 17232
rect 7483 15258 7539 15260
rect 7563 15258 7619 15260
rect 7643 15258 7699 15260
rect 7723 15258 7779 15260
rect 7483 15206 7529 15258
rect 7529 15206 7539 15258
rect 7563 15206 7593 15258
rect 7593 15206 7605 15258
rect 7605 15206 7619 15258
rect 7643 15206 7657 15258
rect 7657 15206 7669 15258
rect 7669 15206 7699 15258
rect 7723 15206 7733 15258
rect 7733 15206 7779 15258
rect 7483 15204 7539 15206
rect 7563 15204 7619 15206
rect 7643 15204 7699 15206
rect 7723 15204 7779 15206
rect 7930 15156 7986 15192
rect 7930 15136 7932 15156
rect 7932 15136 7984 15156
rect 7984 15136 7986 15156
rect 7286 14592 7342 14648
rect 7654 14456 7710 14512
rect 7194 14320 7250 14376
rect 7102 13912 7158 13968
rect 7483 14170 7539 14172
rect 7563 14170 7619 14172
rect 7643 14170 7699 14172
rect 7723 14170 7779 14172
rect 7483 14118 7529 14170
rect 7529 14118 7539 14170
rect 7563 14118 7593 14170
rect 7593 14118 7605 14170
rect 7605 14118 7619 14170
rect 7643 14118 7657 14170
rect 7657 14118 7669 14170
rect 7669 14118 7699 14170
rect 7723 14118 7733 14170
rect 7733 14118 7779 14170
rect 7483 14116 7539 14118
rect 7563 14116 7619 14118
rect 7643 14116 7699 14118
rect 7723 14116 7779 14118
rect 7654 13524 7710 13560
rect 7654 13504 7656 13524
rect 7656 13504 7708 13524
rect 7708 13504 7710 13524
rect 7483 13082 7539 13084
rect 7563 13082 7619 13084
rect 7643 13082 7699 13084
rect 7723 13082 7779 13084
rect 7483 13030 7529 13082
rect 7529 13030 7539 13082
rect 7563 13030 7593 13082
rect 7593 13030 7605 13082
rect 7605 13030 7619 13082
rect 7643 13030 7657 13082
rect 7657 13030 7669 13082
rect 7669 13030 7699 13082
rect 7723 13030 7733 13082
rect 7733 13030 7779 13082
rect 7483 13028 7539 13030
rect 7563 13028 7619 13030
rect 7643 13028 7699 13030
rect 7723 13028 7779 13030
rect 7194 12824 7250 12880
rect 6918 12688 6974 12744
rect 5851 6010 5907 6012
rect 5931 6010 5987 6012
rect 6011 6010 6067 6012
rect 6091 6010 6147 6012
rect 5851 5958 5897 6010
rect 5897 5958 5907 6010
rect 5931 5958 5961 6010
rect 5961 5958 5973 6010
rect 5973 5958 5987 6010
rect 6011 5958 6025 6010
rect 6025 5958 6037 6010
rect 6037 5958 6067 6010
rect 6091 5958 6101 6010
rect 6101 5958 6147 6010
rect 5851 5956 5907 5958
rect 5931 5956 5987 5958
rect 6011 5956 6067 5958
rect 6091 5956 6147 5958
rect 7286 11192 7342 11248
rect 7483 11994 7539 11996
rect 7563 11994 7619 11996
rect 7643 11994 7699 11996
rect 7723 11994 7779 11996
rect 7483 11942 7529 11994
rect 7529 11942 7539 11994
rect 7563 11942 7593 11994
rect 7593 11942 7605 11994
rect 7605 11942 7619 11994
rect 7643 11942 7657 11994
rect 7657 11942 7669 11994
rect 7669 11942 7699 11994
rect 7723 11942 7733 11994
rect 7733 11942 7779 11994
rect 7483 11940 7539 11942
rect 7563 11940 7619 11942
rect 7643 11940 7699 11942
rect 7723 11940 7779 11942
rect 8114 13368 8170 13424
rect 9494 73516 9496 73536
rect 9496 73516 9548 73536
rect 9548 73516 9550 73536
rect 9494 73480 9550 73516
rect 9115 73466 9171 73468
rect 9195 73466 9251 73468
rect 9275 73466 9331 73468
rect 9355 73466 9411 73468
rect 9115 73414 9161 73466
rect 9161 73414 9171 73466
rect 9195 73414 9225 73466
rect 9225 73414 9237 73466
rect 9237 73414 9251 73466
rect 9275 73414 9289 73466
rect 9289 73414 9301 73466
rect 9301 73414 9331 73466
rect 9355 73414 9365 73466
rect 9365 73414 9411 73466
rect 9115 73412 9171 73414
rect 9195 73412 9251 73414
rect 9275 73412 9331 73414
rect 9355 73412 9411 73414
rect 10046 75384 10102 75440
rect 10966 74876 10968 74896
rect 10968 74876 11020 74896
rect 11020 74876 11022 74896
rect 10966 74840 11022 74876
rect 10138 74432 10194 74488
rect 10046 73888 10102 73944
rect 10046 72936 10102 72992
rect 9310 72548 9366 72584
rect 9310 72528 9312 72548
rect 9312 72528 9364 72548
rect 9364 72528 9366 72548
rect 9115 72378 9171 72380
rect 9195 72378 9251 72380
rect 9275 72378 9331 72380
rect 9355 72378 9411 72380
rect 9115 72326 9161 72378
rect 9161 72326 9171 72378
rect 9195 72326 9225 72378
rect 9225 72326 9237 72378
rect 9237 72326 9251 72378
rect 9275 72326 9289 72378
rect 9289 72326 9301 72378
rect 9301 72326 9331 72378
rect 9355 72326 9365 72378
rect 9365 72326 9411 72378
rect 9115 72324 9171 72326
rect 9195 72324 9251 72326
rect 9275 72324 9331 72326
rect 9355 72324 9411 72326
rect 9310 71984 9366 72040
rect 9115 71290 9171 71292
rect 9195 71290 9251 71292
rect 9275 71290 9331 71292
rect 9355 71290 9411 71292
rect 9115 71238 9161 71290
rect 9161 71238 9171 71290
rect 9195 71238 9225 71290
rect 9225 71238 9237 71290
rect 9237 71238 9251 71290
rect 9275 71238 9289 71290
rect 9289 71238 9301 71290
rect 9301 71238 9331 71290
rect 9355 71238 9365 71290
rect 9365 71238 9411 71290
rect 9115 71236 9171 71238
rect 9195 71236 9251 71238
rect 9275 71236 9331 71238
rect 9355 71236 9411 71238
rect 9115 70202 9171 70204
rect 9195 70202 9251 70204
rect 9275 70202 9331 70204
rect 9355 70202 9411 70204
rect 9115 70150 9161 70202
rect 9161 70150 9171 70202
rect 9195 70150 9225 70202
rect 9225 70150 9237 70202
rect 9237 70150 9251 70202
rect 9275 70150 9289 70202
rect 9289 70150 9301 70202
rect 9301 70150 9331 70202
rect 9355 70150 9365 70202
rect 9365 70150 9411 70202
rect 9115 70148 9171 70150
rect 9195 70148 9251 70150
rect 9275 70148 9331 70150
rect 9355 70148 9411 70150
rect 9034 69264 9090 69320
rect 9494 69128 9550 69184
rect 9115 69114 9171 69116
rect 9195 69114 9251 69116
rect 9275 69114 9331 69116
rect 9355 69114 9411 69116
rect 9115 69062 9161 69114
rect 9161 69062 9171 69114
rect 9195 69062 9225 69114
rect 9225 69062 9237 69114
rect 9237 69062 9251 69114
rect 9275 69062 9289 69114
rect 9289 69062 9301 69114
rect 9301 69062 9331 69114
rect 9355 69062 9365 69114
rect 9365 69062 9411 69114
rect 9115 69060 9171 69062
rect 9195 69060 9251 69062
rect 9275 69060 9331 69062
rect 9355 69060 9411 69062
rect 10138 71576 10194 71632
rect 10046 71032 10102 71088
rect 10138 70624 10194 70680
rect 10046 70080 10102 70136
rect 9586 68312 9642 68368
rect 8758 67768 8814 67824
rect 9115 68026 9171 68028
rect 9195 68026 9251 68028
rect 9275 68026 9331 68028
rect 9355 68026 9411 68028
rect 9115 67974 9161 68026
rect 9161 67974 9171 68026
rect 9195 67974 9225 68026
rect 9225 67974 9237 68026
rect 9237 67974 9251 68026
rect 9275 67974 9289 68026
rect 9289 67974 9301 68026
rect 9301 67974 9331 68026
rect 9355 67974 9365 68026
rect 9365 67974 9411 68026
rect 9115 67972 9171 67974
rect 9195 67972 9251 67974
rect 9275 67972 9331 67974
rect 9355 67972 9411 67974
rect 9402 67632 9458 67688
rect 10414 69672 10470 69728
rect 9115 66938 9171 66940
rect 9195 66938 9251 66940
rect 9275 66938 9331 66940
rect 9355 66938 9411 66940
rect 9115 66886 9161 66938
rect 9161 66886 9171 66938
rect 9195 66886 9225 66938
rect 9225 66886 9237 66938
rect 9237 66886 9251 66938
rect 9275 66886 9289 66938
rect 9289 66886 9301 66938
rect 9301 66886 9331 66938
rect 9355 66886 9365 66938
rect 9365 66886 9411 66938
rect 9115 66884 9171 66886
rect 9195 66884 9251 66886
rect 9275 66884 9331 66886
rect 9355 66884 9411 66886
rect 9494 66816 9550 66872
rect 9402 66580 9404 66600
rect 9404 66580 9456 66600
rect 9456 66580 9458 66600
rect 9402 66544 9458 66580
rect 9494 65900 9496 65920
rect 9496 65900 9548 65920
rect 9548 65900 9550 65920
rect 9494 65864 9550 65900
rect 9115 65850 9171 65852
rect 9195 65850 9251 65852
rect 9275 65850 9331 65852
rect 9355 65850 9411 65852
rect 9115 65798 9161 65850
rect 9161 65798 9171 65850
rect 9195 65798 9225 65850
rect 9225 65798 9237 65850
rect 9237 65798 9251 65850
rect 9275 65798 9289 65850
rect 9289 65798 9301 65850
rect 9301 65798 9331 65850
rect 9355 65798 9365 65850
rect 9365 65798 9411 65850
rect 9115 65796 9171 65798
rect 9195 65796 9251 65798
rect 9275 65796 9331 65798
rect 9355 65796 9411 65798
rect 8758 64504 8814 64560
rect 8666 60152 8722 60208
rect 8574 55800 8630 55856
rect 8574 53488 8630 53544
rect 10046 66408 10102 66464
rect 10046 65456 10102 65512
rect 9115 64762 9171 64764
rect 9195 64762 9251 64764
rect 9275 64762 9331 64764
rect 9355 64762 9411 64764
rect 9115 64710 9161 64762
rect 9161 64710 9171 64762
rect 9195 64710 9225 64762
rect 9225 64710 9237 64762
rect 9237 64710 9251 64762
rect 9275 64710 9289 64762
rect 9289 64710 9301 64762
rect 9301 64710 9331 64762
rect 9355 64710 9365 64762
rect 9365 64710 9411 64762
rect 9115 64708 9171 64710
rect 9195 64708 9251 64710
rect 9275 64708 9331 64710
rect 9355 64708 9411 64710
rect 10046 64932 10102 64968
rect 10046 64912 10048 64932
rect 10048 64912 10100 64932
rect 10100 64912 10102 64932
rect 9586 63960 9642 64016
rect 9115 63674 9171 63676
rect 9195 63674 9251 63676
rect 9275 63674 9331 63676
rect 9355 63674 9411 63676
rect 9115 63622 9161 63674
rect 9161 63622 9171 63674
rect 9195 63622 9225 63674
rect 9225 63622 9237 63674
rect 9237 63622 9251 63674
rect 9275 63622 9289 63674
rect 9289 63622 9301 63674
rect 9301 63622 9331 63674
rect 9355 63622 9365 63674
rect 9365 63622 9411 63674
rect 9115 63620 9171 63622
rect 9195 63620 9251 63622
rect 9275 63620 9331 63622
rect 9355 63620 9411 63622
rect 9494 63552 9550 63608
rect 9115 62586 9171 62588
rect 9195 62586 9251 62588
rect 9275 62586 9331 62588
rect 9355 62586 9411 62588
rect 9115 62534 9161 62586
rect 9161 62534 9171 62586
rect 9195 62534 9225 62586
rect 9225 62534 9237 62586
rect 9237 62534 9251 62586
rect 9275 62534 9289 62586
rect 9289 62534 9301 62586
rect 9301 62534 9331 62586
rect 9355 62534 9365 62586
rect 9365 62534 9411 62586
rect 9115 62532 9171 62534
rect 9195 62532 9251 62534
rect 9275 62532 9331 62534
rect 9355 62532 9411 62534
rect 9310 61648 9366 61704
rect 9115 61498 9171 61500
rect 9195 61498 9251 61500
rect 9275 61498 9331 61500
rect 9355 61498 9411 61500
rect 9115 61446 9161 61498
rect 9161 61446 9171 61498
rect 9195 61446 9225 61498
rect 9225 61446 9237 61498
rect 9237 61446 9251 61498
rect 9275 61446 9289 61498
rect 9289 61446 9301 61498
rect 9301 61446 9331 61498
rect 9355 61446 9365 61498
rect 9365 61446 9411 61498
rect 9115 61444 9171 61446
rect 9195 61444 9251 61446
rect 9275 61444 9331 61446
rect 9355 61444 9411 61446
rect 9310 60716 9366 60752
rect 9310 60696 9312 60716
rect 9312 60696 9364 60716
rect 9364 60696 9366 60716
rect 9586 61104 9642 61160
rect 10138 63008 10194 63064
rect 10230 62600 10286 62656
rect 10138 62056 10194 62112
rect 9115 60410 9171 60412
rect 9195 60410 9251 60412
rect 9275 60410 9331 60412
rect 9355 60410 9411 60412
rect 9115 60358 9161 60410
rect 9161 60358 9171 60410
rect 9195 60358 9225 60410
rect 9225 60358 9237 60410
rect 9237 60358 9251 60410
rect 9275 60358 9289 60410
rect 9289 60358 9301 60410
rect 9301 60358 9331 60410
rect 9355 60358 9365 60410
rect 9365 60358 9411 60410
rect 9115 60356 9171 60358
rect 9195 60356 9251 60358
rect 9275 60356 9331 60358
rect 9355 60356 9411 60358
rect 9218 59744 9274 59800
rect 9115 59322 9171 59324
rect 9195 59322 9251 59324
rect 9275 59322 9331 59324
rect 9355 59322 9411 59324
rect 9115 59270 9161 59322
rect 9161 59270 9171 59322
rect 9195 59270 9225 59322
rect 9225 59270 9237 59322
rect 9237 59270 9251 59322
rect 9275 59270 9289 59322
rect 9289 59270 9301 59322
rect 9301 59270 9331 59322
rect 9355 59270 9365 59322
rect 9365 59270 9411 59322
rect 9115 59268 9171 59270
rect 9195 59268 9251 59270
rect 9275 59268 9331 59270
rect 9355 59268 9411 59270
rect 9115 58234 9171 58236
rect 9195 58234 9251 58236
rect 9275 58234 9331 58236
rect 9355 58234 9411 58236
rect 9115 58182 9161 58234
rect 9161 58182 9171 58234
rect 9195 58182 9225 58234
rect 9225 58182 9237 58234
rect 9237 58182 9251 58234
rect 9275 58182 9289 58234
rect 9289 58182 9301 58234
rect 9301 58182 9331 58234
rect 9355 58182 9365 58234
rect 9365 58182 9411 58234
rect 9115 58180 9171 58182
rect 9195 58180 9251 58182
rect 9275 58180 9331 58182
rect 9355 58180 9411 58182
rect 8942 51040 8998 51096
rect 8666 49836 8722 49872
rect 8666 49816 8668 49836
rect 8668 49816 8720 49836
rect 8720 49816 8722 49836
rect 9218 57296 9274 57352
rect 9115 57146 9171 57148
rect 9195 57146 9251 57148
rect 9275 57146 9331 57148
rect 9355 57146 9411 57148
rect 9115 57094 9161 57146
rect 9161 57094 9171 57146
rect 9195 57094 9225 57146
rect 9225 57094 9237 57146
rect 9237 57094 9251 57146
rect 9275 57094 9289 57146
rect 9289 57094 9301 57146
rect 9301 57094 9331 57146
rect 9355 57094 9365 57146
rect 9365 57094 9411 57146
rect 9115 57092 9171 57094
rect 9195 57092 9251 57094
rect 9275 57092 9331 57094
rect 9355 57092 9411 57094
rect 10046 59200 10102 59256
rect 9954 58792 10010 58848
rect 9954 57840 10010 57896
rect 9586 56480 9642 56536
rect 9115 56058 9171 56060
rect 9195 56058 9251 56060
rect 9275 56058 9331 56060
rect 9355 56058 9411 56060
rect 9115 56006 9161 56058
rect 9161 56006 9171 56058
rect 9195 56006 9225 56058
rect 9225 56006 9237 56058
rect 9237 56006 9251 56058
rect 9275 56006 9289 56058
rect 9289 56006 9301 56058
rect 9301 56006 9331 56058
rect 9355 56006 9365 56058
rect 9365 56006 9411 56058
rect 9115 56004 9171 56006
rect 9195 56004 9251 56006
rect 9275 56004 9331 56006
rect 9355 56004 9411 56006
rect 9115 54970 9171 54972
rect 9195 54970 9251 54972
rect 9275 54970 9331 54972
rect 9355 54970 9411 54972
rect 9115 54918 9161 54970
rect 9161 54918 9171 54970
rect 9195 54918 9225 54970
rect 9225 54918 9237 54970
rect 9237 54918 9251 54970
rect 9275 54918 9289 54970
rect 9289 54918 9301 54970
rect 9301 54918 9331 54970
rect 9355 54918 9365 54970
rect 9365 54918 9411 54970
rect 9115 54916 9171 54918
rect 9195 54916 9251 54918
rect 9275 54916 9331 54918
rect 9355 54916 9411 54918
rect 9862 55936 9918 55992
rect 9862 55528 9918 55584
rect 9862 54984 9918 55040
rect 9954 54596 10010 54632
rect 9954 54576 9956 54596
rect 9956 54576 10008 54596
rect 10008 54576 10010 54596
rect 9115 53882 9171 53884
rect 9195 53882 9251 53884
rect 9275 53882 9331 53884
rect 9355 53882 9411 53884
rect 9115 53830 9161 53882
rect 9161 53830 9171 53882
rect 9195 53830 9225 53882
rect 9225 53830 9237 53882
rect 9237 53830 9251 53882
rect 9275 53830 9289 53882
rect 9289 53830 9301 53882
rect 9301 53830 9331 53882
rect 9355 53830 9365 53882
rect 9365 53830 9411 53882
rect 9115 53828 9171 53830
rect 9195 53828 9251 53830
rect 9275 53828 9331 53830
rect 9355 53828 9411 53830
rect 9586 54032 9642 54088
rect 9494 53624 9550 53680
rect 9115 52794 9171 52796
rect 9195 52794 9251 52796
rect 9275 52794 9331 52796
rect 9355 52794 9411 52796
rect 9115 52742 9161 52794
rect 9161 52742 9171 52794
rect 9195 52742 9225 52794
rect 9225 52742 9237 52794
rect 9237 52742 9251 52794
rect 9275 52742 9289 52794
rect 9289 52742 9301 52794
rect 9301 52742 9331 52794
rect 9355 52742 9365 52794
rect 9365 52742 9411 52794
rect 9115 52740 9171 52742
rect 9195 52740 9251 52742
rect 9275 52740 9331 52742
rect 9355 52740 9411 52742
rect 9126 52128 9182 52184
rect 9494 51720 9550 51776
rect 9115 51706 9171 51708
rect 9195 51706 9251 51708
rect 9275 51706 9331 51708
rect 9355 51706 9411 51708
rect 9115 51654 9161 51706
rect 9161 51654 9171 51706
rect 9195 51654 9225 51706
rect 9225 51654 9237 51706
rect 9237 51654 9251 51706
rect 9275 51654 9289 51706
rect 9289 51654 9301 51706
rect 9301 51654 9331 51706
rect 9355 51654 9365 51706
rect 9365 51654 9411 51706
rect 9115 51652 9171 51654
rect 9195 51652 9251 51654
rect 9275 51652 9331 51654
rect 9355 51652 9411 51654
rect 10230 60596 10232 60616
rect 10232 60596 10284 60616
rect 10284 60596 10286 60616
rect 10230 60560 10286 60596
rect 10230 58248 10286 58304
rect 10322 56888 10378 56944
rect 9954 53080 10010 53136
rect 9862 52672 9918 52728
rect 9115 50618 9171 50620
rect 9195 50618 9251 50620
rect 9275 50618 9331 50620
rect 9355 50618 9411 50620
rect 9115 50566 9161 50618
rect 9161 50566 9171 50618
rect 9195 50566 9225 50618
rect 9225 50566 9237 50618
rect 9237 50566 9251 50618
rect 9275 50566 9289 50618
rect 9289 50566 9301 50618
rect 9301 50566 9331 50618
rect 9355 50566 9365 50618
rect 9365 50566 9411 50618
rect 9115 50564 9171 50566
rect 9195 50564 9251 50566
rect 9275 50564 9331 50566
rect 9355 50564 9411 50566
rect 9126 50360 9182 50416
rect 9115 49530 9171 49532
rect 9195 49530 9251 49532
rect 9275 49530 9331 49532
rect 9355 49530 9411 49532
rect 9115 49478 9161 49530
rect 9161 49478 9171 49530
rect 9195 49478 9225 49530
rect 9225 49478 9237 49530
rect 9237 49478 9251 49530
rect 9275 49478 9289 49530
rect 9289 49478 9301 49530
rect 9301 49478 9331 49530
rect 9355 49478 9365 49530
rect 9365 49478 9411 49530
rect 9115 49476 9171 49478
rect 9195 49476 9251 49478
rect 9275 49476 9331 49478
rect 9355 49476 9411 49478
rect 9862 50768 9918 50824
rect 9954 50088 10010 50144
rect 8850 48456 8906 48512
rect 8574 42744 8630 42800
rect 8482 41248 8538 41304
rect 8298 18536 8354 18592
rect 8574 40704 8630 40760
rect 8758 41520 8814 41576
rect 9115 48442 9171 48444
rect 9195 48442 9251 48444
rect 9275 48442 9331 48444
rect 9355 48442 9411 48444
rect 9115 48390 9161 48442
rect 9161 48390 9171 48442
rect 9195 48390 9225 48442
rect 9225 48390 9237 48442
rect 9237 48390 9251 48442
rect 9275 48390 9289 48442
rect 9289 48390 9301 48442
rect 9301 48390 9331 48442
rect 9355 48390 9365 48442
rect 9365 48390 9411 48442
rect 9115 48388 9171 48390
rect 9195 48388 9251 48390
rect 9275 48388 9331 48390
rect 9355 48388 9411 48390
rect 8666 39344 8722 39400
rect 8850 36080 8906 36136
rect 8850 35980 8852 36000
rect 8852 35980 8904 36000
rect 8904 35980 8906 36000
rect 8850 35944 8906 35980
rect 8850 35536 8906 35592
rect 8666 34448 8722 34504
rect 8574 33360 8630 33416
rect 8574 33088 8630 33144
rect 8390 18400 8446 18456
rect 8298 14728 8354 14784
rect 8390 13912 8446 13968
rect 7483 10906 7539 10908
rect 7563 10906 7619 10908
rect 7643 10906 7699 10908
rect 7723 10906 7779 10908
rect 7483 10854 7529 10906
rect 7529 10854 7539 10906
rect 7563 10854 7593 10906
rect 7593 10854 7605 10906
rect 7605 10854 7619 10906
rect 7643 10854 7657 10906
rect 7657 10854 7669 10906
rect 7669 10854 7699 10906
rect 7723 10854 7733 10906
rect 7733 10854 7779 10906
rect 7483 10852 7539 10854
rect 7563 10852 7619 10854
rect 7643 10852 7699 10854
rect 7723 10852 7779 10854
rect 8022 10512 8078 10568
rect 4219 5466 4275 5468
rect 4299 5466 4355 5468
rect 4379 5466 4435 5468
rect 4459 5466 4515 5468
rect 4219 5414 4265 5466
rect 4265 5414 4275 5466
rect 4299 5414 4329 5466
rect 4329 5414 4341 5466
rect 4341 5414 4355 5466
rect 4379 5414 4393 5466
rect 4393 5414 4405 5466
rect 4405 5414 4435 5466
rect 4459 5414 4469 5466
rect 4469 5414 4515 5466
rect 4219 5412 4275 5414
rect 4299 5412 4355 5414
rect 4379 5412 4435 5414
rect 4459 5412 4515 5414
rect 1582 4972 1584 4992
rect 1584 4972 1636 4992
rect 1636 4972 1638 4992
rect 1582 4936 1638 4972
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 4219 4378 4275 4380
rect 4299 4378 4355 4380
rect 4379 4378 4435 4380
rect 4459 4378 4515 4380
rect 4219 4326 4265 4378
rect 4265 4326 4275 4378
rect 4299 4326 4329 4378
rect 4329 4326 4341 4378
rect 4341 4326 4355 4378
rect 4379 4326 4393 4378
rect 4393 4326 4405 4378
rect 4405 4326 4435 4378
rect 4459 4326 4469 4378
rect 4469 4326 4515 4378
rect 4219 4324 4275 4326
rect 4299 4324 4355 4326
rect 4379 4324 4435 4326
rect 4459 4324 4515 4326
rect 1582 4256 1638 4312
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 1582 3576 1638 3632
rect 4219 3290 4275 3292
rect 4299 3290 4355 3292
rect 4379 3290 4435 3292
rect 4459 3290 4515 3292
rect 4219 3238 4265 3290
rect 4265 3238 4275 3290
rect 4299 3238 4329 3290
rect 4329 3238 4341 3290
rect 4341 3238 4355 3290
rect 4379 3238 4393 3290
rect 4393 3238 4405 3290
rect 4405 3238 4435 3290
rect 4459 3238 4469 3290
rect 4469 3238 4515 3290
rect 4219 3236 4275 3238
rect 4299 3236 4355 3238
rect 4379 3236 4435 3238
rect 4459 3236 4515 3238
rect 1582 2896 1638 2952
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 5851 4922 5907 4924
rect 5931 4922 5987 4924
rect 6011 4922 6067 4924
rect 6091 4922 6147 4924
rect 5851 4870 5897 4922
rect 5897 4870 5907 4922
rect 5931 4870 5961 4922
rect 5961 4870 5973 4922
rect 5973 4870 5987 4922
rect 6011 4870 6025 4922
rect 6025 4870 6037 4922
rect 6037 4870 6067 4922
rect 6091 4870 6101 4922
rect 6101 4870 6147 4922
rect 5851 4868 5907 4870
rect 5931 4868 5987 4870
rect 6011 4868 6067 4870
rect 6091 4868 6147 4870
rect 5851 3834 5907 3836
rect 5931 3834 5987 3836
rect 6011 3834 6067 3836
rect 6091 3834 6147 3836
rect 5851 3782 5897 3834
rect 5897 3782 5907 3834
rect 5931 3782 5961 3834
rect 5961 3782 5973 3834
rect 5973 3782 5987 3834
rect 6011 3782 6025 3834
rect 6025 3782 6037 3834
rect 6037 3782 6067 3834
rect 6091 3782 6101 3834
rect 6101 3782 6147 3834
rect 5851 3780 5907 3782
rect 5931 3780 5987 3782
rect 6011 3780 6067 3782
rect 6091 3780 6147 3782
rect 5851 2746 5907 2748
rect 5931 2746 5987 2748
rect 6011 2746 6067 2748
rect 6091 2746 6147 2748
rect 5851 2694 5897 2746
rect 5897 2694 5907 2746
rect 5931 2694 5961 2746
rect 5961 2694 5973 2746
rect 5973 2694 5987 2746
rect 6011 2694 6025 2746
rect 6025 2694 6037 2746
rect 6037 2694 6067 2746
rect 6091 2694 6101 2746
rect 6101 2694 6147 2746
rect 5851 2692 5907 2694
rect 5931 2692 5987 2694
rect 6011 2692 6067 2694
rect 6091 2692 6147 2694
rect 7483 9818 7539 9820
rect 7563 9818 7619 9820
rect 7643 9818 7699 9820
rect 7723 9818 7779 9820
rect 7483 9766 7529 9818
rect 7529 9766 7539 9818
rect 7563 9766 7593 9818
rect 7593 9766 7605 9818
rect 7605 9766 7619 9818
rect 7643 9766 7657 9818
rect 7657 9766 7669 9818
rect 7669 9766 7699 9818
rect 7723 9766 7733 9818
rect 7733 9766 7779 9818
rect 7483 9764 7539 9766
rect 7563 9764 7619 9766
rect 7643 9764 7699 9766
rect 7723 9764 7779 9766
rect 7838 9424 7894 9480
rect 7483 8730 7539 8732
rect 7563 8730 7619 8732
rect 7643 8730 7699 8732
rect 7723 8730 7779 8732
rect 7483 8678 7529 8730
rect 7529 8678 7539 8730
rect 7563 8678 7593 8730
rect 7593 8678 7605 8730
rect 7605 8678 7619 8730
rect 7643 8678 7657 8730
rect 7657 8678 7669 8730
rect 7669 8678 7699 8730
rect 7723 8678 7733 8730
rect 7733 8678 7779 8730
rect 7483 8676 7539 8678
rect 7563 8676 7619 8678
rect 7643 8676 7699 8678
rect 7723 8676 7779 8678
rect 7483 7642 7539 7644
rect 7563 7642 7619 7644
rect 7643 7642 7699 7644
rect 7723 7642 7779 7644
rect 7483 7590 7529 7642
rect 7529 7590 7539 7642
rect 7563 7590 7593 7642
rect 7593 7590 7605 7642
rect 7605 7590 7619 7642
rect 7643 7590 7657 7642
rect 7657 7590 7669 7642
rect 7669 7590 7699 7642
rect 7723 7590 7733 7642
rect 7733 7590 7779 7642
rect 7483 7588 7539 7590
rect 7563 7588 7619 7590
rect 7643 7588 7699 7590
rect 7723 7588 7779 7590
rect 7483 6554 7539 6556
rect 7563 6554 7619 6556
rect 7643 6554 7699 6556
rect 7723 6554 7779 6556
rect 7483 6502 7529 6554
rect 7529 6502 7539 6554
rect 7563 6502 7593 6554
rect 7593 6502 7605 6554
rect 7605 6502 7619 6554
rect 7643 6502 7657 6554
rect 7657 6502 7669 6554
rect 7669 6502 7699 6554
rect 7723 6502 7733 6554
rect 7733 6502 7779 6554
rect 7483 6500 7539 6502
rect 7563 6500 7619 6502
rect 7643 6500 7699 6502
rect 7723 6500 7779 6502
rect 7483 5466 7539 5468
rect 7563 5466 7619 5468
rect 7643 5466 7699 5468
rect 7723 5466 7779 5468
rect 7483 5414 7529 5466
rect 7529 5414 7539 5466
rect 7563 5414 7593 5466
rect 7593 5414 7605 5466
rect 7605 5414 7619 5466
rect 7643 5414 7657 5466
rect 7657 5414 7669 5466
rect 7669 5414 7699 5466
rect 7723 5414 7733 5466
rect 7733 5414 7779 5466
rect 7483 5412 7539 5414
rect 7563 5412 7619 5414
rect 7643 5412 7699 5414
rect 7723 5412 7779 5414
rect 7483 4378 7539 4380
rect 7563 4378 7619 4380
rect 7643 4378 7699 4380
rect 7723 4378 7779 4380
rect 7483 4326 7529 4378
rect 7529 4326 7539 4378
rect 7563 4326 7593 4378
rect 7593 4326 7605 4378
rect 7605 4326 7619 4378
rect 7643 4326 7657 4378
rect 7657 4326 7669 4378
rect 7669 4326 7699 4378
rect 7723 4326 7733 4378
rect 7733 4326 7779 4378
rect 7483 4324 7539 4326
rect 7563 4324 7619 4326
rect 7643 4324 7699 4326
rect 7723 4324 7779 4326
rect 8114 5072 8170 5128
rect 8114 3476 8116 3496
rect 8116 3476 8168 3496
rect 8168 3476 8170 3496
rect 8114 3440 8170 3476
rect 7483 3290 7539 3292
rect 7563 3290 7619 3292
rect 7643 3290 7699 3292
rect 7723 3290 7779 3292
rect 7483 3238 7529 3290
rect 7529 3238 7539 3290
rect 7563 3238 7593 3290
rect 7593 3238 7605 3290
rect 7605 3238 7619 3290
rect 7643 3238 7657 3290
rect 7657 3238 7669 3290
rect 7669 3238 7699 3290
rect 7723 3238 7733 3290
rect 7733 3238 7779 3290
rect 7483 3236 7539 3238
rect 7563 3236 7619 3238
rect 7643 3236 7699 3238
rect 7723 3236 7779 3238
rect 7838 2916 7894 2952
rect 7838 2896 7840 2916
rect 7840 2896 7892 2916
rect 7892 2896 7894 2916
rect 2318 2252 2320 2272
rect 2320 2252 2372 2272
rect 2372 2252 2374 2272
rect 1398 1536 1454 1592
rect 2318 2216 2374 2252
rect 1582 856 1638 912
rect 4219 2202 4275 2204
rect 4299 2202 4355 2204
rect 4379 2202 4435 2204
rect 4459 2202 4515 2204
rect 4219 2150 4265 2202
rect 4265 2150 4275 2202
rect 4299 2150 4329 2202
rect 4329 2150 4341 2202
rect 4341 2150 4355 2202
rect 4379 2150 4393 2202
rect 4393 2150 4405 2202
rect 4405 2150 4435 2202
rect 4459 2150 4469 2202
rect 4469 2150 4515 2202
rect 4219 2148 4275 2150
rect 4299 2148 4355 2150
rect 4379 2148 4435 2150
rect 4459 2148 4515 2150
rect 7483 2202 7539 2204
rect 7563 2202 7619 2204
rect 7643 2202 7699 2204
rect 7723 2202 7779 2204
rect 7483 2150 7529 2202
rect 7529 2150 7539 2202
rect 7563 2150 7593 2202
rect 7593 2150 7605 2202
rect 7605 2150 7619 2202
rect 7643 2150 7657 2202
rect 7657 2150 7669 2202
rect 7669 2150 7699 2202
rect 7723 2150 7733 2202
rect 7733 2150 7779 2202
rect 7483 2148 7539 2150
rect 7563 2148 7619 2150
rect 7643 2148 7699 2150
rect 7723 2148 7779 2150
rect 7930 1536 7986 1592
rect 2870 312 2926 368
rect 8390 11056 8446 11112
rect 8850 31864 8906 31920
rect 9218 47640 9274 47696
rect 9126 47504 9182 47560
rect 9494 47368 9550 47424
rect 9115 47354 9171 47356
rect 9195 47354 9251 47356
rect 9275 47354 9331 47356
rect 9355 47354 9411 47356
rect 9115 47302 9161 47354
rect 9161 47302 9171 47354
rect 9195 47302 9225 47354
rect 9225 47302 9237 47354
rect 9237 47302 9251 47354
rect 9275 47302 9289 47354
rect 9289 47302 9301 47354
rect 9301 47302 9331 47354
rect 9355 47302 9365 47354
rect 9365 47302 9411 47354
rect 9115 47300 9171 47302
rect 9195 47300 9251 47302
rect 9275 47300 9331 47302
rect 9355 47300 9411 47302
rect 9586 46552 9642 46608
rect 9494 46452 9496 46472
rect 9496 46452 9548 46472
rect 9548 46452 9550 46472
rect 9494 46416 9550 46452
rect 9115 46266 9171 46268
rect 9195 46266 9251 46268
rect 9275 46266 9331 46268
rect 9355 46266 9411 46268
rect 9115 46214 9161 46266
rect 9161 46214 9171 46266
rect 9195 46214 9225 46266
rect 9225 46214 9237 46266
rect 9237 46214 9251 46266
rect 9275 46214 9289 46266
rect 9289 46214 9301 46266
rect 9301 46214 9331 46266
rect 9355 46214 9365 46266
rect 9365 46214 9411 46266
rect 9115 46212 9171 46214
rect 9195 46212 9251 46214
rect 9275 46212 9331 46214
rect 9355 46212 9411 46214
rect 9494 46144 9550 46200
rect 9115 45178 9171 45180
rect 9195 45178 9251 45180
rect 9275 45178 9331 45180
rect 9355 45178 9411 45180
rect 9115 45126 9161 45178
rect 9161 45126 9171 45178
rect 9195 45126 9225 45178
rect 9225 45126 9237 45178
rect 9237 45126 9251 45178
rect 9275 45126 9289 45178
rect 9289 45126 9301 45178
rect 9301 45126 9331 45178
rect 9355 45126 9365 45178
rect 9365 45126 9411 45178
rect 9115 45124 9171 45126
rect 9195 45124 9251 45126
rect 9275 45124 9331 45126
rect 9355 45124 9411 45126
rect 9402 44820 9404 44840
rect 9404 44820 9456 44840
rect 9456 44820 9458 44840
rect 9402 44784 9458 44820
rect 9402 44512 9458 44568
rect 9218 44240 9274 44296
rect 9115 44090 9171 44092
rect 9195 44090 9251 44092
rect 9275 44090 9331 44092
rect 9355 44090 9411 44092
rect 9115 44038 9161 44090
rect 9161 44038 9171 44090
rect 9195 44038 9225 44090
rect 9225 44038 9237 44090
rect 9237 44038 9251 44090
rect 9275 44038 9289 44090
rect 9289 44038 9301 44090
rect 9301 44038 9331 44090
rect 9355 44038 9365 44090
rect 9365 44038 9411 44090
rect 9115 44036 9171 44038
rect 9195 44036 9251 44038
rect 9275 44036 9331 44038
rect 9355 44036 9411 44038
rect 9126 43696 9182 43752
rect 9115 43002 9171 43004
rect 9195 43002 9251 43004
rect 9275 43002 9331 43004
rect 9355 43002 9411 43004
rect 9115 42950 9161 43002
rect 9161 42950 9171 43002
rect 9195 42950 9225 43002
rect 9225 42950 9237 43002
rect 9237 42950 9251 43002
rect 9275 42950 9289 43002
rect 9289 42950 9301 43002
rect 9301 42950 9331 43002
rect 9355 42950 9365 43002
rect 9365 42950 9411 43002
rect 9115 42948 9171 42950
rect 9195 42948 9251 42950
rect 9275 42948 9331 42950
rect 9355 42948 9411 42950
rect 9126 42220 9182 42256
rect 9126 42200 9128 42220
rect 9128 42200 9180 42220
rect 9180 42200 9182 42220
rect 9115 41914 9171 41916
rect 9195 41914 9251 41916
rect 9275 41914 9331 41916
rect 9355 41914 9411 41916
rect 9115 41862 9161 41914
rect 9161 41862 9171 41914
rect 9195 41862 9225 41914
rect 9225 41862 9237 41914
rect 9237 41862 9251 41914
rect 9275 41862 9289 41914
rect 9289 41862 9301 41914
rect 9301 41862 9331 41914
rect 9355 41862 9365 41914
rect 9365 41862 9411 41914
rect 9115 41860 9171 41862
rect 9195 41860 9251 41862
rect 9275 41860 9331 41862
rect 9355 41860 9411 41862
rect 9586 43832 9642 43888
rect 9115 40826 9171 40828
rect 9195 40826 9251 40828
rect 9275 40826 9331 40828
rect 9355 40826 9411 40828
rect 9115 40774 9161 40826
rect 9161 40774 9171 40826
rect 9195 40774 9225 40826
rect 9225 40774 9237 40826
rect 9237 40774 9251 40826
rect 9275 40774 9289 40826
rect 9289 40774 9301 40826
rect 9301 40774 9331 40826
rect 9355 40774 9365 40826
rect 9365 40774 9411 40826
rect 9115 40772 9171 40774
rect 9195 40772 9251 40774
rect 9275 40772 9331 40774
rect 9355 40772 9411 40774
rect 9310 39888 9366 39944
rect 9115 39738 9171 39740
rect 9195 39738 9251 39740
rect 9275 39738 9331 39740
rect 9355 39738 9411 39740
rect 9115 39686 9161 39738
rect 9161 39686 9171 39738
rect 9195 39686 9225 39738
rect 9225 39686 9237 39738
rect 9237 39686 9251 39738
rect 9275 39686 9289 39738
rect 9289 39686 9301 39738
rect 9301 39686 9331 39738
rect 9355 39686 9365 39738
rect 9365 39686 9411 39738
rect 9115 39684 9171 39686
rect 9195 39684 9251 39686
rect 9275 39684 9331 39686
rect 9355 39684 9411 39686
rect 9402 39480 9458 39536
rect 9126 38820 9182 38856
rect 9126 38800 9128 38820
rect 9128 38800 9180 38820
rect 9180 38800 9182 38820
rect 9115 38650 9171 38652
rect 9195 38650 9251 38652
rect 9275 38650 9331 38652
rect 9355 38650 9411 38652
rect 9115 38598 9161 38650
rect 9161 38598 9171 38650
rect 9195 38598 9225 38650
rect 9225 38598 9237 38650
rect 9237 38598 9251 38650
rect 9275 38598 9289 38650
rect 9289 38598 9301 38650
rect 9301 38598 9331 38650
rect 9355 38598 9365 38650
rect 9365 38598 9411 38650
rect 9115 38596 9171 38598
rect 9195 38596 9251 38598
rect 9275 38596 9331 38598
rect 9355 38596 9411 38598
rect 9126 38256 9182 38312
rect 9218 38156 9220 38176
rect 9220 38156 9272 38176
rect 9272 38156 9274 38176
rect 9218 38120 9274 38156
rect 9954 46316 9956 46336
rect 9956 46316 10008 46336
rect 10008 46316 10010 46336
rect 9954 46280 10010 46316
rect 10230 46280 10286 46336
rect 9310 37848 9366 37904
rect 9862 44376 9918 44432
rect 9862 43152 9918 43208
rect 9954 41792 10010 41848
rect 9954 41248 10010 41304
rect 9954 40840 10010 40896
rect 10138 42608 10194 42664
rect 10138 42336 10194 42392
rect 10138 42064 10194 42120
rect 9862 39616 9918 39672
rect 10138 40432 10194 40488
rect 9770 38528 9826 38584
rect 9115 37562 9171 37564
rect 9195 37562 9251 37564
rect 9275 37562 9331 37564
rect 9355 37562 9411 37564
rect 9115 37510 9161 37562
rect 9161 37510 9171 37562
rect 9195 37510 9225 37562
rect 9225 37510 9237 37562
rect 9237 37510 9251 37562
rect 9275 37510 9289 37562
rect 9289 37510 9301 37562
rect 9301 37510 9331 37562
rect 9355 37510 9365 37562
rect 9365 37510 9411 37562
rect 9115 37508 9171 37510
rect 9195 37508 9251 37510
rect 9275 37508 9331 37510
rect 9355 37508 9411 37510
rect 9586 37440 9642 37496
rect 9115 36474 9171 36476
rect 9195 36474 9251 36476
rect 9275 36474 9331 36476
rect 9355 36474 9411 36476
rect 9115 36422 9161 36474
rect 9161 36422 9171 36474
rect 9195 36422 9225 36474
rect 9225 36422 9237 36474
rect 9237 36422 9251 36474
rect 9275 36422 9289 36474
rect 9289 36422 9301 36474
rect 9301 36422 9331 36474
rect 9355 36422 9365 36474
rect 9365 36422 9411 36474
rect 9115 36420 9171 36422
rect 9195 36420 9251 36422
rect 9275 36420 9331 36422
rect 9355 36420 9411 36422
rect 9402 36236 9458 36272
rect 9402 36216 9404 36236
rect 9404 36216 9456 36236
rect 9456 36216 9458 36236
rect 9115 35386 9171 35388
rect 9195 35386 9251 35388
rect 9275 35386 9331 35388
rect 9355 35386 9411 35388
rect 9115 35334 9161 35386
rect 9161 35334 9171 35386
rect 9195 35334 9225 35386
rect 9225 35334 9237 35386
rect 9237 35334 9251 35386
rect 9275 35334 9289 35386
rect 9289 35334 9301 35386
rect 9301 35334 9331 35386
rect 9355 35334 9365 35386
rect 9365 35334 9411 35386
rect 9115 35332 9171 35334
rect 9195 35332 9251 35334
rect 9275 35332 9331 35334
rect 9355 35332 9411 35334
rect 9115 34298 9171 34300
rect 9195 34298 9251 34300
rect 9275 34298 9331 34300
rect 9355 34298 9411 34300
rect 9115 34246 9161 34298
rect 9161 34246 9171 34298
rect 9195 34246 9225 34298
rect 9225 34246 9237 34298
rect 9237 34246 9251 34298
rect 9275 34246 9289 34298
rect 9289 34246 9301 34298
rect 9301 34246 9331 34298
rect 9355 34246 9365 34298
rect 9365 34246 9411 34298
rect 9115 34244 9171 34246
rect 9195 34244 9251 34246
rect 9275 34244 9331 34246
rect 9355 34244 9411 34246
rect 9310 33804 9312 33824
rect 9312 33804 9364 33824
rect 9364 33804 9366 33824
rect 9310 33768 9366 33804
rect 9115 33210 9171 33212
rect 9195 33210 9251 33212
rect 9275 33210 9331 33212
rect 9355 33210 9411 33212
rect 9115 33158 9161 33210
rect 9161 33158 9171 33210
rect 9195 33158 9225 33210
rect 9225 33158 9237 33210
rect 9237 33158 9251 33210
rect 9275 33158 9289 33210
rect 9289 33158 9301 33210
rect 9301 33158 9331 33210
rect 9355 33158 9365 33210
rect 9365 33158 9411 33210
rect 9115 33156 9171 33158
rect 9195 33156 9251 33158
rect 9275 33156 9331 33158
rect 9355 33156 9411 33158
rect 10046 38936 10102 38992
rect 9586 33496 9642 33552
rect 9586 33224 9642 33280
rect 9218 32272 9274 32328
rect 9115 32122 9171 32124
rect 9195 32122 9251 32124
rect 9275 32122 9331 32124
rect 9355 32122 9411 32124
rect 9115 32070 9161 32122
rect 9161 32070 9171 32122
rect 9195 32070 9225 32122
rect 9225 32070 9237 32122
rect 9237 32070 9251 32122
rect 9275 32070 9289 32122
rect 9289 32070 9301 32122
rect 9301 32070 9331 32122
rect 9355 32070 9365 32122
rect 9365 32070 9411 32122
rect 9115 32068 9171 32070
rect 9195 32068 9251 32070
rect 9275 32068 9331 32070
rect 9355 32068 9411 32070
rect 9115 31034 9171 31036
rect 9195 31034 9251 31036
rect 9275 31034 9331 31036
rect 9355 31034 9411 31036
rect 9115 30982 9161 31034
rect 9161 30982 9171 31034
rect 9195 30982 9225 31034
rect 9225 30982 9237 31034
rect 9237 30982 9251 31034
rect 9275 30982 9289 31034
rect 9289 30982 9301 31034
rect 9301 30982 9331 31034
rect 9355 30982 9365 31034
rect 9365 30982 9411 31034
rect 9115 30980 9171 30982
rect 9195 30980 9251 30982
rect 9275 30980 9331 30982
rect 9355 30980 9411 30982
rect 9115 29946 9171 29948
rect 9195 29946 9251 29948
rect 9275 29946 9331 29948
rect 9355 29946 9411 29948
rect 9115 29894 9161 29946
rect 9161 29894 9171 29946
rect 9195 29894 9225 29946
rect 9225 29894 9237 29946
rect 9237 29894 9251 29946
rect 9275 29894 9289 29946
rect 9289 29894 9301 29946
rect 9301 29894 9331 29946
rect 9355 29894 9365 29946
rect 9365 29894 9411 29946
rect 9115 29892 9171 29894
rect 9195 29892 9251 29894
rect 9275 29892 9331 29894
rect 9355 29892 9411 29894
rect 9310 29452 9312 29472
rect 9312 29452 9364 29472
rect 9364 29452 9366 29472
rect 9310 29416 9366 29452
rect 9126 29028 9182 29064
rect 9126 29008 9128 29028
rect 9128 29008 9180 29028
rect 9180 29008 9182 29028
rect 9115 28858 9171 28860
rect 9195 28858 9251 28860
rect 9275 28858 9331 28860
rect 9355 28858 9411 28860
rect 9115 28806 9161 28858
rect 9161 28806 9171 28858
rect 9195 28806 9225 28858
rect 9225 28806 9237 28858
rect 9237 28806 9251 28858
rect 9275 28806 9289 28858
rect 9289 28806 9301 28858
rect 9301 28806 9331 28858
rect 9355 28806 9365 28858
rect 9365 28806 9411 28858
rect 9115 28804 9171 28806
rect 9195 28804 9251 28806
rect 9275 28804 9331 28806
rect 9355 28804 9411 28806
rect 9310 28056 9366 28112
rect 9115 27770 9171 27772
rect 9195 27770 9251 27772
rect 9275 27770 9331 27772
rect 9355 27770 9411 27772
rect 9115 27718 9161 27770
rect 9161 27718 9171 27770
rect 9195 27718 9225 27770
rect 9225 27718 9237 27770
rect 9237 27718 9251 27770
rect 9275 27718 9289 27770
rect 9289 27718 9301 27770
rect 9301 27718 9331 27770
rect 9355 27718 9365 27770
rect 9365 27718 9411 27770
rect 9115 27716 9171 27718
rect 9195 27716 9251 27718
rect 9275 27716 9331 27718
rect 9355 27716 9411 27718
rect 8758 22888 8814 22944
rect 9115 26682 9171 26684
rect 9195 26682 9251 26684
rect 9275 26682 9331 26684
rect 9355 26682 9411 26684
rect 9115 26630 9161 26682
rect 9161 26630 9171 26682
rect 9195 26630 9225 26682
rect 9225 26630 9237 26682
rect 9237 26630 9251 26682
rect 9275 26630 9289 26682
rect 9289 26630 9301 26682
rect 9301 26630 9331 26682
rect 9355 26630 9365 26682
rect 9365 26630 9411 26682
rect 9115 26628 9171 26630
rect 9195 26628 9251 26630
rect 9275 26628 9331 26630
rect 9355 26628 9411 26630
rect 9494 25644 9496 25664
rect 9496 25644 9548 25664
rect 9548 25644 9550 25664
rect 9494 25608 9550 25644
rect 9115 25594 9171 25596
rect 9195 25594 9251 25596
rect 9275 25594 9331 25596
rect 9355 25594 9411 25596
rect 9115 25542 9161 25594
rect 9161 25542 9171 25594
rect 9195 25542 9225 25594
rect 9225 25542 9237 25594
rect 9237 25542 9251 25594
rect 9275 25542 9289 25594
rect 9289 25542 9301 25594
rect 9301 25542 9331 25594
rect 9355 25542 9365 25594
rect 9365 25542 9411 25594
rect 9115 25540 9171 25542
rect 9195 25540 9251 25542
rect 9275 25540 9331 25542
rect 9355 25540 9411 25542
rect 9115 24506 9171 24508
rect 9195 24506 9251 24508
rect 9275 24506 9331 24508
rect 9355 24506 9411 24508
rect 9115 24454 9161 24506
rect 9161 24454 9171 24506
rect 9195 24454 9225 24506
rect 9225 24454 9237 24506
rect 9237 24454 9251 24506
rect 9275 24454 9289 24506
rect 9289 24454 9301 24506
rect 9301 24454 9331 24506
rect 9355 24454 9365 24506
rect 9365 24454 9411 24506
rect 9115 24452 9171 24454
rect 9195 24452 9251 24454
rect 9275 24452 9331 24454
rect 9355 24452 9411 24454
rect 9494 24248 9550 24304
rect 9126 23704 9182 23760
rect 9115 23418 9171 23420
rect 9195 23418 9251 23420
rect 9275 23418 9331 23420
rect 9355 23418 9411 23420
rect 9115 23366 9161 23418
rect 9161 23366 9171 23418
rect 9195 23366 9225 23418
rect 9225 23366 9237 23418
rect 9237 23366 9251 23418
rect 9275 23366 9289 23418
rect 9289 23366 9301 23418
rect 9301 23366 9331 23418
rect 9355 23366 9365 23418
rect 9365 23366 9411 23418
rect 9115 23364 9171 23366
rect 9195 23364 9251 23366
rect 9275 23364 9331 23366
rect 9355 23364 9411 23366
rect 9115 22330 9171 22332
rect 9195 22330 9251 22332
rect 9275 22330 9331 22332
rect 9355 22330 9411 22332
rect 9115 22278 9161 22330
rect 9161 22278 9171 22330
rect 9195 22278 9225 22330
rect 9225 22278 9237 22330
rect 9237 22278 9251 22330
rect 9275 22278 9289 22330
rect 9289 22278 9301 22330
rect 9301 22278 9331 22330
rect 9355 22278 9365 22330
rect 9365 22278 9411 22330
rect 9115 22276 9171 22278
rect 9195 22276 9251 22278
rect 9275 22276 9331 22278
rect 9355 22276 9411 22278
rect 9310 21392 9366 21448
rect 9115 21242 9171 21244
rect 9195 21242 9251 21244
rect 9275 21242 9331 21244
rect 9355 21242 9411 21244
rect 9115 21190 9161 21242
rect 9161 21190 9171 21242
rect 9195 21190 9225 21242
rect 9225 21190 9237 21242
rect 9237 21190 9251 21242
rect 9275 21190 9289 21242
rect 9289 21190 9301 21242
rect 9301 21190 9331 21242
rect 9355 21190 9365 21242
rect 9365 21190 9411 21242
rect 9115 21188 9171 21190
rect 9195 21188 9251 21190
rect 9275 21188 9331 21190
rect 9355 21188 9411 21190
rect 10138 34584 10194 34640
rect 10046 34176 10102 34232
rect 10046 32816 10102 32872
rect 9862 29300 9918 29336
rect 9862 29280 9864 29300
rect 9864 29280 9916 29300
rect 9916 29280 9918 29300
rect 10138 30504 10194 30560
rect 10046 30368 10102 30424
rect 10046 29996 10048 30016
rect 10048 29996 10100 30016
rect 10100 29996 10102 30016
rect 10046 29960 10102 29996
rect 10046 29708 10102 29744
rect 10046 29688 10048 29708
rect 10048 29688 10100 29708
rect 10100 29688 10102 29708
rect 10138 29572 10194 29608
rect 10138 29552 10140 29572
rect 10140 29552 10192 29572
rect 10192 29552 10194 29572
rect 10046 28464 10102 28520
rect 10230 28212 10286 28248
rect 10230 28192 10232 28212
rect 10232 28192 10284 28212
rect 10284 28192 10286 28212
rect 10138 27512 10194 27568
rect 10046 27104 10102 27160
rect 10138 26560 10194 26616
rect 10046 26152 10102 26208
rect 9494 20984 9550 21040
rect 9310 20440 9366 20496
rect 9115 20154 9171 20156
rect 9195 20154 9251 20156
rect 9275 20154 9331 20156
rect 9355 20154 9411 20156
rect 9115 20102 9161 20154
rect 9161 20102 9171 20154
rect 9195 20102 9225 20154
rect 9225 20102 9237 20154
rect 9237 20102 9251 20154
rect 9275 20102 9289 20154
rect 9289 20102 9301 20154
rect 9301 20102 9331 20154
rect 9355 20102 9365 20154
rect 9365 20102 9411 20154
rect 9115 20100 9171 20102
rect 9195 20100 9251 20102
rect 9275 20100 9331 20102
rect 9355 20100 9411 20102
rect 8666 17584 8722 17640
rect 9115 19066 9171 19068
rect 9195 19066 9251 19068
rect 9275 19066 9331 19068
rect 9355 19066 9411 19068
rect 9115 19014 9161 19066
rect 9161 19014 9171 19066
rect 9195 19014 9225 19066
rect 9225 19014 9237 19066
rect 9237 19014 9251 19066
rect 9275 19014 9289 19066
rect 9289 19014 9301 19066
rect 9301 19014 9331 19066
rect 9355 19014 9365 19066
rect 9365 19014 9411 19066
rect 9115 19012 9171 19014
rect 9195 19012 9251 19014
rect 9275 19012 9331 19014
rect 9355 19012 9411 19014
rect 9115 17978 9171 17980
rect 9195 17978 9251 17980
rect 9275 17978 9331 17980
rect 9355 17978 9411 17980
rect 9115 17926 9161 17978
rect 9161 17926 9171 17978
rect 9195 17926 9225 17978
rect 9225 17926 9237 17978
rect 9237 17926 9251 17978
rect 9275 17926 9289 17978
rect 9289 17926 9301 17978
rect 9301 17926 9331 17978
rect 9355 17926 9365 17978
rect 9365 17926 9411 17978
rect 9115 17924 9171 17926
rect 9195 17924 9251 17926
rect 9275 17924 9331 17926
rect 9355 17924 9411 17926
rect 9115 16890 9171 16892
rect 9195 16890 9251 16892
rect 9275 16890 9331 16892
rect 9355 16890 9411 16892
rect 9115 16838 9161 16890
rect 9161 16838 9171 16890
rect 9195 16838 9225 16890
rect 9225 16838 9237 16890
rect 9237 16838 9251 16890
rect 9275 16838 9289 16890
rect 9289 16838 9301 16890
rect 9301 16838 9331 16890
rect 9355 16838 9365 16890
rect 9365 16838 9411 16890
rect 9115 16836 9171 16838
rect 9195 16836 9251 16838
rect 9275 16836 9331 16838
rect 9355 16836 9411 16838
rect 9115 15802 9171 15804
rect 9195 15802 9251 15804
rect 9275 15802 9331 15804
rect 9355 15802 9411 15804
rect 9115 15750 9161 15802
rect 9161 15750 9171 15802
rect 9195 15750 9225 15802
rect 9225 15750 9237 15802
rect 9237 15750 9251 15802
rect 9275 15750 9289 15802
rect 9289 15750 9301 15802
rect 9301 15750 9331 15802
rect 9355 15750 9365 15802
rect 9365 15750 9411 15802
rect 9115 15748 9171 15750
rect 9195 15748 9251 15750
rect 9275 15748 9331 15750
rect 9355 15748 9411 15750
rect 8850 15156 8906 15192
rect 8850 15136 8852 15156
rect 8852 15136 8904 15156
rect 8904 15136 8906 15156
rect 9115 14714 9171 14716
rect 9195 14714 9251 14716
rect 9275 14714 9331 14716
rect 9355 14714 9411 14716
rect 9115 14662 9161 14714
rect 9161 14662 9171 14714
rect 9195 14662 9225 14714
rect 9225 14662 9237 14714
rect 9237 14662 9251 14714
rect 9275 14662 9289 14714
rect 9289 14662 9301 14714
rect 9301 14662 9331 14714
rect 9355 14662 9365 14714
rect 9365 14662 9411 14714
rect 9115 14660 9171 14662
rect 9195 14660 9251 14662
rect 9275 14660 9331 14662
rect 9355 14660 9411 14662
rect 8942 7248 8998 7304
rect 9115 13626 9171 13628
rect 9195 13626 9251 13628
rect 9275 13626 9331 13628
rect 9355 13626 9411 13628
rect 9115 13574 9161 13626
rect 9161 13574 9171 13626
rect 9195 13574 9225 13626
rect 9225 13574 9237 13626
rect 9237 13574 9251 13626
rect 9275 13574 9289 13626
rect 9289 13574 9301 13626
rect 9301 13574 9331 13626
rect 9355 13574 9365 13626
rect 9365 13574 9411 13626
rect 9115 13572 9171 13574
rect 9195 13572 9251 13574
rect 9275 13572 9331 13574
rect 9355 13572 9411 13574
rect 9862 24656 9918 24712
rect 9954 23296 10010 23352
rect 10690 52400 10746 52456
rect 10966 53216 11022 53272
rect 10966 51448 11022 51504
rect 10782 51040 10838 51096
rect 10966 51348 10968 51368
rect 10968 51348 11020 51368
rect 11020 51348 11022 51368
rect 10966 51312 11022 51348
rect 10690 41656 10746 41712
rect 10966 49308 10968 49328
rect 10968 49308 11020 49328
rect 11020 49308 11022 49328
rect 10966 49272 11022 49308
rect 10782 41384 10838 41440
rect 11702 56208 11758 56264
rect 11794 54304 11850 54360
rect 11334 50496 11390 50552
rect 11426 43424 11482 43480
rect 11518 42472 11574 42528
rect 10782 40160 10838 40216
rect 10598 36760 10654 36816
rect 10506 36624 10562 36680
rect 10414 33360 10470 33416
rect 10598 33108 10654 33144
rect 10598 33088 10600 33108
rect 10600 33088 10652 33108
rect 10652 33088 10654 33108
rect 10506 32000 10562 32056
rect 10414 30912 10470 30968
rect 10414 30796 10470 30832
rect 10414 30776 10416 30796
rect 10416 30776 10468 30796
rect 10468 30776 10470 30796
rect 10046 22344 10102 22400
rect 9586 19080 9642 19136
rect 10598 31184 10654 31240
rect 11610 38664 11666 38720
rect 11610 36796 11612 36816
rect 11612 36796 11664 36816
rect 11664 36796 11666 36816
rect 11610 36760 11666 36796
rect 11886 39616 11942 39672
rect 10874 31592 10930 31648
rect 10966 25236 10968 25256
rect 10968 25236 11020 25256
rect 11020 25236 11022 25256
rect 10966 25200 11022 25236
rect 10966 22208 11022 22264
rect 11886 32544 11942 32600
rect 11886 29708 11942 29744
rect 11886 29688 11888 29708
rect 11888 29688 11940 29708
rect 11940 29688 11942 29708
rect 11058 16260 11060 16280
rect 11060 16260 11112 16280
rect 11112 16260 11114 16280
rect 11058 16224 11114 16260
rect 9115 12538 9171 12540
rect 9195 12538 9251 12540
rect 9275 12538 9331 12540
rect 9355 12538 9411 12540
rect 9115 12486 9161 12538
rect 9161 12486 9171 12538
rect 9195 12486 9225 12538
rect 9225 12486 9237 12538
rect 9237 12486 9251 12538
rect 9275 12486 9289 12538
rect 9289 12486 9301 12538
rect 9301 12486 9331 12538
rect 9355 12486 9365 12538
rect 9365 12486 9411 12538
rect 9115 12484 9171 12486
rect 9195 12484 9251 12486
rect 9275 12484 9331 12486
rect 9355 12484 9411 12486
rect 9115 11450 9171 11452
rect 9195 11450 9251 11452
rect 9275 11450 9331 11452
rect 9355 11450 9411 11452
rect 9115 11398 9161 11450
rect 9161 11398 9171 11450
rect 9195 11398 9225 11450
rect 9225 11398 9237 11450
rect 9237 11398 9251 11450
rect 9275 11398 9289 11450
rect 9289 11398 9301 11450
rect 9301 11398 9331 11450
rect 9355 11398 9365 11450
rect 9365 11398 9411 11450
rect 9115 11396 9171 11398
rect 9195 11396 9251 11398
rect 9275 11396 9331 11398
rect 9355 11396 9411 11398
rect 9115 10362 9171 10364
rect 9195 10362 9251 10364
rect 9275 10362 9331 10364
rect 9355 10362 9411 10364
rect 9115 10310 9161 10362
rect 9161 10310 9171 10362
rect 9195 10310 9225 10362
rect 9225 10310 9237 10362
rect 9237 10310 9251 10362
rect 9275 10310 9289 10362
rect 9289 10310 9301 10362
rect 9301 10310 9331 10362
rect 9355 10310 9365 10362
rect 9365 10310 9411 10362
rect 9115 10308 9171 10310
rect 9195 10308 9251 10310
rect 9275 10308 9331 10310
rect 9355 10308 9411 10310
rect 9218 10104 9274 10160
rect 9115 9274 9171 9276
rect 9195 9274 9251 9276
rect 9275 9274 9331 9276
rect 9355 9274 9411 9276
rect 9115 9222 9161 9274
rect 9161 9222 9171 9274
rect 9195 9222 9225 9274
rect 9225 9222 9237 9274
rect 9237 9222 9251 9274
rect 9275 9222 9289 9274
rect 9289 9222 9301 9274
rect 9301 9222 9331 9274
rect 9355 9222 9365 9274
rect 9365 9222 9411 9274
rect 9115 9220 9171 9222
rect 9195 9220 9251 9222
rect 9275 9220 9331 9222
rect 9355 9220 9411 9222
rect 9126 8608 9182 8664
rect 9115 8186 9171 8188
rect 9195 8186 9251 8188
rect 9275 8186 9331 8188
rect 9355 8186 9411 8188
rect 9115 8134 9161 8186
rect 9161 8134 9171 8186
rect 9195 8134 9225 8186
rect 9225 8134 9237 8186
rect 9237 8134 9251 8186
rect 9275 8134 9289 8186
rect 9289 8134 9301 8186
rect 9301 8134 9331 8186
rect 9355 8134 9365 8186
rect 9365 8134 9411 8186
rect 9115 8132 9171 8134
rect 9195 8132 9251 8134
rect 9275 8132 9331 8134
rect 9355 8132 9411 8134
rect 9115 7098 9171 7100
rect 9195 7098 9251 7100
rect 9275 7098 9331 7100
rect 9355 7098 9411 7100
rect 9115 7046 9161 7098
rect 9161 7046 9171 7098
rect 9195 7046 9225 7098
rect 9225 7046 9237 7098
rect 9237 7046 9251 7098
rect 9275 7046 9289 7098
rect 9289 7046 9301 7098
rect 9301 7046 9331 7098
rect 9355 7046 9365 7098
rect 9365 7046 9411 7098
rect 9115 7044 9171 7046
rect 9195 7044 9251 7046
rect 9275 7044 9331 7046
rect 9355 7044 9411 7046
rect 8942 4392 8998 4448
rect 9115 6010 9171 6012
rect 9195 6010 9251 6012
rect 9275 6010 9331 6012
rect 9355 6010 9411 6012
rect 9115 5958 9161 6010
rect 9161 5958 9171 6010
rect 9195 5958 9225 6010
rect 9225 5958 9237 6010
rect 9237 5958 9251 6010
rect 9275 5958 9289 6010
rect 9289 5958 9301 6010
rect 9301 5958 9331 6010
rect 9355 5958 9365 6010
rect 9365 5958 9411 6010
rect 9115 5956 9171 5958
rect 9195 5956 9251 5958
rect 9275 5956 9331 5958
rect 9355 5956 9411 5958
rect 9115 4922 9171 4924
rect 9195 4922 9251 4924
rect 9275 4922 9331 4924
rect 9355 4922 9411 4924
rect 9115 4870 9161 4922
rect 9161 4870 9171 4922
rect 9195 4870 9225 4922
rect 9225 4870 9237 4922
rect 9237 4870 9251 4922
rect 9275 4870 9289 4922
rect 9289 4870 9301 4922
rect 9301 4870 9331 4922
rect 9355 4870 9365 4922
rect 9365 4870 9411 4922
rect 9115 4868 9171 4870
rect 9195 4868 9251 4870
rect 9275 4868 9331 4870
rect 9355 4868 9411 4870
rect 10414 10104 10470 10160
rect 9770 9580 9826 9616
rect 9770 9560 9772 9580
rect 9772 9560 9824 9580
rect 9824 9560 9826 9580
rect 9862 8200 9918 8256
rect 10230 7656 10286 7712
rect 9770 6296 9826 6352
rect 10966 6740 10968 6760
rect 10968 6740 11020 6760
rect 11020 6740 11022 6760
rect 10966 6704 11022 6740
rect 9126 3984 9182 4040
rect 9115 3834 9171 3836
rect 9195 3834 9251 3836
rect 9275 3834 9331 3836
rect 9355 3834 9411 3836
rect 9115 3782 9161 3834
rect 9161 3782 9171 3834
rect 9195 3782 9225 3834
rect 9225 3782 9237 3834
rect 9237 3782 9251 3834
rect 9275 3782 9289 3834
rect 9289 3782 9301 3834
rect 9301 3782 9331 3834
rect 9355 3782 9365 3834
rect 9365 3782 9411 3834
rect 9115 3780 9171 3782
rect 9195 3780 9251 3782
rect 9275 3780 9331 3782
rect 9355 3780 9411 3782
rect 9115 2746 9171 2748
rect 9195 2746 9251 2748
rect 9275 2746 9331 2748
rect 9355 2746 9411 2748
rect 9115 2694 9161 2746
rect 9161 2694 9171 2746
rect 9195 2694 9225 2746
rect 9225 2694 9237 2746
rect 9237 2694 9251 2746
rect 9275 2694 9289 2746
rect 9289 2694 9301 2746
rect 9301 2694 9331 2746
rect 9355 2694 9365 2746
rect 9365 2694 9411 2746
rect 9115 2692 9171 2694
rect 9195 2692 9251 2694
rect 9275 2692 9331 2694
rect 9355 2692 9411 2694
rect 9586 2488 9642 2544
rect 9494 1944 9550 2000
rect 9310 992 9366 1048
rect 8206 584 8262 640
rect 8114 176 8170 232
<< metal3 >>
rect 0 79658 800 79688
rect 3233 79658 3299 79661
rect 0 79656 3299 79658
rect 0 79600 3238 79656
rect 3294 79600 3299 79656
rect 0 79598 3299 79600
rect 0 79568 800 79598
rect 3233 79595 3299 79598
rect 7557 79658 7623 79661
rect 11200 79658 12000 79688
rect 7557 79656 12000 79658
rect 7557 79600 7562 79656
rect 7618 79600 12000 79656
rect 7557 79598 12000 79600
rect 7557 79595 7623 79598
rect 11200 79568 12000 79598
rect 8569 79250 8635 79253
rect 11200 79250 12000 79280
rect 8569 79248 12000 79250
rect 8569 79192 8574 79248
rect 8630 79192 12000 79248
rect 8569 79190 12000 79192
rect 8569 79187 8635 79190
rect 11200 79160 12000 79190
rect 0 78978 800 79008
rect 1393 78978 1459 78981
rect 0 78976 1459 78978
rect 0 78920 1398 78976
rect 1454 78920 1459 78976
rect 0 78918 1459 78920
rect 0 78888 800 78918
rect 1393 78915 1459 78918
rect 9489 78706 9555 78709
rect 11200 78706 12000 78736
rect 9489 78704 12000 78706
rect 9489 78648 9494 78704
rect 9550 78648 12000 78704
rect 9489 78646 12000 78648
rect 9489 78643 9555 78646
rect 11200 78616 12000 78646
rect 0 78298 800 78328
rect 2957 78298 3023 78301
rect 0 78296 3023 78298
rect 0 78240 2962 78296
rect 3018 78240 3023 78296
rect 0 78238 3023 78240
rect 0 78208 800 78238
rect 2957 78235 3023 78238
rect 8201 78298 8267 78301
rect 11200 78298 12000 78328
rect 8201 78296 12000 78298
rect 8201 78240 8206 78296
rect 8262 78240 12000 78296
rect 8201 78238 12000 78240
rect 8201 78235 8267 78238
rect 11200 78208 12000 78238
rect 2576 77824 2896 77825
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 77759 2896 77760
rect 5839 77824 6159 77825
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 77759 6159 77760
rect 9103 77824 9423 77825
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 77759 9423 77760
rect 9581 77754 9647 77757
rect 11200 77754 12000 77784
rect 9581 77752 12000 77754
rect 9581 77696 9586 77752
rect 9642 77696 12000 77752
rect 9581 77694 12000 77696
rect 9581 77691 9647 77694
rect 11200 77664 12000 77694
rect 0 77618 800 77648
rect 2865 77618 2931 77621
rect 0 77616 2931 77618
rect 0 77560 2870 77616
rect 2926 77560 2931 77616
rect 0 77558 2931 77560
rect 0 77528 800 77558
rect 2865 77555 2931 77558
rect 9305 77346 9371 77349
rect 11200 77346 12000 77376
rect 9305 77344 12000 77346
rect 9305 77288 9310 77344
rect 9366 77288 12000 77344
rect 9305 77286 12000 77288
rect 9305 77283 9371 77286
rect 4207 77280 4527 77281
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 77215 4527 77216
rect 7471 77280 7791 77281
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 11200 77256 12000 77286
rect 7471 77215 7791 77216
rect 0 76938 800 76968
rect 1577 76938 1643 76941
rect 0 76936 1643 76938
rect 0 76880 1582 76936
rect 1638 76880 1643 76936
rect 0 76878 1643 76880
rect 0 76848 800 76878
rect 1577 76875 1643 76878
rect 10133 76802 10199 76805
rect 11200 76802 12000 76832
rect 10133 76800 12000 76802
rect 10133 76744 10138 76800
rect 10194 76744 12000 76800
rect 10133 76742 12000 76744
rect 10133 76739 10199 76742
rect 2576 76736 2896 76737
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 76671 2896 76672
rect 5839 76736 6159 76737
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 76671 6159 76672
rect 9103 76736 9423 76737
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 11200 76712 12000 76742
rect 9103 76671 9423 76672
rect 10041 76394 10107 76397
rect 11200 76394 12000 76424
rect 10041 76392 12000 76394
rect 10041 76336 10046 76392
rect 10102 76336 12000 76392
rect 10041 76334 12000 76336
rect 10041 76331 10107 76334
rect 11200 76304 12000 76334
rect 0 76258 800 76288
rect 1577 76258 1643 76261
rect 0 76256 1643 76258
rect 0 76200 1582 76256
rect 1638 76200 1643 76256
rect 0 76198 1643 76200
rect 0 76168 800 76198
rect 1577 76195 1643 76198
rect 4207 76192 4527 76193
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 76127 4527 76128
rect 7471 76192 7791 76193
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 76127 7791 76128
rect 9305 75850 9371 75853
rect 11200 75850 12000 75880
rect 9305 75848 12000 75850
rect 9305 75792 9310 75848
rect 9366 75792 12000 75848
rect 9305 75790 12000 75792
rect 9305 75787 9371 75790
rect 11200 75760 12000 75790
rect 2576 75648 2896 75649
rect 0 75578 800 75608
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 75583 2896 75584
rect 5839 75648 6159 75649
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 75583 6159 75584
rect 9103 75648 9423 75649
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 9103 75583 9423 75584
rect 1393 75578 1459 75581
rect 0 75576 1459 75578
rect 0 75520 1398 75576
rect 1454 75520 1459 75576
rect 0 75518 1459 75520
rect 0 75488 800 75518
rect 1393 75515 1459 75518
rect 10041 75442 10107 75445
rect 11200 75442 12000 75472
rect 10041 75440 12000 75442
rect 10041 75384 10046 75440
rect 10102 75384 12000 75440
rect 10041 75382 12000 75384
rect 10041 75379 10107 75382
rect 11200 75352 12000 75382
rect 4207 75104 4527 75105
rect 0 75034 800 75064
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 75039 4527 75040
rect 7471 75104 7791 75105
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 75039 7791 75040
rect 1853 75034 1919 75037
rect 0 75032 1919 75034
rect 0 74976 1858 75032
rect 1914 74976 1919 75032
rect 0 74974 1919 74976
rect 0 74944 800 74974
rect 1853 74971 1919 74974
rect 10961 74898 11027 74901
rect 11200 74898 12000 74928
rect 10961 74896 12000 74898
rect 10961 74840 10966 74896
rect 11022 74840 12000 74896
rect 10961 74838 12000 74840
rect 10961 74835 11027 74838
rect 11200 74808 12000 74838
rect 2576 74560 2896 74561
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 74495 2896 74496
rect 5839 74560 6159 74561
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 74495 6159 74496
rect 9103 74560 9423 74561
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 74495 9423 74496
rect 10133 74490 10199 74493
rect 11200 74490 12000 74520
rect 10133 74488 12000 74490
rect 10133 74432 10138 74488
rect 10194 74432 12000 74488
rect 10133 74430 12000 74432
rect 10133 74427 10199 74430
rect 11200 74400 12000 74430
rect 0 74354 800 74384
rect 2221 74354 2287 74357
rect 0 74352 2287 74354
rect 0 74296 2226 74352
rect 2282 74296 2287 74352
rect 0 74294 2287 74296
rect 0 74264 800 74294
rect 2221 74291 2287 74294
rect 4207 74016 4527 74017
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 73951 4527 73952
rect 7471 74016 7791 74017
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 73951 7791 73952
rect 10041 73946 10107 73949
rect 11200 73946 12000 73976
rect 10041 73944 12000 73946
rect 10041 73888 10046 73944
rect 10102 73888 12000 73944
rect 10041 73886 12000 73888
rect 10041 73883 10107 73886
rect 11200 73856 12000 73886
rect 0 73674 800 73704
rect 1577 73674 1643 73677
rect 0 73672 1643 73674
rect 0 73616 1582 73672
rect 1638 73616 1643 73672
rect 0 73614 1643 73616
rect 0 73584 800 73614
rect 1577 73611 1643 73614
rect 9489 73538 9555 73541
rect 11200 73538 12000 73568
rect 9489 73536 12000 73538
rect 9489 73480 9494 73536
rect 9550 73480 12000 73536
rect 9489 73478 12000 73480
rect 9489 73475 9555 73478
rect 2576 73472 2896 73473
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 73407 2896 73408
rect 5839 73472 6159 73473
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 73407 6159 73408
rect 9103 73472 9423 73473
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 11200 73448 12000 73478
rect 9103 73407 9423 73408
rect 0 72994 800 73024
rect 2865 72994 2931 72997
rect 0 72992 2931 72994
rect 0 72936 2870 72992
rect 2926 72936 2931 72992
rect 0 72934 2931 72936
rect 0 72904 800 72934
rect 2865 72931 2931 72934
rect 10041 72994 10107 72997
rect 11200 72994 12000 73024
rect 10041 72992 12000 72994
rect 10041 72936 10046 72992
rect 10102 72936 12000 72992
rect 10041 72934 12000 72936
rect 10041 72931 10107 72934
rect 4207 72928 4527 72929
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 72863 4527 72864
rect 7471 72928 7791 72929
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 11200 72904 12000 72934
rect 7471 72863 7791 72864
rect 9305 72586 9371 72589
rect 11200 72586 12000 72616
rect 9305 72584 12000 72586
rect 9305 72528 9310 72584
rect 9366 72528 12000 72584
rect 9305 72526 12000 72528
rect 9305 72523 9371 72526
rect 11200 72496 12000 72526
rect 2576 72384 2896 72385
rect 0 72314 800 72344
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 72319 2896 72320
rect 5839 72384 6159 72385
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 72319 6159 72320
rect 9103 72384 9423 72385
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 72319 9423 72320
rect 2221 72314 2287 72317
rect 0 72312 2287 72314
rect 0 72256 2226 72312
rect 2282 72256 2287 72312
rect 0 72254 2287 72256
rect 0 72224 800 72254
rect 2221 72251 2287 72254
rect 9305 72042 9371 72045
rect 11200 72042 12000 72072
rect 9305 72040 12000 72042
rect 9305 71984 9310 72040
rect 9366 71984 12000 72040
rect 9305 71982 12000 71984
rect 9305 71979 9371 71982
rect 11200 71952 12000 71982
rect 8569 71908 8635 71909
rect 8518 71906 8524 71908
rect 8478 71846 8524 71906
rect 8588 71904 8635 71908
rect 8630 71848 8635 71904
rect 8518 71844 8524 71846
rect 8588 71844 8635 71848
rect 8569 71843 8635 71844
rect 4207 71840 4527 71841
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 71775 4527 71776
rect 7471 71840 7791 71841
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 71775 7791 71776
rect 0 71634 800 71664
rect 1577 71634 1643 71637
rect 0 71632 1643 71634
rect 0 71576 1582 71632
rect 1638 71576 1643 71632
rect 0 71574 1643 71576
rect 0 71544 800 71574
rect 1577 71571 1643 71574
rect 10133 71634 10199 71637
rect 11200 71634 12000 71664
rect 10133 71632 12000 71634
rect 10133 71576 10138 71632
rect 10194 71576 12000 71632
rect 10133 71574 12000 71576
rect 10133 71571 10199 71574
rect 11200 71544 12000 71574
rect 2576 71296 2896 71297
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 71231 2896 71232
rect 5839 71296 6159 71297
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 71231 6159 71232
rect 9103 71296 9423 71297
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 71231 9423 71232
rect 10041 71090 10107 71093
rect 11200 71090 12000 71120
rect 10041 71088 12000 71090
rect 10041 71032 10046 71088
rect 10102 71032 12000 71088
rect 10041 71030 12000 71032
rect 10041 71027 10107 71030
rect 11200 71000 12000 71030
rect 0 70954 800 70984
rect 1393 70954 1459 70957
rect 0 70952 1459 70954
rect 0 70896 1398 70952
rect 1454 70896 1459 70952
rect 0 70894 1459 70896
rect 0 70864 800 70894
rect 1393 70891 1459 70894
rect 4207 70752 4527 70753
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 70687 4527 70688
rect 7471 70752 7791 70753
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 70687 7791 70688
rect 10133 70682 10199 70685
rect 11200 70682 12000 70712
rect 10133 70680 12000 70682
rect 10133 70624 10138 70680
rect 10194 70624 12000 70680
rect 10133 70622 12000 70624
rect 10133 70619 10199 70622
rect 11200 70592 12000 70622
rect 1485 70546 1551 70549
rect 798 70544 1551 70546
rect 798 70488 1490 70544
rect 1546 70488 1551 70544
rect 798 70486 1551 70488
rect 798 70440 858 70486
rect 1485 70483 1551 70486
rect 0 70350 858 70440
rect 0 70320 800 70350
rect 2576 70208 2896 70209
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2576 70143 2896 70144
rect 5839 70208 6159 70209
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 70143 6159 70144
rect 9103 70208 9423 70209
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 70143 9423 70144
rect 10041 70138 10107 70141
rect 11200 70138 12000 70168
rect 10041 70136 12000 70138
rect 10041 70080 10046 70136
rect 10102 70080 12000 70136
rect 10041 70078 12000 70080
rect 10041 70075 10107 70078
rect 11200 70048 12000 70078
rect 0 69730 800 69760
rect 3969 69730 4035 69733
rect 0 69728 4035 69730
rect 0 69672 3974 69728
rect 4030 69672 4035 69728
rect 0 69670 4035 69672
rect 0 69640 800 69670
rect 3969 69667 4035 69670
rect 10409 69730 10475 69733
rect 11200 69730 12000 69760
rect 10409 69728 12000 69730
rect 10409 69672 10414 69728
rect 10470 69672 12000 69728
rect 10409 69670 12000 69672
rect 10409 69667 10475 69670
rect 4207 69664 4527 69665
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 69599 4527 69600
rect 7471 69664 7791 69665
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 11200 69640 12000 69670
rect 7471 69599 7791 69600
rect 2865 69322 2931 69325
rect 1534 69320 2931 69322
rect 1534 69264 2870 69320
rect 2926 69264 2931 69320
rect 1534 69262 2931 69264
rect 0 69050 800 69080
rect 1534 69050 1594 69262
rect 2865 69259 2931 69262
rect 8886 69260 8892 69324
rect 8956 69322 8962 69324
rect 9029 69322 9095 69325
rect 8956 69320 9095 69322
rect 8956 69264 9034 69320
rect 9090 69264 9095 69320
rect 8956 69262 9095 69264
rect 8956 69260 8962 69262
rect 9029 69259 9095 69262
rect 9489 69186 9555 69189
rect 11200 69186 12000 69216
rect 9489 69184 12000 69186
rect 9489 69128 9494 69184
rect 9550 69128 12000 69184
rect 9489 69126 12000 69128
rect 9489 69123 9555 69126
rect 2576 69120 2896 69121
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 69055 2896 69056
rect 5839 69120 6159 69121
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 69055 6159 69056
rect 9103 69120 9423 69121
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 11200 69096 12000 69126
rect 9103 69055 9423 69056
rect 0 68990 1594 69050
rect 0 68960 800 68990
rect 8201 68778 8267 68781
rect 11200 68778 12000 68808
rect 8201 68776 12000 68778
rect 8201 68720 8206 68776
rect 8262 68720 12000 68776
rect 8201 68718 12000 68720
rect 8201 68715 8267 68718
rect 11200 68688 12000 68718
rect 4207 68576 4527 68577
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 68511 4527 68512
rect 7471 68576 7791 68577
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 68511 7791 68512
rect 0 68370 800 68400
rect 1577 68370 1643 68373
rect 0 68368 1643 68370
rect 0 68312 1582 68368
rect 1638 68312 1643 68368
rect 0 68310 1643 68312
rect 0 68280 800 68310
rect 1577 68307 1643 68310
rect 9581 68370 9647 68373
rect 11200 68370 12000 68400
rect 9581 68368 12000 68370
rect 9581 68312 9586 68368
rect 9642 68312 12000 68368
rect 9581 68310 12000 68312
rect 9581 68307 9647 68310
rect 11200 68280 12000 68310
rect 2576 68032 2896 68033
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 67967 2896 67968
rect 5839 68032 6159 68033
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 67967 6159 67968
rect 9103 68032 9423 68033
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 67967 9423 67968
rect 8753 67826 8819 67829
rect 11200 67826 12000 67856
rect 8753 67824 12000 67826
rect 8753 67768 8758 67824
rect 8814 67768 12000 67824
rect 8753 67766 12000 67768
rect 8753 67763 8819 67766
rect 11200 67736 12000 67766
rect 0 67690 800 67720
rect 1393 67690 1459 67693
rect 0 67688 1459 67690
rect 0 67632 1398 67688
rect 1454 67632 1459 67688
rect 0 67630 1459 67632
rect 0 67600 800 67630
rect 1393 67627 1459 67630
rect 8702 67628 8708 67692
rect 8772 67690 8778 67692
rect 9397 67690 9463 67693
rect 8772 67688 9463 67690
rect 8772 67632 9402 67688
rect 9458 67632 9463 67688
rect 8772 67630 9463 67632
rect 8772 67628 8778 67630
rect 9397 67627 9463 67630
rect 4207 67488 4527 67489
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 67423 4527 67424
rect 7471 67488 7791 67489
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 67423 7791 67424
rect 8293 67418 8359 67421
rect 11200 67418 12000 67448
rect 8293 67416 12000 67418
rect 8293 67360 8298 67416
rect 8354 67360 12000 67416
rect 8293 67358 12000 67360
rect 8293 67355 8359 67358
rect 11200 67328 12000 67358
rect 0 67010 800 67040
rect 1485 67010 1551 67013
rect 0 67008 1551 67010
rect 0 66952 1490 67008
rect 1546 66952 1551 67008
rect 0 66950 1551 66952
rect 0 66920 800 66950
rect 1485 66947 1551 66950
rect 2576 66944 2896 66945
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 66879 2896 66880
rect 5839 66944 6159 66945
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 66879 6159 66880
rect 9103 66944 9423 66945
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 66879 9423 66880
rect 9489 66874 9555 66877
rect 11200 66874 12000 66904
rect 9489 66872 12000 66874
rect 9489 66816 9494 66872
rect 9550 66816 12000 66872
rect 9489 66814 12000 66816
rect 9489 66811 9555 66814
rect 11200 66784 12000 66814
rect 9397 66602 9463 66605
rect 9622 66602 9628 66604
rect 9397 66600 9628 66602
rect 9397 66544 9402 66600
rect 9458 66544 9628 66600
rect 9397 66542 9628 66544
rect 9397 66539 9463 66542
rect 9622 66540 9628 66542
rect 9692 66540 9698 66604
rect 10041 66466 10107 66469
rect 11200 66466 12000 66496
rect 10041 66464 12000 66466
rect 10041 66408 10046 66464
rect 10102 66408 12000 66464
rect 10041 66406 12000 66408
rect 10041 66403 10107 66406
rect 4207 66400 4527 66401
rect 0 66330 800 66360
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 66335 4527 66336
rect 7471 66400 7791 66401
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 11200 66376 12000 66406
rect 7471 66335 7791 66336
rect 2957 66330 3023 66333
rect 0 66328 3023 66330
rect 0 66272 2962 66328
rect 3018 66272 3023 66328
rect 0 66270 3023 66272
rect 0 66240 800 66270
rect 2957 66267 3023 66270
rect 8293 66332 8359 66333
rect 8293 66328 8340 66332
rect 8404 66330 8410 66332
rect 8293 66272 8298 66328
rect 8293 66268 8340 66272
rect 8404 66270 8450 66330
rect 8404 66268 8410 66270
rect 8293 66267 8359 66268
rect 9489 65922 9555 65925
rect 11200 65922 12000 65952
rect 9489 65920 12000 65922
rect 9489 65864 9494 65920
rect 9550 65864 12000 65920
rect 9489 65862 12000 65864
rect 9489 65859 9555 65862
rect 2576 65856 2896 65857
rect 0 65786 800 65816
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 65791 2896 65792
rect 5839 65856 6159 65857
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 65791 6159 65792
rect 9103 65856 9423 65857
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 11200 65832 12000 65862
rect 9103 65791 9423 65792
rect 1577 65786 1643 65789
rect 0 65784 1643 65786
rect 0 65728 1582 65784
rect 1638 65728 1643 65784
rect 0 65726 1643 65728
rect 0 65696 800 65726
rect 1577 65723 1643 65726
rect 10041 65514 10107 65517
rect 11200 65514 12000 65544
rect 10041 65512 12000 65514
rect 10041 65456 10046 65512
rect 10102 65456 12000 65512
rect 10041 65454 12000 65456
rect 10041 65451 10107 65454
rect 11200 65424 12000 65454
rect 4207 65312 4527 65313
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 65247 4527 65248
rect 7471 65312 7791 65313
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 65247 7791 65248
rect 0 65106 800 65136
rect 2221 65106 2287 65109
rect 0 65104 2287 65106
rect 0 65048 2226 65104
rect 2282 65048 2287 65104
rect 0 65046 2287 65048
rect 0 65016 800 65046
rect 2221 65043 2287 65046
rect 10041 64970 10107 64973
rect 11200 64970 12000 65000
rect 10041 64968 12000 64970
rect 10041 64912 10046 64968
rect 10102 64912 12000 64968
rect 10041 64910 12000 64912
rect 10041 64907 10107 64910
rect 11200 64880 12000 64910
rect 2576 64768 2896 64769
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 64703 2896 64704
rect 5839 64768 6159 64769
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 64703 6159 64704
rect 9103 64768 9423 64769
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 64703 9423 64704
rect 8753 64562 8819 64565
rect 11200 64562 12000 64592
rect 8753 64560 12000 64562
rect 8753 64504 8758 64560
rect 8814 64504 12000 64560
rect 8753 64502 12000 64504
rect 8753 64499 8819 64502
rect 11200 64472 12000 64502
rect 0 64426 800 64456
rect 1853 64426 1919 64429
rect 0 64424 1919 64426
rect 0 64368 1858 64424
rect 1914 64368 1919 64424
rect 0 64366 1919 64368
rect 0 64336 800 64366
rect 1853 64363 1919 64366
rect 4207 64224 4527 64225
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 64159 4527 64160
rect 7471 64224 7791 64225
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 64159 7791 64160
rect 9581 64018 9647 64021
rect 11200 64018 12000 64048
rect 9581 64016 12000 64018
rect 9581 63960 9586 64016
rect 9642 63960 12000 64016
rect 9581 63958 12000 63960
rect 9581 63955 9647 63958
rect 11200 63928 12000 63958
rect 0 63746 800 63776
rect 1393 63746 1459 63749
rect 0 63744 1459 63746
rect 0 63688 1398 63744
rect 1454 63688 1459 63744
rect 0 63686 1459 63688
rect 0 63656 800 63686
rect 1393 63683 1459 63686
rect 2576 63680 2896 63681
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 63615 2896 63616
rect 5839 63680 6159 63681
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 63615 6159 63616
rect 9103 63680 9423 63681
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 63615 9423 63616
rect 9489 63610 9555 63613
rect 11200 63610 12000 63640
rect 9489 63608 12000 63610
rect 9489 63552 9494 63608
rect 9550 63552 12000 63608
rect 9489 63550 12000 63552
rect 9489 63547 9555 63550
rect 11200 63520 12000 63550
rect 4207 63136 4527 63137
rect 0 63066 800 63096
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 63071 4527 63072
rect 7471 63136 7791 63137
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 63071 7791 63072
rect 1025 63066 1091 63069
rect 0 63064 1091 63066
rect 0 63008 1030 63064
rect 1086 63008 1091 63064
rect 0 63006 1091 63008
rect 0 62976 800 63006
rect 1025 63003 1091 63006
rect 10133 63066 10199 63069
rect 11200 63066 12000 63096
rect 10133 63064 12000 63066
rect 10133 63008 10138 63064
rect 10194 63008 12000 63064
rect 10133 63006 12000 63008
rect 10133 63003 10199 63006
rect 11200 62976 12000 63006
rect 2589 62794 2655 62797
rect 3550 62794 3556 62796
rect 2589 62792 3556 62794
rect 2589 62736 2594 62792
rect 2650 62736 3556 62792
rect 2589 62734 3556 62736
rect 2589 62731 2655 62734
rect 3550 62732 3556 62734
rect 3620 62732 3626 62796
rect 10225 62658 10291 62661
rect 11200 62658 12000 62688
rect 10225 62656 12000 62658
rect 10225 62600 10230 62656
rect 10286 62600 12000 62656
rect 10225 62598 12000 62600
rect 10225 62595 10291 62598
rect 2576 62592 2896 62593
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 62527 2896 62528
rect 5839 62592 6159 62593
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 62527 6159 62528
rect 9103 62592 9423 62593
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 11200 62568 12000 62598
rect 9103 62527 9423 62528
rect 0 62386 800 62416
rect 1393 62386 1459 62389
rect 0 62384 1459 62386
rect 0 62328 1398 62384
rect 1454 62328 1459 62384
rect 0 62326 1459 62328
rect 0 62296 800 62326
rect 1393 62323 1459 62326
rect 10133 62114 10199 62117
rect 11200 62114 12000 62144
rect 10133 62112 12000 62114
rect 10133 62056 10138 62112
rect 10194 62056 12000 62112
rect 10133 62054 12000 62056
rect 10133 62051 10199 62054
rect 4207 62048 4527 62049
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 61983 4527 61984
rect 7471 62048 7791 62049
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 11200 62024 12000 62054
rect 7471 61983 7791 61984
rect 0 61706 800 61736
rect 1853 61706 1919 61709
rect 0 61704 1919 61706
rect 0 61648 1858 61704
rect 1914 61648 1919 61704
rect 0 61646 1919 61648
rect 0 61616 800 61646
rect 1853 61643 1919 61646
rect 9305 61706 9371 61709
rect 11200 61706 12000 61736
rect 9305 61704 12000 61706
rect 9305 61648 9310 61704
rect 9366 61648 12000 61704
rect 9305 61646 12000 61648
rect 9305 61643 9371 61646
rect 11200 61616 12000 61646
rect 2576 61504 2896 61505
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2576 61439 2896 61440
rect 5839 61504 6159 61505
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 61439 6159 61440
rect 9103 61504 9423 61505
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 61439 9423 61440
rect 8150 61236 8156 61300
rect 8220 61298 8226 61300
rect 9622 61298 9628 61300
rect 8220 61238 9628 61298
rect 8220 61236 8226 61238
rect 9622 61236 9628 61238
rect 9692 61236 9698 61300
rect 0 61162 800 61192
rect 1393 61162 1459 61165
rect 0 61160 1459 61162
rect 0 61104 1398 61160
rect 1454 61104 1459 61160
rect 0 61102 1459 61104
rect 0 61072 800 61102
rect 1393 61099 1459 61102
rect 9581 61162 9647 61165
rect 11200 61162 12000 61192
rect 9581 61160 12000 61162
rect 9581 61104 9586 61160
rect 9642 61104 12000 61160
rect 9581 61102 12000 61104
rect 9581 61099 9647 61102
rect 11200 61072 12000 61102
rect 8293 61026 8359 61029
rect 8158 61024 8359 61026
rect 8158 60968 8298 61024
rect 8354 60968 8359 61024
rect 8158 60966 8359 60968
rect 4207 60960 4527 60961
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 60895 4527 60896
rect 7471 60960 7791 60961
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 60895 7791 60896
rect 8158 60757 8218 60966
rect 8293 60963 8359 60966
rect 8109 60752 8218 60757
rect 8109 60696 8114 60752
rect 8170 60696 8218 60752
rect 8109 60694 8218 60696
rect 9305 60754 9371 60757
rect 11200 60754 12000 60784
rect 9305 60752 12000 60754
rect 9305 60696 9310 60752
rect 9366 60696 12000 60752
rect 9305 60694 12000 60696
rect 8109 60691 8175 60694
rect 9305 60691 9371 60694
rect 11200 60664 12000 60694
rect 2773 60618 2839 60621
rect 10225 60620 10291 60621
rect 1350 60616 2839 60618
rect 1350 60560 2778 60616
rect 2834 60560 2839 60616
rect 1350 60558 2839 60560
rect 0 60482 800 60512
rect 1350 60482 1410 60558
rect 2773 60555 2839 60558
rect 8150 60556 8156 60620
rect 8220 60618 8226 60620
rect 9622 60618 9628 60620
rect 8220 60558 9628 60618
rect 8220 60556 8226 60558
rect 9622 60556 9628 60558
rect 9692 60556 9698 60620
rect 10174 60618 10180 60620
rect 10134 60558 10180 60618
rect 10244 60616 10291 60620
rect 10286 60560 10291 60616
rect 10174 60556 10180 60558
rect 10244 60556 10291 60560
rect 10225 60555 10291 60556
rect 0 60422 1410 60482
rect 0 60392 800 60422
rect 2576 60416 2896 60417
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2576 60351 2896 60352
rect 5839 60416 6159 60417
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 60351 6159 60352
rect 9103 60416 9423 60417
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 60351 9423 60352
rect 8661 60210 8727 60213
rect 11200 60210 12000 60240
rect 8661 60208 12000 60210
rect 8661 60152 8666 60208
rect 8722 60152 12000 60208
rect 8661 60150 12000 60152
rect 8661 60147 8727 60150
rect 11200 60120 12000 60150
rect 4207 59872 4527 59873
rect 0 59802 800 59832
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 59807 4527 59808
rect 7471 59872 7791 59873
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 59807 7791 59808
rect 1853 59802 1919 59805
rect 0 59800 1919 59802
rect 0 59744 1858 59800
rect 1914 59744 1919 59800
rect 0 59742 1919 59744
rect 0 59712 800 59742
rect 1853 59739 1919 59742
rect 9213 59802 9279 59805
rect 11200 59802 12000 59832
rect 9213 59800 12000 59802
rect 9213 59744 9218 59800
rect 9274 59744 12000 59800
rect 9213 59742 12000 59744
rect 9213 59739 9279 59742
rect 11200 59712 12000 59742
rect 1577 59530 1643 59533
rect 3366 59530 3372 59532
rect 1577 59528 3372 59530
rect 1577 59472 1582 59528
rect 1638 59472 3372 59528
rect 1577 59470 3372 59472
rect 1577 59467 1643 59470
rect 3366 59468 3372 59470
rect 3436 59468 3442 59532
rect 2576 59328 2896 59329
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 59263 2896 59264
rect 5839 59328 6159 59329
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 59263 6159 59264
rect 9103 59328 9423 59329
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 59263 9423 59264
rect 10041 59258 10107 59261
rect 11200 59258 12000 59288
rect 10041 59256 12000 59258
rect 10041 59200 10046 59256
rect 10102 59200 12000 59256
rect 10041 59198 12000 59200
rect 10041 59195 10107 59198
rect 11200 59168 12000 59198
rect 0 59122 800 59152
rect 1853 59122 1919 59125
rect 0 59120 1919 59122
rect 0 59064 1858 59120
rect 1914 59064 1919 59120
rect 0 59062 1919 59064
rect 0 59032 800 59062
rect 1853 59059 1919 59062
rect 9949 58850 10015 58853
rect 11200 58850 12000 58880
rect 9949 58848 12000 58850
rect 9949 58792 9954 58848
rect 10010 58792 12000 58848
rect 9949 58790 12000 58792
rect 9949 58787 10015 58790
rect 4207 58784 4527 58785
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 58719 4527 58720
rect 7471 58784 7791 58785
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 11200 58760 12000 58790
rect 7471 58719 7791 58720
rect 0 58442 800 58472
rect 1577 58442 1643 58445
rect 0 58440 1643 58442
rect 0 58384 1582 58440
rect 1638 58384 1643 58440
rect 0 58382 1643 58384
rect 0 58352 800 58382
rect 1577 58379 1643 58382
rect 10225 58306 10291 58309
rect 11200 58306 12000 58336
rect 10225 58304 12000 58306
rect 10225 58248 10230 58304
rect 10286 58248 12000 58304
rect 10225 58246 12000 58248
rect 10225 58243 10291 58246
rect 2576 58240 2896 58241
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 58175 2896 58176
rect 5839 58240 6159 58241
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 58175 6159 58176
rect 9103 58240 9423 58241
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 11200 58216 12000 58246
rect 9103 58175 9423 58176
rect 9949 57898 10015 57901
rect 11200 57898 12000 57928
rect 9949 57896 12000 57898
rect 9949 57840 9954 57896
rect 10010 57840 12000 57896
rect 9949 57838 12000 57840
rect 9949 57835 10015 57838
rect 11200 57808 12000 57838
rect 0 57762 800 57792
rect 1577 57762 1643 57765
rect 0 57760 1643 57762
rect 0 57704 1582 57760
rect 1638 57704 1643 57760
rect 0 57702 1643 57704
rect 0 57672 800 57702
rect 1577 57699 1643 57702
rect 4207 57696 4527 57697
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 4207 57631 4527 57632
rect 7471 57696 7791 57697
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 57631 7791 57632
rect 9213 57354 9279 57357
rect 11200 57354 12000 57384
rect 9213 57352 12000 57354
rect 9213 57296 9218 57352
rect 9274 57296 12000 57352
rect 9213 57294 12000 57296
rect 9213 57291 9279 57294
rect 11200 57264 12000 57294
rect 2576 57152 2896 57153
rect 0 57082 800 57112
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 57087 2896 57088
rect 5839 57152 6159 57153
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 57087 6159 57088
rect 9103 57152 9423 57153
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 57087 9423 57088
rect 1577 57082 1643 57085
rect 0 57080 1643 57082
rect 0 57024 1582 57080
rect 1638 57024 1643 57080
rect 0 57022 1643 57024
rect 0 56992 800 57022
rect 1577 57019 1643 57022
rect 10317 56946 10383 56949
rect 11200 56946 12000 56976
rect 10317 56944 12000 56946
rect 10317 56888 10322 56944
rect 10378 56888 12000 56944
rect 10317 56886 12000 56888
rect 10317 56883 10383 56886
rect 11200 56856 12000 56886
rect 4207 56608 4527 56609
rect 0 56538 800 56568
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 56543 4527 56544
rect 7471 56608 7791 56609
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 56543 7791 56544
rect 1577 56538 1643 56541
rect 0 56536 1643 56538
rect 0 56480 1582 56536
rect 1638 56480 1643 56536
rect 0 56478 1643 56480
rect 0 56448 800 56478
rect 1577 56475 1643 56478
rect 9581 56538 9647 56541
rect 11200 56538 12000 56568
rect 9581 56536 12000 56538
rect 9581 56480 9586 56536
rect 9642 56480 12000 56536
rect 9581 56478 12000 56480
rect 9581 56475 9647 56478
rect 11200 56448 12000 56478
rect 10726 56204 10732 56268
rect 10796 56266 10802 56268
rect 11697 56266 11763 56269
rect 10796 56264 11763 56266
rect 10796 56208 11702 56264
rect 11758 56208 11763 56264
rect 10796 56206 11763 56208
rect 10796 56204 10802 56206
rect 11697 56203 11763 56206
rect 2576 56064 2896 56065
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 55999 2896 56000
rect 5839 56064 6159 56065
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 55999 6159 56000
rect 9103 56064 9423 56065
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 55999 9423 56000
rect 9857 55994 9923 55997
rect 11200 55994 12000 56024
rect 9857 55992 12000 55994
rect 9857 55936 9862 55992
rect 9918 55936 12000 55992
rect 9857 55934 12000 55936
rect 9857 55931 9923 55934
rect 11200 55904 12000 55934
rect 0 55858 800 55888
rect 1577 55858 1643 55861
rect 0 55856 1643 55858
rect 0 55800 1582 55856
rect 1638 55800 1643 55856
rect 0 55798 1643 55800
rect 0 55768 800 55798
rect 1577 55795 1643 55798
rect 7966 55796 7972 55860
rect 8036 55858 8042 55860
rect 8569 55858 8635 55861
rect 8036 55856 8635 55858
rect 8036 55800 8574 55856
rect 8630 55800 8635 55856
rect 8036 55798 8635 55800
rect 8036 55796 8042 55798
rect 8569 55795 8635 55798
rect 9857 55586 9923 55589
rect 11200 55586 12000 55616
rect 9857 55584 12000 55586
rect 9857 55528 9862 55584
rect 9918 55528 12000 55584
rect 9857 55526 12000 55528
rect 9857 55523 9923 55526
rect 4207 55520 4527 55521
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 55455 4527 55456
rect 7471 55520 7791 55521
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 11200 55496 12000 55526
rect 7471 55455 7791 55456
rect 0 55178 800 55208
rect 1577 55178 1643 55181
rect 0 55176 1643 55178
rect 0 55120 1582 55176
rect 1638 55120 1643 55176
rect 0 55118 1643 55120
rect 0 55088 800 55118
rect 1577 55115 1643 55118
rect 9857 55042 9923 55045
rect 11200 55042 12000 55072
rect 9857 55040 12000 55042
rect 9857 54984 9862 55040
rect 9918 54984 12000 55040
rect 9857 54982 12000 54984
rect 9857 54979 9923 54982
rect 2576 54976 2896 54977
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 54911 2896 54912
rect 5839 54976 6159 54977
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 54911 6159 54912
rect 9103 54976 9423 54977
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 11200 54952 12000 54982
rect 9103 54911 9423 54912
rect 9949 54634 10015 54637
rect 11200 54634 12000 54664
rect 9949 54632 12000 54634
rect 9949 54576 9954 54632
rect 10010 54576 12000 54632
rect 9949 54574 12000 54576
rect 9949 54571 10015 54574
rect 11200 54544 12000 54574
rect 0 54498 800 54528
rect 1577 54498 1643 54501
rect 0 54496 1643 54498
rect 0 54440 1582 54496
rect 1638 54440 1643 54496
rect 0 54438 1643 54440
rect 0 54408 800 54438
rect 1577 54435 1643 54438
rect 4207 54432 4527 54433
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 54367 4527 54368
rect 7471 54432 7791 54433
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 54367 7791 54368
rect 11462 54300 11468 54364
rect 11532 54362 11538 54364
rect 11789 54362 11855 54365
rect 11532 54360 11855 54362
rect 11532 54304 11794 54360
rect 11850 54304 11855 54360
rect 11532 54302 11855 54304
rect 11532 54300 11538 54302
rect 11789 54299 11855 54302
rect 9581 54090 9647 54093
rect 11200 54090 12000 54120
rect 9581 54088 12000 54090
rect 9581 54032 9586 54088
rect 9642 54032 12000 54088
rect 9581 54030 12000 54032
rect 9581 54027 9647 54030
rect 11200 54000 12000 54030
rect 2576 53888 2896 53889
rect 0 53818 800 53848
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 53823 2896 53824
rect 5839 53888 6159 53889
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 53823 6159 53824
rect 9103 53888 9423 53889
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 53823 9423 53824
rect 1577 53818 1643 53821
rect 0 53816 1643 53818
rect 0 53760 1582 53816
rect 1638 53760 1643 53816
rect 0 53758 1643 53760
rect 0 53728 800 53758
rect 1577 53755 1643 53758
rect 9489 53682 9555 53685
rect 11200 53682 12000 53712
rect 9489 53680 12000 53682
rect 9489 53624 9494 53680
rect 9550 53624 12000 53680
rect 9489 53622 12000 53624
rect 9489 53619 9555 53622
rect 11200 53592 12000 53622
rect 8150 53484 8156 53548
rect 8220 53546 8226 53548
rect 8569 53546 8635 53549
rect 8220 53544 8635 53546
rect 8220 53488 8574 53544
rect 8630 53488 8635 53544
rect 8220 53486 8635 53488
rect 8220 53484 8226 53486
rect 8569 53483 8635 53486
rect 4207 53344 4527 53345
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 53279 4527 53280
rect 7471 53344 7791 53345
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 53279 7791 53280
rect 10358 53212 10364 53276
rect 10428 53274 10434 53276
rect 10961 53274 11027 53277
rect 10428 53272 11027 53274
rect 10428 53216 10966 53272
rect 11022 53216 11027 53272
rect 10428 53214 11027 53216
rect 10428 53212 10434 53214
rect 10961 53211 11027 53214
rect 0 53138 800 53168
rect 1577 53138 1643 53141
rect 0 53136 1643 53138
rect 0 53080 1582 53136
rect 1638 53080 1643 53136
rect 0 53078 1643 53080
rect 0 53048 800 53078
rect 1577 53075 1643 53078
rect 9949 53138 10015 53141
rect 11200 53138 12000 53168
rect 9949 53136 12000 53138
rect 9949 53080 9954 53136
rect 10010 53080 12000 53136
rect 9949 53078 12000 53080
rect 9949 53075 10015 53078
rect 11200 53048 12000 53078
rect 2576 52800 2896 52801
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 52735 2896 52736
rect 5839 52800 6159 52801
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 52735 6159 52736
rect 9103 52800 9423 52801
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 52735 9423 52736
rect 9857 52730 9923 52733
rect 11200 52730 12000 52760
rect 9857 52728 12000 52730
rect 9857 52672 9862 52728
rect 9918 52672 12000 52728
rect 9857 52670 12000 52672
rect 9857 52667 9923 52670
rect 11200 52640 12000 52670
rect 0 52458 800 52488
rect 2773 52458 2839 52461
rect 0 52456 2839 52458
rect 0 52400 2778 52456
rect 2834 52400 2839 52456
rect 0 52398 2839 52400
rect 0 52368 800 52398
rect 2773 52395 2839 52398
rect 10685 52458 10751 52461
rect 10910 52458 10916 52460
rect 10685 52456 10916 52458
rect 10685 52400 10690 52456
rect 10746 52400 10916 52456
rect 10685 52398 10916 52400
rect 10685 52395 10751 52398
rect 10910 52396 10916 52398
rect 10980 52396 10986 52460
rect 4207 52256 4527 52257
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 52191 4527 52192
rect 7471 52256 7791 52257
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 52191 7791 52192
rect 9121 52186 9187 52189
rect 11200 52186 12000 52216
rect 9121 52184 12000 52186
rect 9121 52128 9126 52184
rect 9182 52128 12000 52184
rect 9121 52126 12000 52128
rect 9121 52123 9187 52126
rect 11200 52096 12000 52126
rect 0 51914 800 51944
rect 1853 51914 1919 51917
rect 0 51912 1919 51914
rect 0 51856 1858 51912
rect 1914 51856 1919 51912
rect 0 51854 1919 51856
rect 0 51824 800 51854
rect 1853 51851 1919 51854
rect 9489 51778 9555 51781
rect 11200 51778 12000 51808
rect 9489 51776 12000 51778
rect 9489 51720 9494 51776
rect 9550 51720 12000 51776
rect 9489 51718 12000 51720
rect 9489 51715 9555 51718
rect 2576 51712 2896 51713
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 51647 2896 51648
rect 5839 51712 6159 51713
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 51647 6159 51648
rect 9103 51712 9423 51713
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 11200 51688 12000 51718
rect 9103 51647 9423 51648
rect 7046 51444 7052 51508
rect 7116 51506 7122 51508
rect 7189 51506 7255 51509
rect 10961 51506 11027 51509
rect 7116 51504 7255 51506
rect 7116 51448 7194 51504
rect 7250 51448 7255 51504
rect 7116 51446 7255 51448
rect 7116 51444 7122 51446
rect 7189 51443 7255 51446
rect 10780 51504 11027 51506
rect 10780 51448 10966 51504
rect 11022 51448 11027 51504
rect 10780 51446 11027 51448
rect 8293 51370 8359 51373
rect 7238 51368 8359 51370
rect 7238 51312 8298 51368
rect 8354 51312 8359 51368
rect 7238 51310 8359 51312
rect 0 51234 800 51264
rect 1393 51234 1459 51237
rect 0 51232 1459 51234
rect 0 51176 1398 51232
rect 1454 51176 1459 51232
rect 0 51174 1459 51176
rect 0 51144 800 51174
rect 1393 51171 1459 51174
rect 3049 51234 3115 51237
rect 3182 51234 3188 51236
rect 3049 51232 3188 51234
rect 3049 51176 3054 51232
rect 3110 51176 3188 51232
rect 3049 51174 3188 51176
rect 3049 51171 3115 51174
rect 3182 51172 3188 51174
rect 3252 51172 3258 51236
rect 6678 51172 6684 51236
rect 6748 51234 6754 51236
rect 7005 51234 7071 51237
rect 6748 51232 7071 51234
rect 6748 51176 7010 51232
rect 7066 51176 7071 51232
rect 6748 51174 7071 51176
rect 6748 51172 6754 51174
rect 7005 51171 7071 51174
rect 4207 51168 4527 51169
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 51103 4527 51104
rect 7005 51098 7071 51101
rect 7238 51098 7298 51310
rect 8293 51307 8359 51310
rect 8150 51172 8156 51236
rect 8220 51234 8226 51236
rect 8293 51234 8359 51237
rect 8220 51232 8359 51234
rect 8220 51176 8298 51232
rect 8354 51176 8359 51232
rect 8220 51174 8359 51176
rect 8220 51172 8226 51174
rect 8293 51171 8359 51174
rect 7471 51168 7791 51169
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 51103 7791 51104
rect 10780 51101 10840 51446
rect 10961 51443 11027 51446
rect 10961 51368 11027 51373
rect 10961 51312 10966 51368
rect 11022 51312 11027 51368
rect 10961 51307 11027 51312
rect 10964 51200 11024 51307
rect 11200 51234 12000 51264
rect 11148 51200 12000 51234
rect 10964 51144 12000 51200
rect 10964 51140 11208 51144
rect 8937 51098 9003 51101
rect 7005 51096 7298 51098
rect 7005 51040 7010 51096
rect 7066 51040 7298 51096
rect 7005 51038 7298 51040
rect 8894 51096 9003 51098
rect 8894 51040 8942 51096
rect 8998 51040 9003 51096
rect 7005 51035 7071 51038
rect 8894 51035 9003 51040
rect 10777 51096 10843 51101
rect 10777 51040 10782 51096
rect 10838 51040 10843 51096
rect 10777 51035 10843 51040
rect 3141 50964 3207 50965
rect 3141 50962 3188 50964
rect 3096 50960 3188 50962
rect 3096 50904 3146 50960
rect 3096 50902 3188 50904
rect 3141 50900 3188 50902
rect 3252 50900 3258 50964
rect 3601 50962 3667 50965
rect 3734 50962 3740 50964
rect 3601 50960 3740 50962
rect 3601 50904 3606 50960
rect 3662 50904 3740 50960
rect 3601 50902 3740 50904
rect 3141 50899 3207 50900
rect 3601 50899 3667 50902
rect 3734 50900 3740 50902
rect 3804 50900 3810 50964
rect 6678 50900 6684 50964
rect 6748 50962 6754 50964
rect 7005 50962 7071 50965
rect 6748 50960 7071 50962
rect 6748 50904 7010 50960
rect 7066 50904 7071 50960
rect 6748 50902 7071 50904
rect 6748 50900 6754 50902
rect 7005 50899 7071 50902
rect 2576 50624 2896 50625
rect 0 50554 800 50584
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 50559 2896 50560
rect 5839 50624 6159 50625
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 50559 6159 50560
rect 1853 50554 1919 50557
rect 0 50552 1919 50554
rect 0 50496 1858 50552
rect 1914 50496 1919 50552
rect 0 50494 1919 50496
rect 0 50464 800 50494
rect 1853 50491 1919 50494
rect 8150 50356 8156 50420
rect 8220 50418 8226 50420
rect 8385 50418 8451 50421
rect 8220 50416 8451 50418
rect 8220 50360 8390 50416
rect 8446 50360 8451 50416
rect 8220 50358 8451 50360
rect 8894 50418 8954 51035
rect 9857 50826 9923 50829
rect 11200 50826 12000 50856
rect 9857 50824 12000 50826
rect 9857 50768 9862 50824
rect 9918 50768 12000 50824
rect 9857 50766 12000 50768
rect 9857 50763 9923 50766
rect 11200 50736 12000 50766
rect 9103 50624 9423 50625
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 50559 9423 50560
rect 11329 50554 11395 50557
rect 11462 50554 11468 50556
rect 11329 50552 11468 50554
rect 11329 50496 11334 50552
rect 11390 50496 11468 50552
rect 11329 50494 11468 50496
rect 11329 50491 11395 50494
rect 11462 50492 11468 50494
rect 11532 50492 11538 50556
rect 9121 50418 9187 50421
rect 8894 50416 9187 50418
rect 8894 50360 9126 50416
rect 9182 50360 9187 50416
rect 8894 50358 9187 50360
rect 8220 50356 8226 50358
rect 8385 50355 8451 50358
rect 9121 50355 9187 50358
rect 8109 50282 8175 50285
rect 11200 50282 12000 50312
rect 8109 50280 12000 50282
rect 8109 50224 8114 50280
rect 8170 50224 12000 50280
rect 8109 50222 12000 50224
rect 8109 50219 8175 50222
rect 11200 50192 12000 50222
rect 9949 50146 10015 50149
rect 10726 50146 10732 50148
rect 9949 50144 10732 50146
rect 9949 50088 9954 50144
rect 10010 50088 10732 50144
rect 9949 50086 10732 50088
rect 9949 50083 10015 50086
rect 10726 50084 10732 50086
rect 10796 50084 10802 50148
rect 4207 50080 4527 50081
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 50015 4527 50016
rect 7471 50080 7791 50081
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7471 50015 7791 50016
rect 0 49874 800 49904
rect 1853 49874 1919 49877
rect 0 49872 1919 49874
rect 0 49816 1858 49872
rect 1914 49816 1919 49872
rect 0 49814 1919 49816
rect 0 49784 800 49814
rect 1853 49811 1919 49814
rect 8661 49874 8727 49877
rect 11200 49874 12000 49904
rect 8661 49872 12000 49874
rect 8661 49816 8666 49872
rect 8722 49816 12000 49872
rect 8661 49814 12000 49816
rect 8661 49811 8727 49814
rect 11200 49784 12000 49814
rect 3693 49738 3759 49741
rect 3693 49736 3986 49738
rect 3693 49680 3698 49736
rect 3754 49680 3986 49736
rect 3693 49678 3986 49680
rect 3693 49675 3759 49678
rect 3601 49602 3667 49605
rect 3785 49602 3851 49605
rect 3601 49600 3851 49602
rect 3601 49544 3606 49600
rect 3662 49544 3790 49600
rect 3846 49544 3851 49600
rect 3601 49542 3851 49544
rect 3601 49539 3667 49542
rect 3785 49539 3851 49542
rect 2576 49536 2896 49537
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 49471 2896 49472
rect 3693 49466 3759 49469
rect 3926 49466 3986 49678
rect 7005 49604 7071 49605
rect 7005 49602 7052 49604
rect 6960 49600 7052 49602
rect 6960 49544 7010 49600
rect 6960 49542 7052 49544
rect 7005 49540 7052 49542
rect 7116 49540 7122 49604
rect 7005 49539 7071 49540
rect 5839 49536 6159 49537
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5839 49471 6159 49472
rect 9103 49536 9423 49537
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 49471 9423 49472
rect 3693 49464 3986 49466
rect 3693 49408 3698 49464
rect 3754 49408 3986 49464
rect 3693 49406 3986 49408
rect 3693 49403 3759 49406
rect 10961 49330 11027 49333
rect 11200 49330 12000 49360
rect 10961 49328 12000 49330
rect 10961 49272 10966 49328
rect 11022 49272 12000 49328
rect 10961 49270 12000 49272
rect 10961 49267 11027 49270
rect 11200 49240 12000 49270
rect 0 49194 800 49224
rect 1853 49194 1919 49197
rect 0 49192 1919 49194
rect 0 49136 1858 49192
rect 1914 49136 1919 49192
rect 0 49134 1919 49136
rect 0 49104 800 49134
rect 1853 49131 1919 49134
rect 4207 48992 4527 48993
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 48927 4527 48928
rect 7471 48992 7791 48993
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7471 48927 7791 48928
rect 8201 48922 8267 48925
rect 11200 48922 12000 48952
rect 8201 48920 12000 48922
rect 8201 48864 8206 48920
rect 8262 48864 12000 48920
rect 8201 48862 12000 48864
rect 8201 48859 8267 48862
rect 11200 48832 12000 48862
rect 7741 48786 7807 48789
rect 8150 48786 8156 48788
rect 7741 48784 8156 48786
rect 7741 48728 7746 48784
rect 7802 48728 8156 48784
rect 7741 48726 8156 48728
rect 7741 48723 7807 48726
rect 8150 48724 8156 48726
rect 8220 48724 8226 48788
rect 8201 48650 8267 48653
rect 8201 48648 9874 48650
rect 8201 48592 8206 48648
rect 8262 48592 9874 48648
rect 8201 48590 9874 48592
rect 8201 48587 8267 48590
rect 0 48514 800 48544
rect 1853 48514 1919 48517
rect 0 48512 1919 48514
rect 0 48456 1858 48512
rect 1914 48456 1919 48512
rect 0 48454 1919 48456
rect 0 48424 800 48454
rect 1853 48451 1919 48454
rect 7966 48452 7972 48516
rect 8036 48514 8042 48516
rect 8845 48514 8911 48517
rect 8036 48512 8911 48514
rect 8036 48456 8850 48512
rect 8906 48456 8911 48512
rect 8036 48454 8911 48456
rect 8036 48452 8042 48454
rect 8845 48451 8911 48454
rect 2576 48448 2896 48449
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 48383 2896 48384
rect 5839 48448 6159 48449
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5839 48383 6159 48384
rect 9103 48448 9423 48449
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 48383 9423 48384
rect 9814 48378 9874 48590
rect 11200 48378 12000 48408
rect 9814 48318 12000 48378
rect 11200 48288 12000 48318
rect 7230 48044 7236 48108
rect 7300 48106 7306 48108
rect 7741 48106 7807 48109
rect 7300 48104 7807 48106
rect 7300 48048 7746 48104
rect 7802 48048 7807 48104
rect 7300 48046 7807 48048
rect 7300 48044 7306 48046
rect 7741 48043 7807 48046
rect 8201 47970 8267 47973
rect 11200 47970 12000 48000
rect 8201 47968 12000 47970
rect 8201 47912 8206 47968
rect 8262 47912 12000 47968
rect 8201 47910 12000 47912
rect 8201 47907 8267 47910
rect 4207 47904 4527 47905
rect 0 47834 800 47864
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 47839 4527 47840
rect 7471 47904 7791 47905
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 11200 47880 12000 47910
rect 7471 47839 7791 47840
rect 1853 47834 1919 47837
rect 0 47832 1919 47834
rect 0 47776 1858 47832
rect 1914 47776 1919 47832
rect 0 47774 1919 47776
rect 0 47744 800 47774
rect 1853 47771 1919 47774
rect 8150 47636 8156 47700
rect 8220 47698 8226 47700
rect 9213 47698 9279 47701
rect 8220 47696 9279 47698
rect 8220 47640 9218 47696
rect 9274 47640 9279 47696
rect 8220 47638 9279 47640
rect 8220 47636 8226 47638
rect 9213 47635 9279 47638
rect 2497 47562 2563 47565
rect 9121 47562 9187 47565
rect 2497 47560 9187 47562
rect 2497 47504 2502 47560
rect 2558 47504 9126 47560
rect 9182 47504 9187 47560
rect 2497 47502 9187 47504
rect 2497 47499 2563 47502
rect 9121 47499 9187 47502
rect 9489 47426 9555 47429
rect 11200 47426 12000 47456
rect 9489 47424 12000 47426
rect 9489 47368 9494 47424
rect 9550 47368 12000 47424
rect 9489 47366 12000 47368
rect 9489 47363 9555 47366
rect 2576 47360 2896 47361
rect 0 47290 800 47320
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 47295 2896 47296
rect 5839 47360 6159 47361
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 47295 6159 47296
rect 9103 47360 9423 47361
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 11200 47336 12000 47366
rect 9103 47295 9423 47296
rect 1853 47290 1919 47293
rect 0 47288 1919 47290
rect 0 47232 1858 47288
rect 1914 47232 1919 47288
rect 0 47230 1919 47232
rect 0 47200 800 47230
rect 1853 47227 1919 47230
rect 8201 47018 8267 47021
rect 11200 47018 12000 47048
rect 8201 47016 12000 47018
rect 8201 46960 8206 47016
rect 8262 46960 12000 47016
rect 8201 46958 12000 46960
rect 8201 46955 8267 46958
rect 11200 46928 12000 46958
rect 4207 46816 4527 46817
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 46751 4527 46752
rect 7471 46816 7791 46817
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 46751 7791 46752
rect 0 46610 800 46640
rect 1853 46610 1919 46613
rect 0 46608 1919 46610
rect 0 46552 1858 46608
rect 1914 46552 1919 46608
rect 0 46550 1919 46552
rect 0 46520 800 46550
rect 1853 46547 1919 46550
rect 9581 46610 9647 46613
rect 9581 46608 9690 46610
rect 9581 46552 9586 46608
rect 9642 46552 9690 46608
rect 9581 46547 9690 46552
rect 9489 46472 9555 46477
rect 9489 46416 9494 46472
rect 9550 46416 9555 46472
rect 9489 46411 9555 46416
rect 9630 46474 9690 46547
rect 11200 46474 12000 46504
rect 9630 46414 12000 46474
rect 7189 46338 7255 46341
rect 8017 46338 8083 46341
rect 7189 46336 8083 46338
rect 7189 46280 7194 46336
rect 7250 46280 8022 46336
rect 8078 46280 8083 46336
rect 7189 46278 8083 46280
rect 7189 46275 7255 46278
rect 8017 46275 8083 46278
rect 2576 46272 2896 46273
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 46207 2896 46208
rect 5839 46272 6159 46273
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 46207 6159 46208
rect 9103 46272 9423 46273
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 46207 9423 46208
rect 9492 46205 9552 46411
rect 11200 46384 12000 46414
rect 9949 46340 10015 46341
rect 9949 46338 9996 46340
rect 9904 46336 9996 46338
rect 9904 46280 9954 46336
rect 9904 46278 9996 46280
rect 9949 46276 9996 46278
rect 10060 46276 10066 46340
rect 10225 46338 10291 46341
rect 10225 46336 10426 46338
rect 10225 46280 10230 46336
rect 10286 46280 10426 46336
rect 10225 46278 10426 46280
rect 9949 46275 10015 46276
rect 10225 46275 10291 46278
rect 9489 46200 9555 46205
rect 9489 46144 9494 46200
rect 9550 46144 9555 46200
rect 9489 46139 9555 46144
rect 10366 46066 10426 46278
rect 11200 46066 12000 46096
rect 10366 46006 12000 46066
rect 11200 45976 12000 46006
rect 0 45930 800 45960
rect 1853 45930 1919 45933
rect 0 45928 1919 45930
rect 0 45872 1858 45928
rect 1914 45872 1919 45928
rect 0 45870 1919 45872
rect 0 45840 800 45870
rect 1853 45867 1919 45870
rect 4207 45728 4527 45729
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 45663 4527 45664
rect 7471 45728 7791 45729
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 45663 7791 45664
rect 11200 45568 12000 45688
rect 3785 45388 3851 45389
rect 3734 45386 3740 45388
rect 3694 45326 3740 45386
rect 3804 45384 3851 45388
rect 3846 45328 3851 45384
rect 3734 45324 3740 45326
rect 3804 45324 3851 45328
rect 3785 45323 3851 45324
rect 0 45250 800 45280
rect 1393 45250 1459 45253
rect 0 45248 1459 45250
rect 0 45192 1398 45248
rect 1454 45192 1459 45248
rect 0 45190 1459 45192
rect 0 45160 800 45190
rect 1393 45187 1459 45190
rect 2576 45184 2896 45185
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 45119 2896 45120
rect 5839 45184 6159 45185
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 45119 6159 45120
rect 9103 45184 9423 45185
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 45119 9423 45120
rect 11200 45024 12000 45144
rect 7966 44780 7972 44844
rect 8036 44842 8042 44844
rect 9397 44842 9463 44845
rect 8036 44840 9463 44842
rect 8036 44784 9402 44840
rect 9458 44784 9463 44840
rect 8036 44782 9463 44784
rect 8036 44780 8042 44782
rect 9397 44779 9463 44782
rect 8201 44706 8267 44709
rect 11200 44706 12000 44736
rect 8201 44704 12000 44706
rect 8201 44648 8206 44704
rect 8262 44648 12000 44704
rect 8201 44646 12000 44648
rect 8201 44643 8267 44646
rect 4207 44640 4527 44641
rect 0 44570 800 44600
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 44575 4527 44576
rect 7471 44640 7791 44641
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 11200 44616 12000 44646
rect 7471 44575 7791 44576
rect 1853 44570 1919 44573
rect 0 44568 1919 44570
rect 0 44512 1858 44568
rect 1914 44512 1919 44568
rect 0 44510 1919 44512
rect 0 44480 800 44510
rect 1853 44507 1919 44510
rect 9397 44570 9463 44573
rect 9397 44568 10058 44570
rect 9397 44512 9402 44568
rect 9458 44512 10058 44568
rect 9397 44510 10058 44512
rect 9397 44507 9463 44510
rect 3550 44372 3556 44436
rect 3620 44434 3626 44436
rect 9857 44434 9923 44437
rect 3620 44432 9923 44434
rect 3620 44376 9862 44432
rect 9918 44376 9923 44432
rect 3620 44374 9923 44376
rect 9998 44434 10058 44510
rect 11094 44434 11100 44436
rect 9998 44374 11100 44434
rect 3620 44372 3626 44374
rect 9857 44371 9923 44374
rect 11094 44372 11100 44374
rect 11164 44372 11170 44436
rect 7230 44236 7236 44300
rect 7300 44298 7306 44300
rect 7557 44298 7623 44301
rect 7300 44296 7623 44298
rect 7300 44240 7562 44296
rect 7618 44240 7623 44296
rect 7300 44238 7623 44240
rect 7300 44236 7306 44238
rect 7557 44235 7623 44238
rect 9213 44298 9279 44301
rect 9213 44296 9690 44298
rect 9213 44240 9218 44296
rect 9274 44240 9690 44296
rect 9213 44238 9690 44240
rect 9213 44235 9279 44238
rect 9630 44162 9690 44238
rect 11200 44162 12000 44192
rect 9630 44102 12000 44162
rect 2576 44096 2896 44097
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 44031 2896 44032
rect 5839 44096 6159 44097
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 44031 6159 44032
rect 9103 44096 9423 44097
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 11200 44072 12000 44102
rect 9103 44031 9423 44032
rect 0 43890 800 43920
rect 1853 43890 1919 43893
rect 0 43888 1919 43890
rect 0 43832 1858 43888
rect 1914 43832 1919 43888
rect 0 43830 1919 43832
rect 0 43800 800 43830
rect 1853 43827 1919 43830
rect 7281 43890 7347 43893
rect 9581 43890 9647 43893
rect 7281 43888 9647 43890
rect 7281 43832 7286 43888
rect 7342 43832 9586 43888
rect 9642 43832 9647 43888
rect 7281 43830 9647 43832
rect 7281 43827 7347 43830
rect 9581 43827 9647 43830
rect 9121 43754 9187 43757
rect 11200 43754 12000 43784
rect 9121 43752 12000 43754
rect 9121 43696 9126 43752
rect 9182 43696 12000 43752
rect 9121 43694 12000 43696
rect 9121 43691 9187 43694
rect 11200 43664 12000 43694
rect 4207 43552 4527 43553
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 43487 4527 43488
rect 7471 43552 7791 43553
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 43487 7791 43488
rect 11421 43484 11487 43485
rect 11421 43482 11468 43484
rect 11376 43480 11468 43482
rect 11376 43424 11426 43480
rect 11376 43422 11468 43424
rect 11421 43420 11468 43422
rect 11532 43420 11538 43484
rect 11421 43419 11487 43420
rect 0 43210 800 43240
rect 1853 43210 1919 43213
rect 0 43208 1919 43210
rect 0 43152 1858 43208
rect 1914 43152 1919 43208
rect 0 43150 1919 43152
rect 0 43120 800 43150
rect 1853 43147 1919 43150
rect 9857 43210 9923 43213
rect 11200 43210 12000 43240
rect 9857 43208 12000 43210
rect 9857 43152 9862 43208
rect 9918 43152 12000 43208
rect 9857 43150 12000 43152
rect 9857 43147 9923 43150
rect 11200 43120 12000 43150
rect 6637 43074 6703 43077
rect 8150 43074 8156 43076
rect 6637 43072 8156 43074
rect 6637 43016 6642 43072
rect 6698 43016 8156 43072
rect 6637 43014 8156 43016
rect 6637 43011 6703 43014
rect 8150 43012 8156 43014
rect 8220 43012 8226 43076
rect 2576 43008 2896 43009
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 42943 2896 42944
rect 5839 43008 6159 43009
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 42943 6159 42944
rect 9103 43008 9423 43009
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 42943 9423 42944
rect 6821 42802 6887 42805
rect 8334 42802 8340 42804
rect 6821 42800 8340 42802
rect 6821 42744 6826 42800
rect 6882 42744 8340 42800
rect 6821 42742 8340 42744
rect 6821 42739 6887 42742
rect 8334 42740 8340 42742
rect 8404 42740 8410 42804
rect 8569 42802 8635 42805
rect 11200 42802 12000 42832
rect 8569 42800 12000 42802
rect 8569 42744 8574 42800
rect 8630 42744 12000 42800
rect 8569 42742 12000 42744
rect 8569 42739 8635 42742
rect 11200 42712 12000 42742
rect 0 42666 800 42696
rect 1393 42666 1459 42669
rect 0 42664 1459 42666
rect 0 42608 1398 42664
rect 1454 42608 1459 42664
rect 0 42606 1459 42608
rect 0 42576 800 42606
rect 1393 42603 1459 42606
rect 5073 42666 5139 42669
rect 6085 42666 6151 42669
rect 6913 42666 6979 42669
rect 5073 42664 6979 42666
rect 5073 42608 5078 42664
rect 5134 42608 6090 42664
rect 6146 42608 6918 42664
rect 6974 42608 6979 42664
rect 5073 42606 6979 42608
rect 5073 42603 5139 42606
rect 6085 42603 6151 42606
rect 6913 42603 6979 42606
rect 10133 42666 10199 42669
rect 10726 42666 10732 42668
rect 10133 42664 10732 42666
rect 10133 42608 10138 42664
rect 10194 42608 10732 42664
rect 10133 42606 10732 42608
rect 10133 42603 10199 42606
rect 10726 42604 10732 42606
rect 10796 42604 10802 42668
rect 10542 42468 10548 42532
rect 10612 42530 10618 42532
rect 11513 42530 11579 42533
rect 10612 42528 11579 42530
rect 10612 42472 11518 42528
rect 11574 42472 11579 42528
rect 10612 42470 11579 42472
rect 10612 42468 10618 42470
rect 11513 42467 11579 42470
rect 4207 42464 4527 42465
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 42399 4527 42400
rect 7471 42464 7791 42465
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 42399 7791 42400
rect 10133 42394 10199 42397
rect 10358 42394 10364 42396
rect 10133 42392 10364 42394
rect 10133 42336 10138 42392
rect 10194 42336 10364 42392
rect 10133 42334 10364 42336
rect 10133 42331 10199 42334
rect 10358 42332 10364 42334
rect 10428 42332 10434 42396
rect 9121 42258 9187 42261
rect 11200 42258 12000 42288
rect 9121 42256 12000 42258
rect 9121 42200 9126 42256
rect 9182 42200 12000 42256
rect 9121 42198 12000 42200
rect 9121 42195 9187 42198
rect 11200 42168 12000 42198
rect 10133 42122 10199 42125
rect 10910 42122 10916 42124
rect 10133 42120 10916 42122
rect 10133 42064 10138 42120
rect 10194 42064 10916 42120
rect 10133 42062 10916 42064
rect 10133 42059 10199 42062
rect 10910 42060 10916 42062
rect 10980 42060 10986 42124
rect 0 41986 800 42016
rect 1393 41986 1459 41989
rect 0 41984 1459 41986
rect 0 41928 1398 41984
rect 1454 41928 1459 41984
rect 0 41926 1459 41928
rect 0 41896 800 41926
rect 1393 41923 1459 41926
rect 2576 41920 2896 41921
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 41855 2896 41856
rect 5839 41920 6159 41921
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5839 41855 6159 41856
rect 9103 41920 9423 41921
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 41855 9423 41856
rect 9949 41850 10015 41853
rect 11200 41850 12000 41880
rect 9949 41848 12000 41850
rect 9949 41792 9954 41848
rect 10010 41792 12000 41848
rect 9949 41790 12000 41792
rect 9949 41787 10015 41790
rect 11200 41760 12000 41790
rect 10685 41714 10751 41717
rect 10685 41712 10794 41714
rect 10685 41656 10690 41712
rect 10746 41656 10794 41712
rect 10685 41651 10794 41656
rect 8150 41516 8156 41580
rect 8220 41578 8226 41580
rect 8753 41578 8819 41581
rect 8220 41576 8819 41578
rect 8220 41520 8758 41576
rect 8814 41520 8819 41576
rect 8220 41518 8819 41520
rect 8220 41516 8226 41518
rect 8753 41515 8819 41518
rect 10734 41445 10794 41651
rect 10734 41440 10843 41445
rect 10734 41384 10782 41440
rect 10838 41384 10843 41440
rect 10734 41382 10843 41384
rect 10777 41379 10843 41382
rect 4207 41376 4527 41377
rect 0 41306 800 41336
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 41311 4527 41312
rect 7471 41376 7791 41377
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 7471 41311 7791 41312
rect 1393 41306 1459 41309
rect 0 41304 1459 41306
rect 0 41248 1398 41304
rect 1454 41248 1459 41304
rect 0 41246 1459 41248
rect 0 41216 800 41246
rect 1393 41243 1459 41246
rect 8150 41244 8156 41308
rect 8220 41306 8226 41308
rect 8477 41306 8543 41309
rect 8220 41304 8543 41306
rect 8220 41248 8482 41304
rect 8538 41248 8543 41304
rect 8220 41246 8543 41248
rect 8220 41244 8226 41246
rect 8477 41243 8543 41246
rect 9949 41304 10015 41309
rect 11200 41306 12000 41336
rect 9949 41248 9954 41304
rect 10010 41248 10015 41304
rect 9949 41243 10015 41248
rect 10918 41246 12000 41306
rect 9952 41170 10012 41243
rect 10918 41170 10978 41246
rect 11200 41216 12000 41246
rect 9952 41110 10978 41170
rect 9949 40898 10015 40901
rect 11200 40898 12000 40928
rect 9949 40896 12000 40898
rect 9949 40840 9954 40896
rect 10010 40840 12000 40896
rect 9949 40838 12000 40840
rect 9949 40835 10015 40838
rect 2576 40832 2896 40833
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2576 40767 2896 40768
rect 5839 40832 6159 40833
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 40767 6159 40768
rect 9103 40832 9423 40833
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 11200 40808 12000 40838
rect 9103 40767 9423 40768
rect 8569 40764 8635 40765
rect 8518 40762 8524 40764
rect 8478 40702 8524 40762
rect 8588 40760 8635 40764
rect 8630 40704 8635 40760
rect 8518 40700 8524 40702
rect 8588 40700 8635 40704
rect 8569 40699 8635 40700
rect 0 40626 800 40656
rect 1853 40626 1919 40629
rect 0 40624 1919 40626
rect 0 40568 1858 40624
rect 1914 40568 1919 40624
rect 0 40566 1919 40568
rect 0 40536 800 40566
rect 1853 40563 1919 40566
rect 5073 40490 5139 40493
rect 10133 40492 10199 40493
rect 7966 40490 7972 40492
rect 5073 40488 7972 40490
rect 5073 40432 5078 40488
rect 5134 40432 7972 40488
rect 5073 40430 7972 40432
rect 5073 40427 5139 40430
rect 7966 40428 7972 40430
rect 8036 40428 8042 40492
rect 10133 40490 10180 40492
rect 10088 40488 10180 40490
rect 10088 40432 10138 40488
rect 10088 40430 10180 40432
rect 10133 40428 10180 40430
rect 10244 40428 10250 40492
rect 10133 40427 10199 40428
rect 8201 40354 8267 40357
rect 11200 40354 12000 40384
rect 8201 40352 12000 40354
rect 8201 40296 8206 40352
rect 8262 40296 12000 40352
rect 8201 40294 12000 40296
rect 8201 40291 8267 40294
rect 4207 40288 4527 40289
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 40223 4527 40224
rect 7471 40288 7791 40289
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 11200 40264 12000 40294
rect 7471 40223 7791 40224
rect 10542 40156 10548 40220
rect 10612 40218 10618 40220
rect 10777 40218 10843 40221
rect 10612 40216 10843 40218
rect 10612 40160 10782 40216
rect 10838 40160 10843 40216
rect 10612 40158 10843 40160
rect 10612 40156 10618 40158
rect 10777 40155 10843 40158
rect 0 39946 800 39976
rect 1393 39946 1459 39949
rect 0 39944 1459 39946
rect 0 39888 1398 39944
rect 1454 39888 1459 39944
rect 0 39886 1459 39888
rect 0 39856 800 39886
rect 1393 39883 1459 39886
rect 9305 39946 9371 39949
rect 11200 39946 12000 39976
rect 9305 39944 12000 39946
rect 9305 39888 9310 39944
rect 9366 39888 12000 39944
rect 9305 39886 12000 39888
rect 9305 39883 9371 39886
rect 11200 39856 12000 39886
rect 2576 39744 2896 39745
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 39679 2896 39680
rect 5839 39744 6159 39745
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 39679 6159 39680
rect 9103 39744 9423 39745
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 39679 9423 39680
rect 9857 39674 9923 39677
rect 10358 39674 10364 39676
rect 9857 39672 10364 39674
rect 9857 39616 9862 39672
rect 9918 39616 10364 39672
rect 9857 39614 10364 39616
rect 9857 39611 9923 39614
rect 10358 39612 10364 39614
rect 10428 39612 10434 39676
rect 10910 39612 10916 39676
rect 10980 39674 10986 39676
rect 11881 39674 11947 39677
rect 10980 39672 11947 39674
rect 10980 39616 11886 39672
rect 11942 39616 11947 39672
rect 10980 39614 11947 39616
rect 10980 39612 10986 39614
rect 11881 39611 11947 39614
rect 2221 39538 2287 39541
rect 8518 39538 8524 39540
rect 2221 39536 8524 39538
rect 2221 39480 2226 39536
rect 2282 39480 8524 39536
rect 2221 39478 8524 39480
rect 2221 39475 2287 39478
rect 8518 39476 8524 39478
rect 8588 39538 8594 39540
rect 9397 39538 9463 39541
rect 8588 39536 9463 39538
rect 8588 39480 9402 39536
rect 9458 39480 9463 39536
rect 8588 39478 9463 39480
rect 8588 39476 8594 39478
rect 9397 39475 9463 39478
rect 7465 39402 7531 39405
rect 6686 39400 7531 39402
rect 6686 39344 7470 39400
rect 7526 39344 7531 39400
rect 6686 39342 7531 39344
rect 0 39266 800 39296
rect 1853 39266 1919 39269
rect 0 39264 1919 39266
rect 0 39208 1858 39264
rect 1914 39208 1919 39264
rect 0 39206 1919 39208
rect 0 39176 800 39206
rect 1853 39203 1919 39206
rect 4207 39200 4527 39201
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 39135 4527 39136
rect 6545 39130 6611 39133
rect 6686 39130 6746 39342
rect 7465 39339 7531 39342
rect 8661 39402 8727 39405
rect 11200 39402 12000 39432
rect 8661 39400 12000 39402
rect 8661 39344 8666 39400
rect 8722 39344 12000 39400
rect 8661 39342 12000 39344
rect 8661 39339 8727 39342
rect 11200 39312 12000 39342
rect 7471 39200 7791 39201
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 39135 7791 39136
rect 6545 39128 6746 39130
rect 6545 39072 6550 39128
rect 6606 39072 6746 39128
rect 6545 39070 6746 39072
rect 6545 39067 6611 39070
rect 10041 38994 10107 38997
rect 11200 38994 12000 39024
rect 10041 38992 12000 38994
rect 10041 38936 10046 38992
rect 10102 38936 12000 38992
rect 10041 38934 12000 38936
rect 10041 38931 10107 38934
rect 11200 38904 12000 38934
rect 8886 38796 8892 38860
rect 8956 38858 8962 38860
rect 9121 38858 9187 38861
rect 8956 38856 9187 38858
rect 8956 38800 9126 38856
rect 9182 38800 9187 38856
rect 8956 38798 9187 38800
rect 8956 38796 8962 38798
rect 9121 38795 9187 38798
rect 11462 38660 11468 38724
rect 11532 38722 11538 38724
rect 11605 38722 11671 38725
rect 11532 38720 11671 38722
rect 11532 38664 11610 38720
rect 11666 38664 11671 38720
rect 11532 38662 11671 38664
rect 11532 38660 11538 38662
rect 11605 38659 11671 38662
rect 2576 38656 2896 38657
rect 0 38586 800 38616
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 38591 2896 38592
rect 5839 38656 6159 38657
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 38591 6159 38592
rect 9103 38656 9423 38657
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 9103 38591 9423 38592
rect 1393 38586 1459 38589
rect 0 38584 1459 38586
rect 0 38528 1398 38584
rect 1454 38528 1459 38584
rect 0 38526 1459 38528
rect 0 38496 800 38526
rect 1393 38523 1459 38526
rect 9765 38588 9831 38589
rect 9765 38584 9812 38588
rect 9876 38586 9882 38588
rect 9765 38528 9770 38584
rect 9765 38524 9812 38528
rect 9876 38526 9922 38586
rect 9876 38524 9882 38526
rect 9765 38523 9831 38524
rect 7005 38450 7071 38453
rect 8109 38450 8175 38453
rect 11200 38450 12000 38480
rect 7005 38448 7114 38450
rect 7005 38392 7010 38448
rect 7066 38392 7114 38448
rect 7005 38387 7114 38392
rect 8109 38448 9506 38450
rect 8109 38392 8114 38448
rect 8170 38416 9506 38448
rect 9630 38416 12000 38450
rect 8170 38392 12000 38416
rect 8109 38390 12000 38392
rect 8109 38387 8175 38390
rect 7054 38181 7114 38387
rect 9446 38356 9690 38390
rect 11200 38360 12000 38390
rect 7741 38314 7807 38317
rect 8334 38314 8340 38316
rect 7741 38312 8340 38314
rect 7741 38256 7746 38312
rect 7802 38256 8340 38312
rect 7741 38254 8340 38256
rect 7741 38251 7807 38254
rect 8334 38252 8340 38254
rect 8404 38252 8410 38316
rect 8518 38252 8524 38316
rect 8588 38314 8594 38316
rect 9121 38314 9187 38317
rect 8588 38312 9187 38314
rect 8588 38256 9126 38312
rect 9182 38256 9187 38312
rect 8588 38254 9187 38256
rect 8588 38252 8594 38254
rect 9121 38251 9187 38254
rect 7005 38176 7114 38181
rect 7005 38120 7010 38176
rect 7066 38120 7114 38176
rect 7005 38118 7114 38120
rect 7005 38115 7071 38118
rect 8886 38116 8892 38180
rect 8956 38178 8962 38180
rect 9213 38178 9279 38181
rect 8956 38176 9279 38178
rect 8956 38120 9218 38176
rect 9274 38120 9279 38176
rect 8956 38118 9279 38120
rect 8956 38116 8962 38118
rect 9213 38115 9279 38118
rect 4207 38112 4527 38113
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 38047 4527 38048
rect 7471 38112 7791 38113
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 38047 7791 38048
rect 8109 38042 8175 38045
rect 11200 38042 12000 38072
rect 8109 38040 12000 38042
rect 8109 37984 8114 38040
rect 8170 37984 12000 38040
rect 8109 37982 12000 37984
rect 8109 37979 8175 37982
rect 11200 37952 12000 37982
rect 0 37906 800 37936
rect 1393 37906 1459 37909
rect 0 37904 1459 37906
rect 0 37848 1398 37904
rect 1454 37848 1459 37904
rect 0 37846 1459 37848
rect 0 37816 800 37846
rect 1393 37843 1459 37846
rect 8518 37844 8524 37908
rect 8588 37906 8594 37908
rect 9305 37906 9371 37909
rect 8588 37904 9371 37906
rect 8588 37848 9310 37904
rect 9366 37848 9371 37904
rect 8588 37846 9371 37848
rect 8588 37844 8594 37846
rect 9305 37843 9371 37846
rect 2681 37770 2747 37773
rect 9622 37770 9628 37772
rect 2681 37768 9628 37770
rect 2681 37712 2686 37768
rect 2742 37712 9628 37768
rect 2681 37710 9628 37712
rect 2681 37707 2747 37710
rect 9622 37708 9628 37710
rect 9692 37708 9698 37772
rect 2576 37568 2896 37569
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 37503 2896 37504
rect 5839 37568 6159 37569
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 37503 6159 37504
rect 9103 37568 9423 37569
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 37503 9423 37504
rect 9581 37498 9647 37501
rect 11200 37498 12000 37528
rect 9581 37496 12000 37498
rect 9581 37440 9586 37496
rect 9642 37440 12000 37496
rect 9581 37438 12000 37440
rect 9581 37435 9647 37438
rect 11200 37408 12000 37438
rect 0 37362 800 37392
rect 1301 37362 1367 37365
rect 0 37360 1367 37362
rect 0 37304 1306 37360
rect 1362 37304 1367 37360
rect 0 37302 1367 37304
rect 0 37272 800 37302
rect 1301 37299 1367 37302
rect 3366 37164 3372 37228
rect 3436 37226 3442 37228
rect 8109 37226 8175 37229
rect 3436 37224 8175 37226
rect 3436 37168 8114 37224
rect 8170 37168 8175 37224
rect 3436 37166 8175 37168
rect 3436 37164 3442 37166
rect 8109 37163 8175 37166
rect 8109 37090 8175 37093
rect 11200 37090 12000 37120
rect 8109 37088 12000 37090
rect 8109 37032 8114 37088
rect 8170 37032 12000 37088
rect 8109 37030 12000 37032
rect 8109 37027 8175 37030
rect 4207 37024 4527 37025
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 36959 4527 36960
rect 7471 37024 7791 37025
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 11200 37000 12000 37030
rect 7471 36959 7791 36960
rect 10593 36820 10659 36821
rect 10542 36818 10548 36820
rect 10502 36758 10548 36818
rect 10612 36816 10659 36820
rect 11605 36820 11671 36821
rect 11605 36818 11652 36820
rect 10654 36760 10659 36816
rect 10542 36756 10548 36758
rect 10612 36756 10659 36760
rect 11560 36816 11652 36818
rect 11560 36760 11610 36816
rect 11560 36758 11652 36760
rect 10593 36755 10659 36756
rect 11605 36756 11652 36758
rect 11716 36756 11722 36820
rect 11605 36755 11671 36756
rect 0 36682 800 36712
rect 1393 36682 1459 36685
rect 0 36680 1459 36682
rect 0 36624 1398 36680
rect 1454 36624 1459 36680
rect 0 36622 1459 36624
rect 0 36592 800 36622
rect 1393 36619 1459 36622
rect 8109 36682 8175 36685
rect 8109 36680 9690 36682
rect 8109 36624 8114 36680
rect 8170 36624 9690 36680
rect 8109 36622 9690 36624
rect 8109 36619 8175 36622
rect 9630 36546 9690 36622
rect 10174 36620 10180 36684
rect 10244 36682 10250 36684
rect 10501 36682 10567 36685
rect 10244 36680 10567 36682
rect 10244 36624 10506 36680
rect 10562 36624 10567 36680
rect 10244 36622 10567 36624
rect 10244 36620 10250 36622
rect 10501 36619 10567 36622
rect 11200 36546 12000 36576
rect 9630 36486 12000 36546
rect 2576 36480 2896 36481
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 36415 2896 36416
rect 5839 36480 6159 36481
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 36415 6159 36416
rect 9103 36480 9423 36481
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 11200 36456 12000 36486
rect 9103 36415 9423 36416
rect 8334 36212 8340 36276
rect 8404 36274 8410 36276
rect 9397 36274 9463 36277
rect 8404 36272 9463 36274
rect 8404 36216 9402 36272
rect 9458 36216 9463 36272
rect 8404 36214 9463 36216
rect 8404 36212 8410 36214
rect 9397 36211 9463 36214
rect 8845 36138 8911 36141
rect 11200 36138 12000 36168
rect 8845 36136 12000 36138
rect 8845 36080 8850 36136
rect 8906 36080 12000 36136
rect 8845 36078 12000 36080
rect 8845 36075 8911 36078
rect 11200 36048 12000 36078
rect 0 36002 800 36032
rect 1577 36002 1643 36005
rect 0 36000 1643 36002
rect 0 35944 1582 36000
rect 1638 35944 1643 36000
rect 0 35942 1643 35944
rect 0 35912 800 35942
rect 1577 35939 1643 35942
rect 8845 36004 8911 36005
rect 8845 36000 8892 36004
rect 8956 36002 8962 36004
rect 8845 35944 8850 36000
rect 8845 35940 8892 35944
rect 8956 35942 9002 36002
rect 8956 35940 8962 35942
rect 8845 35939 8911 35940
rect 4207 35936 4527 35937
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 35871 4527 35872
rect 7471 35936 7791 35937
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 35871 7791 35872
rect 8845 35594 8911 35597
rect 11200 35594 12000 35624
rect 8845 35592 12000 35594
rect 8845 35536 8850 35592
rect 8906 35536 12000 35592
rect 8845 35534 12000 35536
rect 8845 35531 8911 35534
rect 11200 35504 12000 35534
rect 2576 35392 2896 35393
rect 0 35322 800 35352
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 35327 2896 35328
rect 5839 35392 6159 35393
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 35327 6159 35328
rect 9103 35392 9423 35393
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 35327 9423 35328
rect 1577 35322 1643 35325
rect 0 35320 1643 35322
rect 0 35264 1582 35320
rect 1638 35264 1643 35320
rect 0 35262 1643 35264
rect 0 35232 800 35262
rect 1577 35259 1643 35262
rect 8109 35186 8175 35189
rect 11200 35186 12000 35216
rect 8109 35184 12000 35186
rect 8109 35128 8114 35184
rect 8170 35128 12000 35184
rect 8109 35126 12000 35128
rect 8109 35123 8175 35126
rect 11200 35096 12000 35126
rect 4207 34848 4527 34849
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 34783 4527 34784
rect 7471 34848 7791 34849
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 34783 7791 34784
rect 0 34642 800 34672
rect 1577 34642 1643 34645
rect 0 34640 1643 34642
rect 0 34584 1582 34640
rect 1638 34584 1643 34640
rect 0 34582 1643 34584
rect 0 34552 800 34582
rect 1577 34579 1643 34582
rect 10133 34642 10199 34645
rect 11200 34642 12000 34672
rect 10133 34640 12000 34642
rect 10133 34584 10138 34640
rect 10194 34584 12000 34640
rect 10133 34582 12000 34584
rect 10133 34579 10199 34582
rect 11200 34552 12000 34582
rect 8661 34508 8727 34509
rect 8661 34504 8708 34508
rect 8772 34506 8778 34508
rect 8661 34448 8666 34504
rect 8661 34444 8708 34448
rect 8772 34446 8818 34506
rect 8772 34444 8778 34446
rect 8661 34443 8727 34444
rect 2576 34304 2896 34305
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 34239 2896 34240
rect 5839 34304 6159 34305
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 34239 6159 34240
rect 9103 34304 9423 34305
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 34239 9423 34240
rect 10041 34234 10107 34237
rect 11200 34234 12000 34264
rect 10041 34232 12000 34234
rect 10041 34176 10046 34232
rect 10102 34176 12000 34232
rect 10041 34174 12000 34176
rect 10041 34171 10107 34174
rect 11200 34144 12000 34174
rect 0 33962 800 33992
rect 1393 33962 1459 33965
rect 0 33960 1459 33962
rect 0 33904 1398 33960
rect 1454 33904 1459 33960
rect 0 33902 1459 33904
rect 0 33872 800 33902
rect 1393 33899 1459 33902
rect 9305 33826 9371 33829
rect 11200 33826 12000 33856
rect 9305 33824 12000 33826
rect 9305 33768 9310 33824
rect 9366 33768 12000 33824
rect 9305 33766 12000 33768
rect 9305 33763 9371 33766
rect 4207 33760 4527 33761
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 33695 4527 33696
rect 7471 33760 7791 33761
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 11200 33736 12000 33766
rect 7471 33695 7791 33696
rect 8518 33492 8524 33556
rect 8588 33554 8594 33556
rect 9581 33554 9647 33557
rect 8588 33552 9647 33554
rect 8588 33496 9586 33552
rect 9642 33496 9647 33552
rect 8588 33494 9647 33496
rect 8588 33492 8594 33494
rect 9581 33491 9647 33494
rect 8569 33418 8635 33421
rect 8526 33416 8635 33418
rect 8526 33360 8574 33416
rect 8630 33360 8635 33416
rect 8526 33355 8635 33360
rect 10409 33418 10475 33421
rect 10542 33418 10548 33420
rect 10409 33416 10548 33418
rect 10409 33360 10414 33416
rect 10470 33360 10548 33416
rect 10409 33358 10548 33360
rect 10409 33355 10475 33358
rect 10542 33356 10548 33358
rect 10612 33356 10618 33420
rect 0 33282 800 33312
rect 1393 33282 1459 33285
rect 0 33280 1459 33282
rect 0 33224 1398 33280
rect 1454 33224 1459 33280
rect 0 33222 1459 33224
rect 0 33192 800 33222
rect 1393 33219 1459 33222
rect 2576 33216 2896 33217
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 33151 2896 33152
rect 5839 33216 6159 33217
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 33151 6159 33152
rect 8526 33149 8586 33355
rect 9581 33282 9647 33285
rect 11200 33282 12000 33312
rect 9581 33280 12000 33282
rect 9581 33224 9586 33280
rect 9642 33224 12000 33280
rect 9581 33222 12000 33224
rect 9581 33219 9647 33222
rect 9103 33216 9423 33217
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 11200 33192 12000 33222
rect 9103 33151 9423 33152
rect 8526 33144 8635 33149
rect 10593 33148 10659 33149
rect 8526 33088 8574 33144
rect 8630 33088 8635 33144
rect 8526 33086 8635 33088
rect 8569 33083 8635 33086
rect 10542 33084 10548 33148
rect 10612 33146 10659 33148
rect 10612 33144 10704 33146
rect 10654 33088 10704 33144
rect 10612 33086 10704 33088
rect 10612 33084 10659 33086
rect 10593 33083 10659 33084
rect 10041 32874 10107 32877
rect 11200 32874 12000 32904
rect 10041 32872 12000 32874
rect 10041 32816 10046 32872
rect 10102 32816 12000 32872
rect 10041 32814 12000 32816
rect 10041 32811 10107 32814
rect 11200 32784 12000 32814
rect 0 32738 800 32768
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32648 800 32678
rect 1577 32675 1643 32678
rect 4207 32672 4527 32673
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 32607 4527 32608
rect 7471 32672 7791 32673
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 32607 7791 32608
rect 10726 32540 10732 32604
rect 10796 32602 10802 32604
rect 11881 32602 11947 32605
rect 10796 32600 11947 32602
rect 10796 32544 11886 32600
rect 11942 32544 11947 32600
rect 10796 32542 11947 32544
rect 10796 32540 10802 32542
rect 11881 32539 11947 32542
rect 9213 32330 9279 32333
rect 11200 32330 12000 32360
rect 9213 32328 12000 32330
rect 9213 32272 9218 32328
rect 9274 32272 12000 32328
rect 9213 32270 12000 32272
rect 9213 32267 9279 32270
rect 11200 32240 12000 32270
rect 2576 32128 2896 32129
rect 0 32058 800 32088
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 32063 2896 32064
rect 5839 32128 6159 32129
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 32063 6159 32064
rect 9103 32128 9423 32129
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 32063 9423 32064
rect 1577 32058 1643 32061
rect 0 32056 1643 32058
rect 0 32000 1582 32056
rect 1638 32000 1643 32056
rect 0 31998 1643 32000
rect 0 31968 800 31998
rect 1577 31995 1643 31998
rect 10501 32058 10567 32061
rect 10726 32058 10732 32060
rect 10501 32056 10732 32058
rect 10501 32000 10506 32056
rect 10562 32000 10732 32056
rect 10501 31998 10732 32000
rect 10501 31995 10567 31998
rect 10726 31996 10732 31998
rect 10796 31996 10802 32060
rect 8845 31922 8911 31925
rect 11200 31922 12000 31952
rect 8845 31920 12000 31922
rect 8845 31864 8850 31920
rect 8906 31864 12000 31920
rect 8845 31862 12000 31864
rect 8845 31859 8911 31862
rect 11200 31832 12000 31862
rect 10542 31724 10548 31788
rect 10612 31786 10618 31788
rect 10612 31726 11116 31786
rect 10612 31724 10618 31726
rect 10869 31650 10935 31653
rect 10869 31648 10978 31650
rect 10869 31592 10874 31648
rect 10930 31592 10978 31648
rect 10869 31587 10978 31592
rect 4207 31584 4527 31585
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 31519 4527 31520
rect 7471 31584 7791 31585
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 31519 7791 31520
rect 10918 31514 10978 31587
rect 10734 31454 10978 31514
rect 0 31378 800 31408
rect 1577 31378 1643 31381
rect 0 31376 1643 31378
rect 0 31320 1582 31376
rect 1638 31320 1643 31376
rect 0 31318 1643 31320
rect 0 31288 800 31318
rect 1577 31315 1643 31318
rect 10593 31242 10659 31245
rect 10734 31242 10794 31454
rect 11056 31378 11116 31726
rect 11200 31378 12000 31408
rect 11056 31318 12000 31378
rect 11200 31288 12000 31318
rect 10593 31240 10794 31242
rect 10593 31184 10598 31240
rect 10654 31184 10794 31240
rect 10593 31182 10794 31184
rect 10593 31179 10659 31182
rect 2576 31040 2896 31041
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 30975 2896 30976
rect 5839 31040 6159 31041
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 30975 6159 30976
rect 9103 31040 9423 31041
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 30975 9423 30976
rect 10409 30970 10475 30973
rect 11200 30970 12000 31000
rect 10409 30968 12000 30970
rect 10409 30912 10414 30968
rect 10470 30912 12000 30968
rect 10409 30910 12000 30912
rect 10409 30907 10475 30910
rect 11200 30880 12000 30910
rect 9990 30772 9996 30836
rect 10060 30834 10066 30836
rect 10409 30834 10475 30837
rect 10060 30832 10475 30834
rect 10060 30776 10414 30832
rect 10470 30776 10475 30832
rect 10060 30774 10475 30776
rect 10060 30772 10066 30774
rect 10409 30771 10475 30774
rect 0 30698 800 30728
rect 1577 30698 1643 30701
rect 0 30696 1643 30698
rect 0 30640 1582 30696
rect 1638 30640 1643 30696
rect 0 30638 1643 30640
rect 0 30608 800 30638
rect 1577 30635 1643 30638
rect 10133 30562 10199 30565
rect 10726 30562 10732 30564
rect 10133 30560 10732 30562
rect 10133 30504 10138 30560
rect 10194 30504 10732 30560
rect 10133 30502 10732 30504
rect 10133 30499 10199 30502
rect 10726 30500 10732 30502
rect 10796 30500 10802 30564
rect 4207 30496 4527 30497
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 30431 4527 30432
rect 7471 30496 7791 30497
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 30431 7791 30432
rect 10041 30426 10107 30429
rect 11200 30426 12000 30456
rect 10041 30424 12000 30426
rect 10041 30368 10046 30424
rect 10102 30368 12000 30424
rect 10041 30366 12000 30368
rect 10041 30363 10107 30366
rect 11200 30336 12000 30366
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 10041 30018 10107 30021
rect 11200 30018 12000 30048
rect 10041 30016 12000 30018
rect 10041 29960 10046 30016
rect 10102 29960 12000 30016
rect 10041 29958 12000 29960
rect 10041 29955 10107 29958
rect 2576 29952 2896 29953
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 29887 2896 29888
rect 5839 29952 6159 29953
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 29887 6159 29888
rect 9103 29952 9423 29953
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 11200 29928 12000 29958
rect 9103 29887 9423 29888
rect 9806 29684 9812 29748
rect 9876 29746 9882 29748
rect 10041 29746 10107 29749
rect 9876 29744 10107 29746
rect 9876 29688 10046 29744
rect 10102 29688 10107 29744
rect 9876 29686 10107 29688
rect 9876 29684 9882 29686
rect 10041 29683 10107 29686
rect 11646 29684 11652 29748
rect 11716 29746 11722 29748
rect 11881 29746 11947 29749
rect 11716 29744 11947 29746
rect 11716 29688 11886 29744
rect 11942 29688 11947 29744
rect 11716 29686 11947 29688
rect 11716 29684 11722 29686
rect 11881 29683 11947 29686
rect 10133 29612 10199 29613
rect 10133 29610 10180 29612
rect 10088 29608 10180 29610
rect 10088 29552 10138 29608
rect 10088 29550 10180 29552
rect 10133 29548 10180 29550
rect 10244 29548 10250 29612
rect 10133 29547 10199 29548
rect 9305 29474 9371 29477
rect 11200 29474 12000 29504
rect 9305 29472 12000 29474
rect 9305 29416 9310 29472
rect 9366 29416 12000 29472
rect 9305 29414 12000 29416
rect 9305 29411 9371 29414
rect 4207 29408 4527 29409
rect 0 29338 800 29368
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 29343 4527 29344
rect 7471 29408 7791 29409
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 11200 29384 12000 29414
rect 7471 29343 7791 29344
rect 1577 29338 1643 29341
rect 0 29336 1643 29338
rect 0 29280 1582 29336
rect 1638 29280 1643 29336
rect 0 29278 1643 29280
rect 0 29248 800 29278
rect 1577 29275 1643 29278
rect 9857 29338 9923 29341
rect 10910 29338 10916 29340
rect 9857 29336 10916 29338
rect 9857 29280 9862 29336
rect 9918 29280 10916 29336
rect 9857 29278 10916 29280
rect 9857 29275 9923 29278
rect 10910 29276 10916 29278
rect 10980 29276 10986 29340
rect 9121 29066 9187 29069
rect 11200 29066 12000 29096
rect 9121 29064 12000 29066
rect 9121 29008 9126 29064
rect 9182 29008 12000 29064
rect 9121 29006 12000 29008
rect 9121 29003 9187 29006
rect 11200 28976 12000 29006
rect 2576 28864 2896 28865
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 28799 2896 28800
rect 5839 28864 6159 28865
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 28799 6159 28800
rect 9103 28864 9423 28865
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 28799 9423 28800
rect 0 28658 800 28688
rect 1577 28658 1643 28661
rect 0 28656 1643 28658
rect 0 28600 1582 28656
rect 1638 28600 1643 28656
rect 0 28598 1643 28600
rect 0 28568 800 28598
rect 1577 28595 1643 28598
rect 10041 28522 10107 28525
rect 11200 28522 12000 28552
rect 10041 28520 12000 28522
rect 10041 28464 10046 28520
rect 10102 28464 12000 28520
rect 10041 28462 12000 28464
rect 10041 28459 10107 28462
rect 11200 28432 12000 28462
rect 4207 28320 4527 28321
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 28255 4527 28256
rect 7471 28320 7791 28321
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 28255 7791 28256
rect 10225 28250 10291 28253
rect 10358 28250 10364 28252
rect 10225 28248 10364 28250
rect 10225 28192 10230 28248
rect 10286 28192 10364 28248
rect 10225 28190 10364 28192
rect 10225 28187 10291 28190
rect 10358 28188 10364 28190
rect 10428 28188 10434 28252
rect 0 28114 800 28144
rect 1577 28114 1643 28117
rect 0 28112 1643 28114
rect 0 28056 1582 28112
rect 1638 28056 1643 28112
rect 0 28054 1643 28056
rect 0 28024 800 28054
rect 1577 28051 1643 28054
rect 9305 28114 9371 28117
rect 11200 28114 12000 28144
rect 9305 28112 12000 28114
rect 9305 28056 9310 28112
rect 9366 28056 12000 28112
rect 9305 28054 12000 28056
rect 9305 28051 9371 28054
rect 11200 28024 12000 28054
rect 2576 27776 2896 27777
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 27711 2896 27712
rect 5839 27776 6159 27777
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 27711 6159 27712
rect 9103 27776 9423 27777
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 27711 9423 27712
rect 10133 27570 10199 27573
rect 11200 27570 12000 27600
rect 10133 27568 12000 27570
rect 10133 27512 10138 27568
rect 10194 27512 12000 27568
rect 10133 27510 12000 27512
rect 10133 27507 10199 27510
rect 11200 27480 12000 27510
rect 0 27434 800 27464
rect 1577 27434 1643 27437
rect 0 27432 1643 27434
rect 0 27376 1582 27432
rect 1638 27376 1643 27432
rect 0 27374 1643 27376
rect 0 27344 800 27374
rect 1577 27371 1643 27374
rect 4207 27232 4527 27233
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 27167 4527 27168
rect 7471 27232 7791 27233
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 27167 7791 27168
rect 10041 27162 10107 27165
rect 11200 27162 12000 27192
rect 10041 27160 12000 27162
rect 10041 27104 10046 27160
rect 10102 27104 12000 27160
rect 10041 27102 12000 27104
rect 10041 27099 10107 27102
rect 11200 27072 12000 27102
rect 0 26754 800 26784
rect 1577 26754 1643 26757
rect 0 26752 1643 26754
rect 0 26696 1582 26752
rect 1638 26696 1643 26752
rect 0 26694 1643 26696
rect 0 26664 800 26694
rect 1577 26691 1643 26694
rect 2576 26688 2896 26689
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 26623 2896 26624
rect 5839 26688 6159 26689
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 26623 6159 26624
rect 9103 26688 9423 26689
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 26623 9423 26624
rect 10133 26618 10199 26621
rect 11200 26618 12000 26648
rect 10133 26616 12000 26618
rect 10133 26560 10138 26616
rect 10194 26560 12000 26616
rect 10133 26558 12000 26560
rect 10133 26555 10199 26558
rect 11200 26528 12000 26558
rect 10041 26210 10107 26213
rect 11200 26210 12000 26240
rect 10041 26208 12000 26210
rect 10041 26152 10046 26208
rect 10102 26152 12000 26208
rect 10041 26150 12000 26152
rect 10041 26147 10107 26150
rect 4207 26144 4527 26145
rect 0 26074 800 26104
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 26079 4527 26080
rect 7471 26144 7791 26145
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 11200 26120 12000 26150
rect 7471 26079 7791 26080
rect 1577 26074 1643 26077
rect 0 26072 1643 26074
rect 0 26016 1582 26072
rect 1638 26016 1643 26072
rect 0 26014 1643 26016
rect 0 25984 800 26014
rect 1577 26011 1643 26014
rect 9489 25666 9555 25669
rect 11200 25666 12000 25696
rect 9489 25664 12000 25666
rect 9489 25608 9494 25664
rect 9550 25608 12000 25664
rect 9489 25606 12000 25608
rect 9489 25603 9555 25606
rect 2576 25600 2896 25601
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 25535 2896 25536
rect 5839 25600 6159 25601
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 25535 6159 25536
rect 9103 25600 9423 25601
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 11200 25576 12000 25606
rect 9103 25535 9423 25536
rect 0 25394 800 25424
rect 1577 25394 1643 25397
rect 0 25392 1643 25394
rect 0 25336 1582 25392
rect 1638 25336 1643 25392
rect 0 25334 1643 25336
rect 0 25304 800 25334
rect 1577 25331 1643 25334
rect 10961 25258 11027 25261
rect 11200 25258 12000 25288
rect 10961 25256 12000 25258
rect 10961 25200 10966 25256
rect 11022 25200 12000 25256
rect 10961 25198 12000 25200
rect 10961 25195 11027 25198
rect 11200 25168 12000 25198
rect 4207 25056 4527 25057
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 24991 4527 24992
rect 7471 25056 7791 25057
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 24991 7791 24992
rect 0 24714 800 24744
rect 1577 24714 1643 24717
rect 0 24712 1643 24714
rect 0 24656 1582 24712
rect 1638 24656 1643 24712
rect 0 24654 1643 24656
rect 0 24624 800 24654
rect 1577 24651 1643 24654
rect 9857 24714 9923 24717
rect 11200 24714 12000 24744
rect 9857 24712 12000 24714
rect 9857 24656 9862 24712
rect 9918 24656 12000 24712
rect 9857 24654 12000 24656
rect 9857 24651 9923 24654
rect 11200 24624 12000 24654
rect 2576 24512 2896 24513
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2576 24447 2896 24448
rect 5839 24512 6159 24513
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 24447 6159 24448
rect 9103 24512 9423 24513
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 24447 9423 24448
rect 9489 24306 9555 24309
rect 11200 24306 12000 24336
rect 9489 24304 12000 24306
rect 9489 24248 9494 24304
rect 9550 24248 12000 24304
rect 9489 24246 12000 24248
rect 9489 24243 9555 24246
rect 11200 24216 12000 24246
rect 0 24034 800 24064
rect 1577 24034 1643 24037
rect 0 24032 1643 24034
rect 0 23976 1582 24032
rect 1638 23976 1643 24032
rect 0 23974 1643 23976
rect 0 23944 800 23974
rect 1577 23971 1643 23974
rect 4207 23968 4527 23969
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 23903 4527 23904
rect 7471 23968 7791 23969
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 23903 7791 23904
rect 9121 23762 9187 23765
rect 11200 23762 12000 23792
rect 9121 23760 12000 23762
rect 9121 23704 9126 23760
rect 9182 23704 12000 23760
rect 9121 23702 12000 23704
rect 9121 23699 9187 23702
rect 11200 23672 12000 23702
rect 0 23490 800 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 800 23430
rect 1577 23427 1643 23430
rect 2576 23424 2896 23425
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 23359 2896 23360
rect 5839 23424 6159 23425
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 23359 6159 23360
rect 9103 23424 9423 23425
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 23359 9423 23360
rect 9949 23354 10015 23357
rect 11200 23354 12000 23384
rect 9949 23352 12000 23354
rect 9949 23296 9954 23352
rect 10010 23296 12000 23352
rect 9949 23294 12000 23296
rect 9949 23291 10015 23294
rect 11200 23264 12000 23294
rect 8753 22946 8819 22949
rect 11200 22946 12000 22976
rect 8753 22944 12000 22946
rect 8753 22888 8758 22944
rect 8814 22888 12000 22944
rect 8753 22886 12000 22888
rect 8753 22883 8819 22886
rect 4207 22880 4527 22881
rect 0 22810 800 22840
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 22815 4527 22816
rect 7471 22880 7791 22881
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 11200 22856 12000 22886
rect 7471 22815 7791 22816
rect 1577 22810 1643 22813
rect 0 22808 1643 22810
rect 0 22752 1582 22808
rect 1638 22752 1643 22808
rect 0 22750 1643 22752
rect 0 22720 800 22750
rect 1577 22747 1643 22750
rect 10041 22402 10107 22405
rect 11200 22402 12000 22432
rect 10041 22400 12000 22402
rect 10041 22344 10046 22400
rect 10102 22344 12000 22400
rect 10041 22342 12000 22344
rect 10041 22339 10107 22342
rect 2576 22336 2896 22337
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 22271 2896 22272
rect 5839 22336 6159 22337
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 22271 6159 22272
rect 9103 22336 9423 22337
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 11200 22312 12000 22342
rect 9103 22271 9423 22272
rect 10961 22268 11027 22269
rect 10910 22266 10916 22268
rect 10870 22206 10916 22266
rect 10980 22264 11027 22268
rect 11022 22208 11027 22264
rect 10910 22204 10916 22206
rect 10980 22204 11027 22208
rect 10961 22203 11027 22204
rect 0 22130 800 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 800 22070
rect 1577 22067 1643 22070
rect 8109 21994 8175 21997
rect 11200 21994 12000 22024
rect 8109 21992 12000 21994
rect 8109 21936 8114 21992
rect 8170 21936 12000 21992
rect 8109 21934 12000 21936
rect 8109 21931 8175 21934
rect 11200 21904 12000 21934
rect 4207 21792 4527 21793
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 21727 4527 21728
rect 7471 21792 7791 21793
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 21727 7791 21728
rect 0 21450 800 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 800 21390
rect 1577 21387 1643 21390
rect 9305 21450 9371 21453
rect 11200 21450 12000 21480
rect 9305 21448 12000 21450
rect 9305 21392 9310 21448
rect 9366 21392 12000 21448
rect 9305 21390 12000 21392
rect 9305 21387 9371 21390
rect 11200 21360 12000 21390
rect 2576 21248 2896 21249
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 21183 2896 21184
rect 5839 21248 6159 21249
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 21183 6159 21184
rect 9103 21248 9423 21249
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 21183 9423 21184
rect 9489 21042 9555 21045
rect 11200 21042 12000 21072
rect 9489 21040 12000 21042
rect 9489 20984 9494 21040
rect 9550 20984 12000 21040
rect 9489 20982 12000 20984
rect 9489 20979 9555 20982
rect 11200 20952 12000 20982
rect 0 20770 800 20800
rect 1577 20770 1643 20773
rect 0 20768 1643 20770
rect 0 20712 1582 20768
rect 1638 20712 1643 20768
rect 0 20710 1643 20712
rect 0 20680 800 20710
rect 1577 20707 1643 20710
rect 4207 20704 4527 20705
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 20639 4527 20640
rect 7471 20704 7791 20705
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 20639 7791 20640
rect 9305 20498 9371 20501
rect 11200 20498 12000 20528
rect 9305 20496 12000 20498
rect 9305 20440 9310 20496
rect 9366 20440 12000 20496
rect 9305 20438 12000 20440
rect 9305 20435 9371 20438
rect 11200 20408 12000 20438
rect 8109 20362 8175 20365
rect 8109 20360 9874 20362
rect 8109 20304 8114 20360
rect 8170 20304 9874 20360
rect 8109 20302 9874 20304
rect 8109 20299 8175 20302
rect 2576 20160 2896 20161
rect 0 20090 800 20120
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 20095 2896 20096
rect 5839 20160 6159 20161
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 20095 6159 20096
rect 9103 20160 9423 20161
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 20095 9423 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 9814 20090 9874 20302
rect 11200 20090 12000 20120
rect 9814 20030 12000 20090
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 11200 20000 12000 20030
rect 4207 19616 4527 19617
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 19551 4527 19552
rect 7471 19616 7791 19617
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 19551 7791 19552
rect 8109 19546 8175 19549
rect 11200 19546 12000 19576
rect 8109 19544 12000 19546
rect 8109 19488 8114 19544
rect 8170 19488 12000 19544
rect 8109 19486 12000 19488
rect 8109 19483 8175 19486
rect 11200 19456 12000 19486
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 9581 19138 9647 19141
rect 11200 19138 12000 19168
rect 9581 19136 12000 19138
rect 9581 19080 9586 19136
rect 9642 19080 12000 19136
rect 9581 19078 12000 19080
rect 9581 19075 9647 19078
rect 2576 19072 2896 19073
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 19007 2896 19008
rect 5839 19072 6159 19073
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 19007 6159 19008
rect 9103 19072 9423 19073
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 11200 19048 12000 19078
rect 9103 19007 9423 19008
rect 0 18866 800 18896
rect 1577 18866 1643 18869
rect 0 18864 1643 18866
rect 0 18808 1582 18864
rect 1638 18808 1643 18864
rect 0 18806 1643 18808
rect 0 18776 800 18806
rect 1577 18803 1643 18806
rect 8293 18594 8359 18597
rect 11200 18594 12000 18624
rect 8293 18592 12000 18594
rect 8293 18536 8298 18592
rect 8354 18536 12000 18592
rect 8293 18534 12000 18536
rect 8293 18531 8359 18534
rect 4207 18528 4527 18529
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 18463 4527 18464
rect 7471 18528 7791 18529
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 11200 18504 12000 18534
rect 7471 18463 7791 18464
rect 8385 18458 8451 18461
rect 8886 18458 8892 18460
rect 8385 18456 8892 18458
rect 8385 18400 8390 18456
rect 8446 18400 8892 18456
rect 8385 18398 8892 18400
rect 8385 18395 8451 18398
rect 8886 18396 8892 18398
rect 8956 18396 8962 18460
rect 0 18186 800 18216
rect 1577 18186 1643 18189
rect 0 18184 1643 18186
rect 0 18128 1582 18184
rect 1638 18128 1643 18184
rect 0 18126 1643 18128
rect 0 18096 800 18126
rect 1577 18123 1643 18126
rect 7833 18186 7899 18189
rect 11200 18186 12000 18216
rect 7833 18184 12000 18186
rect 7833 18128 7838 18184
rect 7894 18128 12000 18184
rect 7833 18126 12000 18128
rect 7833 18123 7899 18126
rect 11200 18096 12000 18126
rect 2576 17984 2896 17985
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 17919 2896 17920
rect 5839 17984 6159 17985
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 17919 6159 17920
rect 9103 17984 9423 17985
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 17919 9423 17920
rect 8661 17642 8727 17645
rect 11200 17642 12000 17672
rect 8661 17640 12000 17642
rect 8661 17584 8666 17640
rect 8722 17584 12000 17640
rect 8661 17582 12000 17584
rect 8661 17579 8727 17582
rect 11200 17552 12000 17582
rect 0 17506 800 17536
rect 1577 17506 1643 17509
rect 0 17504 1643 17506
rect 0 17448 1582 17504
rect 1638 17448 1643 17504
rect 0 17446 1643 17448
rect 0 17416 800 17446
rect 1577 17443 1643 17446
rect 4207 17440 4527 17441
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 17375 4527 17376
rect 7471 17440 7791 17441
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 17375 7791 17376
rect 7925 17234 7991 17237
rect 11200 17234 12000 17264
rect 7925 17232 12000 17234
rect 7925 17176 7930 17232
rect 7986 17176 12000 17232
rect 7925 17174 12000 17176
rect 7925 17171 7991 17174
rect 11200 17144 12000 17174
rect 2576 16896 2896 16897
rect 0 16826 800 16856
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 16831 2896 16832
rect 5839 16896 6159 16897
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 16831 6159 16832
rect 9103 16896 9423 16897
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 16831 9423 16832
rect 1577 16826 1643 16829
rect 0 16824 1643 16826
rect 0 16768 1582 16824
rect 1638 16768 1643 16824
rect 0 16766 1643 16768
rect 0 16736 800 16766
rect 1577 16763 1643 16766
rect 7281 16690 7347 16693
rect 11200 16690 12000 16720
rect 7281 16688 12000 16690
rect 7281 16632 7286 16688
rect 7342 16632 12000 16688
rect 7281 16630 12000 16632
rect 7281 16627 7347 16630
rect 11200 16600 12000 16630
rect 4207 16352 4527 16353
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 16287 4527 16288
rect 7471 16352 7791 16353
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 16287 7791 16288
rect 11053 16282 11119 16285
rect 11200 16282 12000 16312
rect 11053 16280 12000 16282
rect 11053 16224 11058 16280
rect 11114 16224 12000 16280
rect 11053 16222 12000 16224
rect 11053 16219 11119 16222
rect 11200 16192 12000 16222
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 6913 16010 6979 16013
rect 6913 16008 9690 16010
rect 6913 15952 6918 16008
rect 6974 15952 9690 16008
rect 6913 15950 9690 15952
rect 6913 15947 6979 15950
rect 2576 15808 2896 15809
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 15743 2896 15744
rect 5839 15808 6159 15809
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 15743 6159 15744
rect 9103 15808 9423 15809
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 15743 9423 15744
rect 9630 15738 9690 15950
rect 11200 15738 12000 15768
rect 9630 15678 12000 15738
rect 11200 15648 12000 15678
rect 0 15466 800 15496
rect 1577 15466 1643 15469
rect 0 15464 1643 15466
rect 0 15408 1582 15464
rect 1638 15408 1643 15464
rect 0 15406 1643 15408
rect 0 15376 800 15406
rect 1577 15403 1643 15406
rect 7097 15466 7163 15469
rect 7097 15464 8034 15466
rect 7097 15408 7102 15464
rect 7158 15408 8034 15464
rect 7097 15406 8034 15408
rect 7097 15403 7163 15406
rect 7974 15330 8034 15406
rect 11200 15330 12000 15360
rect 7974 15270 12000 15330
rect 4207 15264 4527 15265
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 15199 4527 15200
rect 7471 15264 7791 15265
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 11200 15240 12000 15270
rect 7471 15199 7791 15200
rect 7925 15194 7991 15197
rect 8845 15194 8911 15197
rect 7925 15192 8911 15194
rect 7925 15136 7930 15192
rect 7986 15136 8850 15192
rect 8906 15136 8911 15192
rect 7925 15134 8911 15136
rect 7925 15131 7991 15134
rect 8845 15131 8911 15134
rect 6913 14922 6979 14925
rect 6913 14920 9690 14922
rect 6913 14864 6918 14920
rect 6974 14864 9690 14920
rect 6913 14862 9690 14864
rect 6913 14859 6979 14862
rect 0 14786 800 14816
rect 1577 14786 1643 14789
rect 0 14784 1643 14786
rect 0 14728 1582 14784
rect 1638 14728 1643 14784
rect 0 14726 1643 14728
rect 0 14696 800 14726
rect 1577 14723 1643 14726
rect 6361 14786 6427 14789
rect 8293 14786 8359 14789
rect 6361 14784 8359 14786
rect 6361 14728 6366 14784
rect 6422 14728 8298 14784
rect 8354 14728 8359 14784
rect 6361 14726 8359 14728
rect 9630 14786 9690 14862
rect 11200 14786 12000 14816
rect 9630 14726 12000 14786
rect 6361 14723 6427 14726
rect 8293 14723 8359 14726
rect 2576 14720 2896 14721
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 14655 2896 14656
rect 5839 14720 6159 14721
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 14655 6159 14656
rect 9103 14720 9423 14721
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 11200 14696 12000 14726
rect 9103 14655 9423 14656
rect 7281 14652 7347 14653
rect 7230 14650 7236 14652
rect 7190 14590 7236 14650
rect 7300 14648 7347 14652
rect 7342 14592 7347 14648
rect 7230 14588 7236 14590
rect 7300 14588 7347 14592
rect 7281 14587 7347 14588
rect 6177 14514 6243 14517
rect 7649 14514 7715 14517
rect 6177 14512 7715 14514
rect 6177 14456 6182 14512
rect 6238 14456 7654 14512
rect 7710 14456 7715 14512
rect 6177 14454 7715 14456
rect 6177 14451 6243 14454
rect 7649 14451 7715 14454
rect 7189 14378 7255 14381
rect 11200 14378 12000 14408
rect 7189 14376 12000 14378
rect 7189 14320 7194 14376
rect 7250 14320 12000 14376
rect 7189 14318 12000 14320
rect 7189 14315 7255 14318
rect 11200 14288 12000 14318
rect 0 14242 800 14272
rect 1577 14242 1643 14245
rect 0 14240 1643 14242
rect 0 14184 1582 14240
rect 1638 14184 1643 14240
rect 0 14182 1643 14184
rect 0 14152 800 14182
rect 1577 14179 1643 14182
rect 4207 14176 4527 14177
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 14111 4527 14112
rect 7471 14176 7791 14177
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 14111 7791 14112
rect 7097 13970 7163 13973
rect 8385 13970 8451 13973
rect 7097 13968 8451 13970
rect 7097 13912 7102 13968
rect 7158 13912 8390 13968
rect 8446 13912 8451 13968
rect 7097 13910 8451 13912
rect 7097 13907 7163 13910
rect 8385 13907 8451 13910
rect 6913 13834 6979 13837
rect 11200 13834 12000 13864
rect 6913 13832 12000 13834
rect 6913 13776 6918 13832
rect 6974 13776 12000 13832
rect 6913 13774 12000 13776
rect 6913 13771 6979 13774
rect 11200 13744 12000 13774
rect 2576 13632 2896 13633
rect 0 13562 800 13592
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 13567 2896 13568
rect 5839 13632 6159 13633
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 13567 6159 13568
rect 9103 13632 9423 13633
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 13567 9423 13568
rect 1577 13562 1643 13565
rect 0 13560 1643 13562
rect 0 13504 1582 13560
rect 1638 13504 1643 13560
rect 0 13502 1643 13504
rect 0 13472 800 13502
rect 1577 13499 1643 13502
rect 7230 13500 7236 13564
rect 7300 13562 7306 13564
rect 7649 13562 7715 13565
rect 7300 13560 7715 13562
rect 7300 13504 7654 13560
rect 7710 13504 7715 13560
rect 7300 13502 7715 13504
rect 7300 13500 7306 13502
rect 5349 13426 5415 13429
rect 7238 13426 7298 13500
rect 7649 13499 7715 13502
rect 5349 13424 7298 13426
rect 5349 13368 5354 13424
rect 5410 13368 7298 13424
rect 5349 13366 7298 13368
rect 8109 13426 8175 13429
rect 11200 13426 12000 13456
rect 8109 13424 12000 13426
rect 8109 13368 8114 13424
rect 8170 13368 12000 13424
rect 8109 13366 12000 13368
rect 5349 13363 5415 13366
rect 4207 13088 4527 13089
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 13023 4527 13024
rect 6318 13021 6378 13366
rect 8109 13363 8175 13366
rect 11200 13336 12000 13366
rect 7471 13088 7791 13089
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 13023 7791 13024
rect 6269 13016 6378 13021
rect 6269 12960 6274 13016
rect 6330 12960 6378 13016
rect 6269 12958 6378 12960
rect 6269 12955 6335 12958
rect 0 12882 800 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 800 12822
rect 1577 12819 1643 12822
rect 7189 12882 7255 12885
rect 11200 12882 12000 12912
rect 7189 12880 12000 12882
rect 7189 12824 7194 12880
rect 7250 12824 12000 12880
rect 7189 12822 12000 12824
rect 7189 12819 7255 12822
rect 11200 12792 12000 12822
rect 6913 12746 6979 12749
rect 6913 12744 9690 12746
rect 6913 12688 6918 12744
rect 6974 12688 9690 12744
rect 6913 12686 9690 12688
rect 6913 12683 6979 12686
rect 2576 12544 2896 12545
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 12479 2896 12480
rect 5839 12544 6159 12545
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 12479 6159 12480
rect 9103 12544 9423 12545
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 12479 9423 12480
rect 9630 12474 9690 12686
rect 11200 12474 12000 12504
rect 9630 12414 12000 12474
rect 11200 12384 12000 12414
rect 0 12202 800 12232
rect 1577 12202 1643 12205
rect 0 12200 1643 12202
rect 0 12144 1582 12200
rect 1638 12144 1643 12200
rect 0 12142 1643 12144
rect 0 12112 800 12142
rect 1577 12139 1643 12142
rect 5901 12202 5967 12205
rect 5901 12200 9690 12202
rect 5901 12144 5906 12200
rect 5962 12144 9690 12200
rect 5901 12142 9690 12144
rect 5901 12139 5967 12142
rect 4207 12000 4527 12001
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 11935 4527 11936
rect 7471 12000 7791 12001
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 11935 7791 11936
rect 9630 11930 9690 12142
rect 11200 11930 12000 11960
rect 9630 11870 12000 11930
rect 11200 11840 12000 11870
rect 0 11522 800 11552
rect 1577 11522 1643 11525
rect 11200 11522 12000 11552
rect 0 11520 1643 11522
rect 0 11464 1582 11520
rect 1638 11464 1643 11520
rect 0 11462 1643 11464
rect 0 11432 800 11462
rect 1577 11459 1643 11462
rect 9584 11462 12000 11522
rect 2576 11456 2896 11457
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5839 11456 6159 11457
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 11391 6159 11392
rect 9103 11456 9423 11457
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 11391 9423 11392
rect 7281 11250 7347 11253
rect 9584 11250 9644 11462
rect 11200 11432 12000 11462
rect 7281 11248 9644 11250
rect 7281 11192 7286 11248
rect 7342 11192 9644 11248
rect 7281 11190 9644 11192
rect 7281 11187 7347 11190
rect 8385 11114 8451 11117
rect 11200 11114 12000 11144
rect 8385 11112 12000 11114
rect 8385 11056 8390 11112
rect 8446 11056 12000 11112
rect 8385 11054 12000 11056
rect 8385 11051 8451 11054
rect 11200 11024 12000 11054
rect 4207 10912 4527 10913
rect 0 10842 800 10872
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 10847 4527 10848
rect 7471 10912 7791 10913
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 10847 7791 10848
rect 1577 10842 1643 10845
rect 0 10840 1643 10842
rect 0 10784 1582 10840
rect 1638 10784 1643 10840
rect 0 10782 1643 10784
rect 0 10752 800 10782
rect 1577 10779 1643 10782
rect 8017 10570 8083 10573
rect 11200 10570 12000 10600
rect 8017 10568 12000 10570
rect 8017 10512 8022 10568
rect 8078 10512 12000 10568
rect 8017 10510 12000 10512
rect 8017 10507 8083 10510
rect 11200 10480 12000 10510
rect 2576 10368 2896 10369
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5839 10368 6159 10369
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 10303 6159 10304
rect 9103 10368 9423 10369
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 10303 9423 10304
rect 0 10162 800 10192
rect 1577 10162 1643 10165
rect 0 10160 1643 10162
rect 0 10104 1582 10160
rect 1638 10104 1643 10160
rect 0 10102 1643 10104
rect 0 10072 800 10102
rect 1577 10099 1643 10102
rect 8886 10100 8892 10164
rect 8956 10162 8962 10164
rect 9213 10162 9279 10165
rect 8956 10160 9279 10162
rect 8956 10104 9218 10160
rect 9274 10104 9279 10160
rect 8956 10102 9279 10104
rect 8956 10100 8962 10102
rect 9213 10099 9279 10102
rect 10409 10162 10475 10165
rect 11200 10162 12000 10192
rect 10409 10160 12000 10162
rect 10409 10104 10414 10160
rect 10470 10104 12000 10160
rect 10409 10102 12000 10104
rect 10409 10099 10475 10102
rect 11200 10072 12000 10102
rect 4207 9824 4527 9825
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 9759 4527 9760
rect 7471 9824 7791 9825
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 9759 7791 9760
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 9765 9618 9831 9621
rect 11200 9618 12000 9648
rect 9765 9616 12000 9618
rect 9765 9560 9770 9616
rect 9826 9560 12000 9616
rect 9765 9558 12000 9560
rect 9765 9555 9831 9558
rect 11200 9528 12000 9558
rect 7833 9482 7899 9485
rect 7833 9480 9644 9482
rect 7833 9424 7838 9480
rect 7894 9424 9644 9480
rect 7833 9422 9644 9424
rect 7833 9419 7899 9422
rect 2576 9280 2896 9281
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5839 9280 6159 9281
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 9215 6159 9216
rect 9103 9280 9423 9281
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 9215 9423 9216
rect 9584 9210 9644 9422
rect 11200 9210 12000 9240
rect 9584 9150 12000 9210
rect 11200 9120 12000 9150
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 4207 8736 4527 8737
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 8671 4527 8672
rect 7471 8736 7791 8737
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 8671 7791 8672
rect 9121 8666 9187 8669
rect 11200 8666 12000 8696
rect 9121 8664 12000 8666
rect 9121 8608 9126 8664
rect 9182 8608 12000 8664
rect 9121 8606 12000 8608
rect 9121 8603 9187 8606
rect 11200 8576 12000 8606
rect 0 8258 800 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 800 8198
rect 1577 8195 1643 8198
rect 9857 8258 9923 8261
rect 11200 8258 12000 8288
rect 9857 8256 12000 8258
rect 9857 8200 9862 8256
rect 9918 8200 12000 8256
rect 9857 8198 12000 8200
rect 9857 8195 9923 8198
rect 2576 8192 2896 8193
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5839 8192 6159 8193
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 8127 6159 8128
rect 9103 8192 9423 8193
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 11200 8168 12000 8198
rect 9103 8127 9423 8128
rect 10225 7714 10291 7717
rect 11200 7714 12000 7744
rect 10225 7712 12000 7714
rect 10225 7656 10230 7712
rect 10286 7656 12000 7712
rect 10225 7654 12000 7656
rect 10225 7651 10291 7654
rect 4207 7648 4527 7649
rect 0 7578 800 7608
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 7583 4527 7584
rect 7471 7648 7791 7649
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 11200 7624 12000 7654
rect 7471 7583 7791 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 8937 7306 9003 7309
rect 11200 7306 12000 7336
rect 8937 7304 12000 7306
rect 8937 7248 8942 7304
rect 8998 7248 12000 7304
rect 8937 7246 12000 7248
rect 8937 7243 9003 7246
rect 11200 7216 12000 7246
rect 2576 7104 2896 7105
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5839 7104 6159 7105
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 7039 6159 7040
rect 9103 7104 9423 7105
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 7039 9423 7040
rect 0 6898 800 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 800 6838
rect 1577 6835 1643 6838
rect 10961 6762 11027 6765
rect 11200 6762 12000 6792
rect 10961 6760 12000 6762
rect 10961 6704 10966 6760
rect 11022 6704 12000 6760
rect 10961 6702 12000 6704
rect 10961 6699 11027 6702
rect 11200 6672 12000 6702
rect 4207 6560 4527 6561
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 6495 4527 6496
rect 7471 6560 7791 6561
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 6495 7791 6496
rect 9765 6354 9831 6357
rect 11200 6354 12000 6384
rect 9765 6352 12000 6354
rect 9765 6296 9770 6352
rect 9826 6296 12000 6352
rect 9765 6294 12000 6296
rect 9765 6291 9831 6294
rect 11200 6264 12000 6294
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 2576 6016 2896 6017
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5839 6016 6159 6017
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 5951 6159 5952
rect 9103 6016 9423 6017
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 5951 9423 5952
rect 11200 5720 12000 5840
rect 0 5538 800 5568
rect 1577 5538 1643 5541
rect 0 5536 1643 5538
rect 0 5480 1582 5536
rect 1638 5480 1643 5536
rect 0 5478 1643 5480
rect 0 5448 800 5478
rect 1577 5475 1643 5478
rect 4207 5472 4527 5473
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 5407 4527 5408
rect 7471 5472 7791 5473
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 5407 7791 5408
rect 11200 5312 12000 5432
rect 8109 5130 8175 5133
rect 8109 5128 9874 5130
rect 8109 5072 8114 5128
rect 8170 5072 9874 5128
rect 8109 5070 9874 5072
rect 8109 5067 8175 5070
rect 0 4994 800 5024
rect 1577 4994 1643 4997
rect 0 4992 1643 4994
rect 0 4936 1582 4992
rect 1638 4936 1643 4992
rect 0 4934 1643 4936
rect 0 4904 800 4934
rect 1577 4931 1643 4934
rect 2576 4928 2896 4929
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5839 4928 6159 4929
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 4863 6159 4864
rect 9103 4928 9423 4929
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 4863 9423 4864
rect 9814 4858 9874 5070
rect 11200 4858 12000 4888
rect 9814 4798 12000 4858
rect 11200 4768 12000 4798
rect 8937 4450 9003 4453
rect 11200 4450 12000 4480
rect 8937 4448 12000 4450
rect 8937 4392 8942 4448
rect 8998 4392 12000 4448
rect 8937 4390 12000 4392
rect 8937 4387 9003 4390
rect 4207 4384 4527 4385
rect 0 4314 800 4344
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 4319 4527 4320
rect 7471 4384 7791 4385
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 11200 4360 12000 4390
rect 7471 4319 7791 4320
rect 1577 4314 1643 4317
rect 0 4312 1643 4314
rect 0 4256 1582 4312
rect 1638 4256 1643 4312
rect 0 4254 1643 4256
rect 0 4224 800 4254
rect 1577 4251 1643 4254
rect 9121 4042 9187 4045
rect 9121 4040 10058 4042
rect 9121 3984 9126 4040
rect 9182 3984 10058 4040
rect 9121 3982 10058 3984
rect 9121 3979 9187 3982
rect 9998 3906 10058 3982
rect 11200 3906 12000 3936
rect 9998 3846 12000 3906
rect 2576 3840 2896 3841
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5839 3840 6159 3841
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 3775 6159 3776
rect 9103 3840 9423 3841
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 11200 3816 12000 3846
rect 9103 3775 9423 3776
rect 0 3634 800 3664
rect 1577 3634 1643 3637
rect 0 3632 1643 3634
rect 0 3576 1582 3632
rect 1638 3576 1643 3632
rect 0 3574 1643 3576
rect 0 3544 800 3574
rect 1577 3571 1643 3574
rect 8109 3498 8175 3501
rect 11200 3498 12000 3528
rect 8109 3496 12000 3498
rect 8109 3440 8114 3496
rect 8170 3440 12000 3496
rect 8109 3438 12000 3440
rect 8109 3435 8175 3438
rect 11200 3408 12000 3438
rect 4207 3296 4527 3297
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 3231 4527 3232
rect 7471 3296 7791 3297
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 7471 3231 7791 3232
rect 0 2954 800 2984
rect 1577 2954 1643 2957
rect 0 2952 1643 2954
rect 0 2896 1582 2952
rect 1638 2896 1643 2952
rect 0 2894 1643 2896
rect 0 2864 800 2894
rect 1577 2891 1643 2894
rect 7833 2954 7899 2957
rect 11200 2954 12000 2984
rect 7833 2952 12000 2954
rect 7833 2896 7838 2952
rect 7894 2896 12000 2952
rect 7833 2894 12000 2896
rect 7833 2891 7899 2894
rect 11200 2864 12000 2894
rect 2576 2752 2896 2753
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5839 2752 6159 2753
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2687 6159 2688
rect 9103 2752 9423 2753
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2687 9423 2688
rect 9581 2546 9647 2549
rect 11200 2546 12000 2576
rect 9581 2544 12000 2546
rect 9581 2488 9586 2544
rect 9642 2488 12000 2544
rect 9581 2486 12000 2488
rect 9581 2483 9647 2486
rect 11200 2456 12000 2486
rect 0 2274 800 2304
rect 2313 2274 2379 2277
rect 0 2272 2379 2274
rect 0 2216 2318 2272
rect 2374 2216 2379 2272
rect 0 2214 2379 2216
rect 0 2184 800 2214
rect 2313 2211 2379 2214
rect 4207 2208 4527 2209
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2143 4527 2144
rect 7471 2208 7791 2209
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2143 7791 2144
rect 9489 2002 9555 2005
rect 11200 2002 12000 2032
rect 9489 2000 12000 2002
rect 9489 1944 9494 2000
rect 9550 1944 12000 2000
rect 9489 1942 12000 1944
rect 9489 1939 9555 1942
rect 11200 1912 12000 1942
rect 0 1594 800 1624
rect 1393 1594 1459 1597
rect 0 1592 1459 1594
rect 0 1536 1398 1592
rect 1454 1536 1459 1592
rect 0 1534 1459 1536
rect 0 1504 800 1534
rect 1393 1531 1459 1534
rect 7925 1594 7991 1597
rect 11200 1594 12000 1624
rect 7925 1592 12000 1594
rect 7925 1536 7930 1592
rect 7986 1536 12000 1592
rect 7925 1534 12000 1536
rect 7925 1531 7991 1534
rect 11200 1504 12000 1534
rect 9305 1050 9371 1053
rect 11200 1050 12000 1080
rect 9305 1048 12000 1050
rect 9305 992 9310 1048
rect 9366 992 12000 1048
rect 9305 990 12000 992
rect 9305 987 9371 990
rect 11200 960 12000 990
rect 0 914 800 944
rect 1577 914 1643 917
rect 0 912 1643 914
rect 0 856 1582 912
rect 1638 856 1643 912
rect 0 854 1643 856
rect 0 824 800 854
rect 1577 851 1643 854
rect 8201 642 8267 645
rect 11200 642 12000 672
rect 8201 640 12000 642
rect 8201 584 8206 640
rect 8262 584 12000 640
rect 8201 582 12000 584
rect 8201 579 8267 582
rect 11200 552 12000 582
rect 0 370 800 400
rect 2865 370 2931 373
rect 0 368 2931 370
rect 0 312 2870 368
rect 2926 312 2931 368
rect 0 310 2931 312
rect 0 280 800 310
rect 2865 307 2931 310
rect 8109 234 8175 237
rect 11200 234 12000 264
rect 8109 232 12000 234
rect 8109 176 8114 232
rect 8170 176 12000 232
rect 8109 174 12000 176
rect 8109 171 8175 174
rect 11200 144 12000 174
<< via3 >>
rect 2584 77820 2648 77824
rect 2584 77764 2588 77820
rect 2588 77764 2644 77820
rect 2644 77764 2648 77820
rect 2584 77760 2648 77764
rect 2664 77820 2728 77824
rect 2664 77764 2668 77820
rect 2668 77764 2724 77820
rect 2724 77764 2728 77820
rect 2664 77760 2728 77764
rect 2744 77820 2808 77824
rect 2744 77764 2748 77820
rect 2748 77764 2804 77820
rect 2804 77764 2808 77820
rect 2744 77760 2808 77764
rect 2824 77820 2888 77824
rect 2824 77764 2828 77820
rect 2828 77764 2884 77820
rect 2884 77764 2888 77820
rect 2824 77760 2888 77764
rect 5847 77820 5911 77824
rect 5847 77764 5851 77820
rect 5851 77764 5907 77820
rect 5907 77764 5911 77820
rect 5847 77760 5911 77764
rect 5927 77820 5991 77824
rect 5927 77764 5931 77820
rect 5931 77764 5987 77820
rect 5987 77764 5991 77820
rect 5927 77760 5991 77764
rect 6007 77820 6071 77824
rect 6007 77764 6011 77820
rect 6011 77764 6067 77820
rect 6067 77764 6071 77820
rect 6007 77760 6071 77764
rect 6087 77820 6151 77824
rect 6087 77764 6091 77820
rect 6091 77764 6147 77820
rect 6147 77764 6151 77820
rect 6087 77760 6151 77764
rect 9111 77820 9175 77824
rect 9111 77764 9115 77820
rect 9115 77764 9171 77820
rect 9171 77764 9175 77820
rect 9111 77760 9175 77764
rect 9191 77820 9255 77824
rect 9191 77764 9195 77820
rect 9195 77764 9251 77820
rect 9251 77764 9255 77820
rect 9191 77760 9255 77764
rect 9271 77820 9335 77824
rect 9271 77764 9275 77820
rect 9275 77764 9331 77820
rect 9331 77764 9335 77820
rect 9271 77760 9335 77764
rect 9351 77820 9415 77824
rect 9351 77764 9355 77820
rect 9355 77764 9411 77820
rect 9411 77764 9415 77820
rect 9351 77760 9415 77764
rect 4215 77276 4279 77280
rect 4215 77220 4219 77276
rect 4219 77220 4275 77276
rect 4275 77220 4279 77276
rect 4215 77216 4279 77220
rect 4295 77276 4359 77280
rect 4295 77220 4299 77276
rect 4299 77220 4355 77276
rect 4355 77220 4359 77276
rect 4295 77216 4359 77220
rect 4375 77276 4439 77280
rect 4375 77220 4379 77276
rect 4379 77220 4435 77276
rect 4435 77220 4439 77276
rect 4375 77216 4439 77220
rect 4455 77276 4519 77280
rect 4455 77220 4459 77276
rect 4459 77220 4515 77276
rect 4515 77220 4519 77276
rect 4455 77216 4519 77220
rect 7479 77276 7543 77280
rect 7479 77220 7483 77276
rect 7483 77220 7539 77276
rect 7539 77220 7543 77276
rect 7479 77216 7543 77220
rect 7559 77276 7623 77280
rect 7559 77220 7563 77276
rect 7563 77220 7619 77276
rect 7619 77220 7623 77276
rect 7559 77216 7623 77220
rect 7639 77276 7703 77280
rect 7639 77220 7643 77276
rect 7643 77220 7699 77276
rect 7699 77220 7703 77276
rect 7639 77216 7703 77220
rect 7719 77276 7783 77280
rect 7719 77220 7723 77276
rect 7723 77220 7779 77276
rect 7779 77220 7783 77276
rect 7719 77216 7783 77220
rect 2584 76732 2648 76736
rect 2584 76676 2588 76732
rect 2588 76676 2644 76732
rect 2644 76676 2648 76732
rect 2584 76672 2648 76676
rect 2664 76732 2728 76736
rect 2664 76676 2668 76732
rect 2668 76676 2724 76732
rect 2724 76676 2728 76732
rect 2664 76672 2728 76676
rect 2744 76732 2808 76736
rect 2744 76676 2748 76732
rect 2748 76676 2804 76732
rect 2804 76676 2808 76732
rect 2744 76672 2808 76676
rect 2824 76732 2888 76736
rect 2824 76676 2828 76732
rect 2828 76676 2884 76732
rect 2884 76676 2888 76732
rect 2824 76672 2888 76676
rect 5847 76732 5911 76736
rect 5847 76676 5851 76732
rect 5851 76676 5907 76732
rect 5907 76676 5911 76732
rect 5847 76672 5911 76676
rect 5927 76732 5991 76736
rect 5927 76676 5931 76732
rect 5931 76676 5987 76732
rect 5987 76676 5991 76732
rect 5927 76672 5991 76676
rect 6007 76732 6071 76736
rect 6007 76676 6011 76732
rect 6011 76676 6067 76732
rect 6067 76676 6071 76732
rect 6007 76672 6071 76676
rect 6087 76732 6151 76736
rect 6087 76676 6091 76732
rect 6091 76676 6147 76732
rect 6147 76676 6151 76732
rect 6087 76672 6151 76676
rect 9111 76732 9175 76736
rect 9111 76676 9115 76732
rect 9115 76676 9171 76732
rect 9171 76676 9175 76732
rect 9111 76672 9175 76676
rect 9191 76732 9255 76736
rect 9191 76676 9195 76732
rect 9195 76676 9251 76732
rect 9251 76676 9255 76732
rect 9191 76672 9255 76676
rect 9271 76732 9335 76736
rect 9271 76676 9275 76732
rect 9275 76676 9331 76732
rect 9331 76676 9335 76732
rect 9271 76672 9335 76676
rect 9351 76732 9415 76736
rect 9351 76676 9355 76732
rect 9355 76676 9411 76732
rect 9411 76676 9415 76732
rect 9351 76672 9415 76676
rect 4215 76188 4279 76192
rect 4215 76132 4219 76188
rect 4219 76132 4275 76188
rect 4275 76132 4279 76188
rect 4215 76128 4279 76132
rect 4295 76188 4359 76192
rect 4295 76132 4299 76188
rect 4299 76132 4355 76188
rect 4355 76132 4359 76188
rect 4295 76128 4359 76132
rect 4375 76188 4439 76192
rect 4375 76132 4379 76188
rect 4379 76132 4435 76188
rect 4435 76132 4439 76188
rect 4375 76128 4439 76132
rect 4455 76188 4519 76192
rect 4455 76132 4459 76188
rect 4459 76132 4515 76188
rect 4515 76132 4519 76188
rect 4455 76128 4519 76132
rect 7479 76188 7543 76192
rect 7479 76132 7483 76188
rect 7483 76132 7539 76188
rect 7539 76132 7543 76188
rect 7479 76128 7543 76132
rect 7559 76188 7623 76192
rect 7559 76132 7563 76188
rect 7563 76132 7619 76188
rect 7619 76132 7623 76188
rect 7559 76128 7623 76132
rect 7639 76188 7703 76192
rect 7639 76132 7643 76188
rect 7643 76132 7699 76188
rect 7699 76132 7703 76188
rect 7639 76128 7703 76132
rect 7719 76188 7783 76192
rect 7719 76132 7723 76188
rect 7723 76132 7779 76188
rect 7779 76132 7783 76188
rect 7719 76128 7783 76132
rect 2584 75644 2648 75648
rect 2584 75588 2588 75644
rect 2588 75588 2644 75644
rect 2644 75588 2648 75644
rect 2584 75584 2648 75588
rect 2664 75644 2728 75648
rect 2664 75588 2668 75644
rect 2668 75588 2724 75644
rect 2724 75588 2728 75644
rect 2664 75584 2728 75588
rect 2744 75644 2808 75648
rect 2744 75588 2748 75644
rect 2748 75588 2804 75644
rect 2804 75588 2808 75644
rect 2744 75584 2808 75588
rect 2824 75644 2888 75648
rect 2824 75588 2828 75644
rect 2828 75588 2884 75644
rect 2884 75588 2888 75644
rect 2824 75584 2888 75588
rect 5847 75644 5911 75648
rect 5847 75588 5851 75644
rect 5851 75588 5907 75644
rect 5907 75588 5911 75644
rect 5847 75584 5911 75588
rect 5927 75644 5991 75648
rect 5927 75588 5931 75644
rect 5931 75588 5987 75644
rect 5987 75588 5991 75644
rect 5927 75584 5991 75588
rect 6007 75644 6071 75648
rect 6007 75588 6011 75644
rect 6011 75588 6067 75644
rect 6067 75588 6071 75644
rect 6007 75584 6071 75588
rect 6087 75644 6151 75648
rect 6087 75588 6091 75644
rect 6091 75588 6147 75644
rect 6147 75588 6151 75644
rect 6087 75584 6151 75588
rect 9111 75644 9175 75648
rect 9111 75588 9115 75644
rect 9115 75588 9171 75644
rect 9171 75588 9175 75644
rect 9111 75584 9175 75588
rect 9191 75644 9255 75648
rect 9191 75588 9195 75644
rect 9195 75588 9251 75644
rect 9251 75588 9255 75644
rect 9191 75584 9255 75588
rect 9271 75644 9335 75648
rect 9271 75588 9275 75644
rect 9275 75588 9331 75644
rect 9331 75588 9335 75644
rect 9271 75584 9335 75588
rect 9351 75644 9415 75648
rect 9351 75588 9355 75644
rect 9355 75588 9411 75644
rect 9411 75588 9415 75644
rect 9351 75584 9415 75588
rect 4215 75100 4279 75104
rect 4215 75044 4219 75100
rect 4219 75044 4275 75100
rect 4275 75044 4279 75100
rect 4215 75040 4279 75044
rect 4295 75100 4359 75104
rect 4295 75044 4299 75100
rect 4299 75044 4355 75100
rect 4355 75044 4359 75100
rect 4295 75040 4359 75044
rect 4375 75100 4439 75104
rect 4375 75044 4379 75100
rect 4379 75044 4435 75100
rect 4435 75044 4439 75100
rect 4375 75040 4439 75044
rect 4455 75100 4519 75104
rect 4455 75044 4459 75100
rect 4459 75044 4515 75100
rect 4515 75044 4519 75100
rect 4455 75040 4519 75044
rect 7479 75100 7543 75104
rect 7479 75044 7483 75100
rect 7483 75044 7539 75100
rect 7539 75044 7543 75100
rect 7479 75040 7543 75044
rect 7559 75100 7623 75104
rect 7559 75044 7563 75100
rect 7563 75044 7619 75100
rect 7619 75044 7623 75100
rect 7559 75040 7623 75044
rect 7639 75100 7703 75104
rect 7639 75044 7643 75100
rect 7643 75044 7699 75100
rect 7699 75044 7703 75100
rect 7639 75040 7703 75044
rect 7719 75100 7783 75104
rect 7719 75044 7723 75100
rect 7723 75044 7779 75100
rect 7779 75044 7783 75100
rect 7719 75040 7783 75044
rect 2584 74556 2648 74560
rect 2584 74500 2588 74556
rect 2588 74500 2644 74556
rect 2644 74500 2648 74556
rect 2584 74496 2648 74500
rect 2664 74556 2728 74560
rect 2664 74500 2668 74556
rect 2668 74500 2724 74556
rect 2724 74500 2728 74556
rect 2664 74496 2728 74500
rect 2744 74556 2808 74560
rect 2744 74500 2748 74556
rect 2748 74500 2804 74556
rect 2804 74500 2808 74556
rect 2744 74496 2808 74500
rect 2824 74556 2888 74560
rect 2824 74500 2828 74556
rect 2828 74500 2884 74556
rect 2884 74500 2888 74556
rect 2824 74496 2888 74500
rect 5847 74556 5911 74560
rect 5847 74500 5851 74556
rect 5851 74500 5907 74556
rect 5907 74500 5911 74556
rect 5847 74496 5911 74500
rect 5927 74556 5991 74560
rect 5927 74500 5931 74556
rect 5931 74500 5987 74556
rect 5987 74500 5991 74556
rect 5927 74496 5991 74500
rect 6007 74556 6071 74560
rect 6007 74500 6011 74556
rect 6011 74500 6067 74556
rect 6067 74500 6071 74556
rect 6007 74496 6071 74500
rect 6087 74556 6151 74560
rect 6087 74500 6091 74556
rect 6091 74500 6147 74556
rect 6147 74500 6151 74556
rect 6087 74496 6151 74500
rect 9111 74556 9175 74560
rect 9111 74500 9115 74556
rect 9115 74500 9171 74556
rect 9171 74500 9175 74556
rect 9111 74496 9175 74500
rect 9191 74556 9255 74560
rect 9191 74500 9195 74556
rect 9195 74500 9251 74556
rect 9251 74500 9255 74556
rect 9191 74496 9255 74500
rect 9271 74556 9335 74560
rect 9271 74500 9275 74556
rect 9275 74500 9331 74556
rect 9331 74500 9335 74556
rect 9271 74496 9335 74500
rect 9351 74556 9415 74560
rect 9351 74500 9355 74556
rect 9355 74500 9411 74556
rect 9411 74500 9415 74556
rect 9351 74496 9415 74500
rect 4215 74012 4279 74016
rect 4215 73956 4219 74012
rect 4219 73956 4275 74012
rect 4275 73956 4279 74012
rect 4215 73952 4279 73956
rect 4295 74012 4359 74016
rect 4295 73956 4299 74012
rect 4299 73956 4355 74012
rect 4355 73956 4359 74012
rect 4295 73952 4359 73956
rect 4375 74012 4439 74016
rect 4375 73956 4379 74012
rect 4379 73956 4435 74012
rect 4435 73956 4439 74012
rect 4375 73952 4439 73956
rect 4455 74012 4519 74016
rect 4455 73956 4459 74012
rect 4459 73956 4515 74012
rect 4515 73956 4519 74012
rect 4455 73952 4519 73956
rect 7479 74012 7543 74016
rect 7479 73956 7483 74012
rect 7483 73956 7539 74012
rect 7539 73956 7543 74012
rect 7479 73952 7543 73956
rect 7559 74012 7623 74016
rect 7559 73956 7563 74012
rect 7563 73956 7619 74012
rect 7619 73956 7623 74012
rect 7559 73952 7623 73956
rect 7639 74012 7703 74016
rect 7639 73956 7643 74012
rect 7643 73956 7699 74012
rect 7699 73956 7703 74012
rect 7639 73952 7703 73956
rect 7719 74012 7783 74016
rect 7719 73956 7723 74012
rect 7723 73956 7779 74012
rect 7779 73956 7783 74012
rect 7719 73952 7783 73956
rect 2584 73468 2648 73472
rect 2584 73412 2588 73468
rect 2588 73412 2644 73468
rect 2644 73412 2648 73468
rect 2584 73408 2648 73412
rect 2664 73468 2728 73472
rect 2664 73412 2668 73468
rect 2668 73412 2724 73468
rect 2724 73412 2728 73468
rect 2664 73408 2728 73412
rect 2744 73468 2808 73472
rect 2744 73412 2748 73468
rect 2748 73412 2804 73468
rect 2804 73412 2808 73468
rect 2744 73408 2808 73412
rect 2824 73468 2888 73472
rect 2824 73412 2828 73468
rect 2828 73412 2884 73468
rect 2884 73412 2888 73468
rect 2824 73408 2888 73412
rect 5847 73468 5911 73472
rect 5847 73412 5851 73468
rect 5851 73412 5907 73468
rect 5907 73412 5911 73468
rect 5847 73408 5911 73412
rect 5927 73468 5991 73472
rect 5927 73412 5931 73468
rect 5931 73412 5987 73468
rect 5987 73412 5991 73468
rect 5927 73408 5991 73412
rect 6007 73468 6071 73472
rect 6007 73412 6011 73468
rect 6011 73412 6067 73468
rect 6067 73412 6071 73468
rect 6007 73408 6071 73412
rect 6087 73468 6151 73472
rect 6087 73412 6091 73468
rect 6091 73412 6147 73468
rect 6147 73412 6151 73468
rect 6087 73408 6151 73412
rect 9111 73468 9175 73472
rect 9111 73412 9115 73468
rect 9115 73412 9171 73468
rect 9171 73412 9175 73468
rect 9111 73408 9175 73412
rect 9191 73468 9255 73472
rect 9191 73412 9195 73468
rect 9195 73412 9251 73468
rect 9251 73412 9255 73468
rect 9191 73408 9255 73412
rect 9271 73468 9335 73472
rect 9271 73412 9275 73468
rect 9275 73412 9331 73468
rect 9331 73412 9335 73468
rect 9271 73408 9335 73412
rect 9351 73468 9415 73472
rect 9351 73412 9355 73468
rect 9355 73412 9411 73468
rect 9411 73412 9415 73468
rect 9351 73408 9415 73412
rect 4215 72924 4279 72928
rect 4215 72868 4219 72924
rect 4219 72868 4275 72924
rect 4275 72868 4279 72924
rect 4215 72864 4279 72868
rect 4295 72924 4359 72928
rect 4295 72868 4299 72924
rect 4299 72868 4355 72924
rect 4355 72868 4359 72924
rect 4295 72864 4359 72868
rect 4375 72924 4439 72928
rect 4375 72868 4379 72924
rect 4379 72868 4435 72924
rect 4435 72868 4439 72924
rect 4375 72864 4439 72868
rect 4455 72924 4519 72928
rect 4455 72868 4459 72924
rect 4459 72868 4515 72924
rect 4515 72868 4519 72924
rect 4455 72864 4519 72868
rect 7479 72924 7543 72928
rect 7479 72868 7483 72924
rect 7483 72868 7539 72924
rect 7539 72868 7543 72924
rect 7479 72864 7543 72868
rect 7559 72924 7623 72928
rect 7559 72868 7563 72924
rect 7563 72868 7619 72924
rect 7619 72868 7623 72924
rect 7559 72864 7623 72868
rect 7639 72924 7703 72928
rect 7639 72868 7643 72924
rect 7643 72868 7699 72924
rect 7699 72868 7703 72924
rect 7639 72864 7703 72868
rect 7719 72924 7783 72928
rect 7719 72868 7723 72924
rect 7723 72868 7779 72924
rect 7779 72868 7783 72924
rect 7719 72864 7783 72868
rect 2584 72380 2648 72384
rect 2584 72324 2588 72380
rect 2588 72324 2644 72380
rect 2644 72324 2648 72380
rect 2584 72320 2648 72324
rect 2664 72380 2728 72384
rect 2664 72324 2668 72380
rect 2668 72324 2724 72380
rect 2724 72324 2728 72380
rect 2664 72320 2728 72324
rect 2744 72380 2808 72384
rect 2744 72324 2748 72380
rect 2748 72324 2804 72380
rect 2804 72324 2808 72380
rect 2744 72320 2808 72324
rect 2824 72380 2888 72384
rect 2824 72324 2828 72380
rect 2828 72324 2884 72380
rect 2884 72324 2888 72380
rect 2824 72320 2888 72324
rect 5847 72380 5911 72384
rect 5847 72324 5851 72380
rect 5851 72324 5907 72380
rect 5907 72324 5911 72380
rect 5847 72320 5911 72324
rect 5927 72380 5991 72384
rect 5927 72324 5931 72380
rect 5931 72324 5987 72380
rect 5987 72324 5991 72380
rect 5927 72320 5991 72324
rect 6007 72380 6071 72384
rect 6007 72324 6011 72380
rect 6011 72324 6067 72380
rect 6067 72324 6071 72380
rect 6007 72320 6071 72324
rect 6087 72380 6151 72384
rect 6087 72324 6091 72380
rect 6091 72324 6147 72380
rect 6147 72324 6151 72380
rect 6087 72320 6151 72324
rect 9111 72380 9175 72384
rect 9111 72324 9115 72380
rect 9115 72324 9171 72380
rect 9171 72324 9175 72380
rect 9111 72320 9175 72324
rect 9191 72380 9255 72384
rect 9191 72324 9195 72380
rect 9195 72324 9251 72380
rect 9251 72324 9255 72380
rect 9191 72320 9255 72324
rect 9271 72380 9335 72384
rect 9271 72324 9275 72380
rect 9275 72324 9331 72380
rect 9331 72324 9335 72380
rect 9271 72320 9335 72324
rect 9351 72380 9415 72384
rect 9351 72324 9355 72380
rect 9355 72324 9411 72380
rect 9411 72324 9415 72380
rect 9351 72320 9415 72324
rect 8524 71904 8588 71908
rect 8524 71848 8574 71904
rect 8574 71848 8588 71904
rect 8524 71844 8588 71848
rect 4215 71836 4279 71840
rect 4215 71780 4219 71836
rect 4219 71780 4275 71836
rect 4275 71780 4279 71836
rect 4215 71776 4279 71780
rect 4295 71836 4359 71840
rect 4295 71780 4299 71836
rect 4299 71780 4355 71836
rect 4355 71780 4359 71836
rect 4295 71776 4359 71780
rect 4375 71836 4439 71840
rect 4375 71780 4379 71836
rect 4379 71780 4435 71836
rect 4435 71780 4439 71836
rect 4375 71776 4439 71780
rect 4455 71836 4519 71840
rect 4455 71780 4459 71836
rect 4459 71780 4515 71836
rect 4515 71780 4519 71836
rect 4455 71776 4519 71780
rect 7479 71836 7543 71840
rect 7479 71780 7483 71836
rect 7483 71780 7539 71836
rect 7539 71780 7543 71836
rect 7479 71776 7543 71780
rect 7559 71836 7623 71840
rect 7559 71780 7563 71836
rect 7563 71780 7619 71836
rect 7619 71780 7623 71836
rect 7559 71776 7623 71780
rect 7639 71836 7703 71840
rect 7639 71780 7643 71836
rect 7643 71780 7699 71836
rect 7699 71780 7703 71836
rect 7639 71776 7703 71780
rect 7719 71836 7783 71840
rect 7719 71780 7723 71836
rect 7723 71780 7779 71836
rect 7779 71780 7783 71836
rect 7719 71776 7783 71780
rect 2584 71292 2648 71296
rect 2584 71236 2588 71292
rect 2588 71236 2644 71292
rect 2644 71236 2648 71292
rect 2584 71232 2648 71236
rect 2664 71292 2728 71296
rect 2664 71236 2668 71292
rect 2668 71236 2724 71292
rect 2724 71236 2728 71292
rect 2664 71232 2728 71236
rect 2744 71292 2808 71296
rect 2744 71236 2748 71292
rect 2748 71236 2804 71292
rect 2804 71236 2808 71292
rect 2744 71232 2808 71236
rect 2824 71292 2888 71296
rect 2824 71236 2828 71292
rect 2828 71236 2884 71292
rect 2884 71236 2888 71292
rect 2824 71232 2888 71236
rect 5847 71292 5911 71296
rect 5847 71236 5851 71292
rect 5851 71236 5907 71292
rect 5907 71236 5911 71292
rect 5847 71232 5911 71236
rect 5927 71292 5991 71296
rect 5927 71236 5931 71292
rect 5931 71236 5987 71292
rect 5987 71236 5991 71292
rect 5927 71232 5991 71236
rect 6007 71292 6071 71296
rect 6007 71236 6011 71292
rect 6011 71236 6067 71292
rect 6067 71236 6071 71292
rect 6007 71232 6071 71236
rect 6087 71292 6151 71296
rect 6087 71236 6091 71292
rect 6091 71236 6147 71292
rect 6147 71236 6151 71292
rect 6087 71232 6151 71236
rect 9111 71292 9175 71296
rect 9111 71236 9115 71292
rect 9115 71236 9171 71292
rect 9171 71236 9175 71292
rect 9111 71232 9175 71236
rect 9191 71292 9255 71296
rect 9191 71236 9195 71292
rect 9195 71236 9251 71292
rect 9251 71236 9255 71292
rect 9191 71232 9255 71236
rect 9271 71292 9335 71296
rect 9271 71236 9275 71292
rect 9275 71236 9331 71292
rect 9331 71236 9335 71292
rect 9271 71232 9335 71236
rect 9351 71292 9415 71296
rect 9351 71236 9355 71292
rect 9355 71236 9411 71292
rect 9411 71236 9415 71292
rect 9351 71232 9415 71236
rect 4215 70748 4279 70752
rect 4215 70692 4219 70748
rect 4219 70692 4275 70748
rect 4275 70692 4279 70748
rect 4215 70688 4279 70692
rect 4295 70748 4359 70752
rect 4295 70692 4299 70748
rect 4299 70692 4355 70748
rect 4355 70692 4359 70748
rect 4295 70688 4359 70692
rect 4375 70748 4439 70752
rect 4375 70692 4379 70748
rect 4379 70692 4435 70748
rect 4435 70692 4439 70748
rect 4375 70688 4439 70692
rect 4455 70748 4519 70752
rect 4455 70692 4459 70748
rect 4459 70692 4515 70748
rect 4515 70692 4519 70748
rect 4455 70688 4519 70692
rect 7479 70748 7543 70752
rect 7479 70692 7483 70748
rect 7483 70692 7539 70748
rect 7539 70692 7543 70748
rect 7479 70688 7543 70692
rect 7559 70748 7623 70752
rect 7559 70692 7563 70748
rect 7563 70692 7619 70748
rect 7619 70692 7623 70748
rect 7559 70688 7623 70692
rect 7639 70748 7703 70752
rect 7639 70692 7643 70748
rect 7643 70692 7699 70748
rect 7699 70692 7703 70748
rect 7639 70688 7703 70692
rect 7719 70748 7783 70752
rect 7719 70692 7723 70748
rect 7723 70692 7779 70748
rect 7779 70692 7783 70748
rect 7719 70688 7783 70692
rect 2584 70204 2648 70208
rect 2584 70148 2588 70204
rect 2588 70148 2644 70204
rect 2644 70148 2648 70204
rect 2584 70144 2648 70148
rect 2664 70204 2728 70208
rect 2664 70148 2668 70204
rect 2668 70148 2724 70204
rect 2724 70148 2728 70204
rect 2664 70144 2728 70148
rect 2744 70204 2808 70208
rect 2744 70148 2748 70204
rect 2748 70148 2804 70204
rect 2804 70148 2808 70204
rect 2744 70144 2808 70148
rect 2824 70204 2888 70208
rect 2824 70148 2828 70204
rect 2828 70148 2884 70204
rect 2884 70148 2888 70204
rect 2824 70144 2888 70148
rect 5847 70204 5911 70208
rect 5847 70148 5851 70204
rect 5851 70148 5907 70204
rect 5907 70148 5911 70204
rect 5847 70144 5911 70148
rect 5927 70204 5991 70208
rect 5927 70148 5931 70204
rect 5931 70148 5987 70204
rect 5987 70148 5991 70204
rect 5927 70144 5991 70148
rect 6007 70204 6071 70208
rect 6007 70148 6011 70204
rect 6011 70148 6067 70204
rect 6067 70148 6071 70204
rect 6007 70144 6071 70148
rect 6087 70204 6151 70208
rect 6087 70148 6091 70204
rect 6091 70148 6147 70204
rect 6147 70148 6151 70204
rect 6087 70144 6151 70148
rect 9111 70204 9175 70208
rect 9111 70148 9115 70204
rect 9115 70148 9171 70204
rect 9171 70148 9175 70204
rect 9111 70144 9175 70148
rect 9191 70204 9255 70208
rect 9191 70148 9195 70204
rect 9195 70148 9251 70204
rect 9251 70148 9255 70204
rect 9191 70144 9255 70148
rect 9271 70204 9335 70208
rect 9271 70148 9275 70204
rect 9275 70148 9331 70204
rect 9331 70148 9335 70204
rect 9271 70144 9335 70148
rect 9351 70204 9415 70208
rect 9351 70148 9355 70204
rect 9355 70148 9411 70204
rect 9411 70148 9415 70204
rect 9351 70144 9415 70148
rect 4215 69660 4279 69664
rect 4215 69604 4219 69660
rect 4219 69604 4275 69660
rect 4275 69604 4279 69660
rect 4215 69600 4279 69604
rect 4295 69660 4359 69664
rect 4295 69604 4299 69660
rect 4299 69604 4355 69660
rect 4355 69604 4359 69660
rect 4295 69600 4359 69604
rect 4375 69660 4439 69664
rect 4375 69604 4379 69660
rect 4379 69604 4435 69660
rect 4435 69604 4439 69660
rect 4375 69600 4439 69604
rect 4455 69660 4519 69664
rect 4455 69604 4459 69660
rect 4459 69604 4515 69660
rect 4515 69604 4519 69660
rect 4455 69600 4519 69604
rect 7479 69660 7543 69664
rect 7479 69604 7483 69660
rect 7483 69604 7539 69660
rect 7539 69604 7543 69660
rect 7479 69600 7543 69604
rect 7559 69660 7623 69664
rect 7559 69604 7563 69660
rect 7563 69604 7619 69660
rect 7619 69604 7623 69660
rect 7559 69600 7623 69604
rect 7639 69660 7703 69664
rect 7639 69604 7643 69660
rect 7643 69604 7699 69660
rect 7699 69604 7703 69660
rect 7639 69600 7703 69604
rect 7719 69660 7783 69664
rect 7719 69604 7723 69660
rect 7723 69604 7779 69660
rect 7779 69604 7783 69660
rect 7719 69600 7783 69604
rect 8892 69260 8956 69324
rect 2584 69116 2648 69120
rect 2584 69060 2588 69116
rect 2588 69060 2644 69116
rect 2644 69060 2648 69116
rect 2584 69056 2648 69060
rect 2664 69116 2728 69120
rect 2664 69060 2668 69116
rect 2668 69060 2724 69116
rect 2724 69060 2728 69116
rect 2664 69056 2728 69060
rect 2744 69116 2808 69120
rect 2744 69060 2748 69116
rect 2748 69060 2804 69116
rect 2804 69060 2808 69116
rect 2744 69056 2808 69060
rect 2824 69116 2888 69120
rect 2824 69060 2828 69116
rect 2828 69060 2884 69116
rect 2884 69060 2888 69116
rect 2824 69056 2888 69060
rect 5847 69116 5911 69120
rect 5847 69060 5851 69116
rect 5851 69060 5907 69116
rect 5907 69060 5911 69116
rect 5847 69056 5911 69060
rect 5927 69116 5991 69120
rect 5927 69060 5931 69116
rect 5931 69060 5987 69116
rect 5987 69060 5991 69116
rect 5927 69056 5991 69060
rect 6007 69116 6071 69120
rect 6007 69060 6011 69116
rect 6011 69060 6067 69116
rect 6067 69060 6071 69116
rect 6007 69056 6071 69060
rect 6087 69116 6151 69120
rect 6087 69060 6091 69116
rect 6091 69060 6147 69116
rect 6147 69060 6151 69116
rect 6087 69056 6151 69060
rect 9111 69116 9175 69120
rect 9111 69060 9115 69116
rect 9115 69060 9171 69116
rect 9171 69060 9175 69116
rect 9111 69056 9175 69060
rect 9191 69116 9255 69120
rect 9191 69060 9195 69116
rect 9195 69060 9251 69116
rect 9251 69060 9255 69116
rect 9191 69056 9255 69060
rect 9271 69116 9335 69120
rect 9271 69060 9275 69116
rect 9275 69060 9331 69116
rect 9331 69060 9335 69116
rect 9271 69056 9335 69060
rect 9351 69116 9415 69120
rect 9351 69060 9355 69116
rect 9355 69060 9411 69116
rect 9411 69060 9415 69116
rect 9351 69056 9415 69060
rect 4215 68572 4279 68576
rect 4215 68516 4219 68572
rect 4219 68516 4275 68572
rect 4275 68516 4279 68572
rect 4215 68512 4279 68516
rect 4295 68572 4359 68576
rect 4295 68516 4299 68572
rect 4299 68516 4355 68572
rect 4355 68516 4359 68572
rect 4295 68512 4359 68516
rect 4375 68572 4439 68576
rect 4375 68516 4379 68572
rect 4379 68516 4435 68572
rect 4435 68516 4439 68572
rect 4375 68512 4439 68516
rect 4455 68572 4519 68576
rect 4455 68516 4459 68572
rect 4459 68516 4515 68572
rect 4515 68516 4519 68572
rect 4455 68512 4519 68516
rect 7479 68572 7543 68576
rect 7479 68516 7483 68572
rect 7483 68516 7539 68572
rect 7539 68516 7543 68572
rect 7479 68512 7543 68516
rect 7559 68572 7623 68576
rect 7559 68516 7563 68572
rect 7563 68516 7619 68572
rect 7619 68516 7623 68572
rect 7559 68512 7623 68516
rect 7639 68572 7703 68576
rect 7639 68516 7643 68572
rect 7643 68516 7699 68572
rect 7699 68516 7703 68572
rect 7639 68512 7703 68516
rect 7719 68572 7783 68576
rect 7719 68516 7723 68572
rect 7723 68516 7779 68572
rect 7779 68516 7783 68572
rect 7719 68512 7783 68516
rect 2584 68028 2648 68032
rect 2584 67972 2588 68028
rect 2588 67972 2644 68028
rect 2644 67972 2648 68028
rect 2584 67968 2648 67972
rect 2664 68028 2728 68032
rect 2664 67972 2668 68028
rect 2668 67972 2724 68028
rect 2724 67972 2728 68028
rect 2664 67968 2728 67972
rect 2744 68028 2808 68032
rect 2744 67972 2748 68028
rect 2748 67972 2804 68028
rect 2804 67972 2808 68028
rect 2744 67968 2808 67972
rect 2824 68028 2888 68032
rect 2824 67972 2828 68028
rect 2828 67972 2884 68028
rect 2884 67972 2888 68028
rect 2824 67968 2888 67972
rect 5847 68028 5911 68032
rect 5847 67972 5851 68028
rect 5851 67972 5907 68028
rect 5907 67972 5911 68028
rect 5847 67968 5911 67972
rect 5927 68028 5991 68032
rect 5927 67972 5931 68028
rect 5931 67972 5987 68028
rect 5987 67972 5991 68028
rect 5927 67968 5991 67972
rect 6007 68028 6071 68032
rect 6007 67972 6011 68028
rect 6011 67972 6067 68028
rect 6067 67972 6071 68028
rect 6007 67968 6071 67972
rect 6087 68028 6151 68032
rect 6087 67972 6091 68028
rect 6091 67972 6147 68028
rect 6147 67972 6151 68028
rect 6087 67968 6151 67972
rect 9111 68028 9175 68032
rect 9111 67972 9115 68028
rect 9115 67972 9171 68028
rect 9171 67972 9175 68028
rect 9111 67968 9175 67972
rect 9191 68028 9255 68032
rect 9191 67972 9195 68028
rect 9195 67972 9251 68028
rect 9251 67972 9255 68028
rect 9191 67968 9255 67972
rect 9271 68028 9335 68032
rect 9271 67972 9275 68028
rect 9275 67972 9331 68028
rect 9331 67972 9335 68028
rect 9271 67968 9335 67972
rect 9351 68028 9415 68032
rect 9351 67972 9355 68028
rect 9355 67972 9411 68028
rect 9411 67972 9415 68028
rect 9351 67968 9415 67972
rect 8708 67628 8772 67692
rect 4215 67484 4279 67488
rect 4215 67428 4219 67484
rect 4219 67428 4275 67484
rect 4275 67428 4279 67484
rect 4215 67424 4279 67428
rect 4295 67484 4359 67488
rect 4295 67428 4299 67484
rect 4299 67428 4355 67484
rect 4355 67428 4359 67484
rect 4295 67424 4359 67428
rect 4375 67484 4439 67488
rect 4375 67428 4379 67484
rect 4379 67428 4435 67484
rect 4435 67428 4439 67484
rect 4375 67424 4439 67428
rect 4455 67484 4519 67488
rect 4455 67428 4459 67484
rect 4459 67428 4515 67484
rect 4515 67428 4519 67484
rect 4455 67424 4519 67428
rect 7479 67484 7543 67488
rect 7479 67428 7483 67484
rect 7483 67428 7539 67484
rect 7539 67428 7543 67484
rect 7479 67424 7543 67428
rect 7559 67484 7623 67488
rect 7559 67428 7563 67484
rect 7563 67428 7619 67484
rect 7619 67428 7623 67484
rect 7559 67424 7623 67428
rect 7639 67484 7703 67488
rect 7639 67428 7643 67484
rect 7643 67428 7699 67484
rect 7699 67428 7703 67484
rect 7639 67424 7703 67428
rect 7719 67484 7783 67488
rect 7719 67428 7723 67484
rect 7723 67428 7779 67484
rect 7779 67428 7783 67484
rect 7719 67424 7783 67428
rect 2584 66940 2648 66944
rect 2584 66884 2588 66940
rect 2588 66884 2644 66940
rect 2644 66884 2648 66940
rect 2584 66880 2648 66884
rect 2664 66940 2728 66944
rect 2664 66884 2668 66940
rect 2668 66884 2724 66940
rect 2724 66884 2728 66940
rect 2664 66880 2728 66884
rect 2744 66940 2808 66944
rect 2744 66884 2748 66940
rect 2748 66884 2804 66940
rect 2804 66884 2808 66940
rect 2744 66880 2808 66884
rect 2824 66940 2888 66944
rect 2824 66884 2828 66940
rect 2828 66884 2884 66940
rect 2884 66884 2888 66940
rect 2824 66880 2888 66884
rect 5847 66940 5911 66944
rect 5847 66884 5851 66940
rect 5851 66884 5907 66940
rect 5907 66884 5911 66940
rect 5847 66880 5911 66884
rect 5927 66940 5991 66944
rect 5927 66884 5931 66940
rect 5931 66884 5987 66940
rect 5987 66884 5991 66940
rect 5927 66880 5991 66884
rect 6007 66940 6071 66944
rect 6007 66884 6011 66940
rect 6011 66884 6067 66940
rect 6067 66884 6071 66940
rect 6007 66880 6071 66884
rect 6087 66940 6151 66944
rect 6087 66884 6091 66940
rect 6091 66884 6147 66940
rect 6147 66884 6151 66940
rect 6087 66880 6151 66884
rect 9111 66940 9175 66944
rect 9111 66884 9115 66940
rect 9115 66884 9171 66940
rect 9171 66884 9175 66940
rect 9111 66880 9175 66884
rect 9191 66940 9255 66944
rect 9191 66884 9195 66940
rect 9195 66884 9251 66940
rect 9251 66884 9255 66940
rect 9191 66880 9255 66884
rect 9271 66940 9335 66944
rect 9271 66884 9275 66940
rect 9275 66884 9331 66940
rect 9331 66884 9335 66940
rect 9271 66880 9335 66884
rect 9351 66940 9415 66944
rect 9351 66884 9355 66940
rect 9355 66884 9411 66940
rect 9411 66884 9415 66940
rect 9351 66880 9415 66884
rect 9628 66540 9692 66604
rect 4215 66396 4279 66400
rect 4215 66340 4219 66396
rect 4219 66340 4275 66396
rect 4275 66340 4279 66396
rect 4215 66336 4279 66340
rect 4295 66396 4359 66400
rect 4295 66340 4299 66396
rect 4299 66340 4355 66396
rect 4355 66340 4359 66396
rect 4295 66336 4359 66340
rect 4375 66396 4439 66400
rect 4375 66340 4379 66396
rect 4379 66340 4435 66396
rect 4435 66340 4439 66396
rect 4375 66336 4439 66340
rect 4455 66396 4519 66400
rect 4455 66340 4459 66396
rect 4459 66340 4515 66396
rect 4515 66340 4519 66396
rect 4455 66336 4519 66340
rect 7479 66396 7543 66400
rect 7479 66340 7483 66396
rect 7483 66340 7539 66396
rect 7539 66340 7543 66396
rect 7479 66336 7543 66340
rect 7559 66396 7623 66400
rect 7559 66340 7563 66396
rect 7563 66340 7619 66396
rect 7619 66340 7623 66396
rect 7559 66336 7623 66340
rect 7639 66396 7703 66400
rect 7639 66340 7643 66396
rect 7643 66340 7699 66396
rect 7699 66340 7703 66396
rect 7639 66336 7703 66340
rect 7719 66396 7783 66400
rect 7719 66340 7723 66396
rect 7723 66340 7779 66396
rect 7779 66340 7783 66396
rect 7719 66336 7783 66340
rect 8340 66328 8404 66332
rect 8340 66272 8354 66328
rect 8354 66272 8404 66328
rect 8340 66268 8404 66272
rect 2584 65852 2648 65856
rect 2584 65796 2588 65852
rect 2588 65796 2644 65852
rect 2644 65796 2648 65852
rect 2584 65792 2648 65796
rect 2664 65852 2728 65856
rect 2664 65796 2668 65852
rect 2668 65796 2724 65852
rect 2724 65796 2728 65852
rect 2664 65792 2728 65796
rect 2744 65852 2808 65856
rect 2744 65796 2748 65852
rect 2748 65796 2804 65852
rect 2804 65796 2808 65852
rect 2744 65792 2808 65796
rect 2824 65852 2888 65856
rect 2824 65796 2828 65852
rect 2828 65796 2884 65852
rect 2884 65796 2888 65852
rect 2824 65792 2888 65796
rect 5847 65852 5911 65856
rect 5847 65796 5851 65852
rect 5851 65796 5907 65852
rect 5907 65796 5911 65852
rect 5847 65792 5911 65796
rect 5927 65852 5991 65856
rect 5927 65796 5931 65852
rect 5931 65796 5987 65852
rect 5987 65796 5991 65852
rect 5927 65792 5991 65796
rect 6007 65852 6071 65856
rect 6007 65796 6011 65852
rect 6011 65796 6067 65852
rect 6067 65796 6071 65852
rect 6007 65792 6071 65796
rect 6087 65852 6151 65856
rect 6087 65796 6091 65852
rect 6091 65796 6147 65852
rect 6147 65796 6151 65852
rect 6087 65792 6151 65796
rect 9111 65852 9175 65856
rect 9111 65796 9115 65852
rect 9115 65796 9171 65852
rect 9171 65796 9175 65852
rect 9111 65792 9175 65796
rect 9191 65852 9255 65856
rect 9191 65796 9195 65852
rect 9195 65796 9251 65852
rect 9251 65796 9255 65852
rect 9191 65792 9255 65796
rect 9271 65852 9335 65856
rect 9271 65796 9275 65852
rect 9275 65796 9331 65852
rect 9331 65796 9335 65852
rect 9271 65792 9335 65796
rect 9351 65852 9415 65856
rect 9351 65796 9355 65852
rect 9355 65796 9411 65852
rect 9411 65796 9415 65852
rect 9351 65792 9415 65796
rect 4215 65308 4279 65312
rect 4215 65252 4219 65308
rect 4219 65252 4275 65308
rect 4275 65252 4279 65308
rect 4215 65248 4279 65252
rect 4295 65308 4359 65312
rect 4295 65252 4299 65308
rect 4299 65252 4355 65308
rect 4355 65252 4359 65308
rect 4295 65248 4359 65252
rect 4375 65308 4439 65312
rect 4375 65252 4379 65308
rect 4379 65252 4435 65308
rect 4435 65252 4439 65308
rect 4375 65248 4439 65252
rect 4455 65308 4519 65312
rect 4455 65252 4459 65308
rect 4459 65252 4515 65308
rect 4515 65252 4519 65308
rect 4455 65248 4519 65252
rect 7479 65308 7543 65312
rect 7479 65252 7483 65308
rect 7483 65252 7539 65308
rect 7539 65252 7543 65308
rect 7479 65248 7543 65252
rect 7559 65308 7623 65312
rect 7559 65252 7563 65308
rect 7563 65252 7619 65308
rect 7619 65252 7623 65308
rect 7559 65248 7623 65252
rect 7639 65308 7703 65312
rect 7639 65252 7643 65308
rect 7643 65252 7699 65308
rect 7699 65252 7703 65308
rect 7639 65248 7703 65252
rect 7719 65308 7783 65312
rect 7719 65252 7723 65308
rect 7723 65252 7779 65308
rect 7779 65252 7783 65308
rect 7719 65248 7783 65252
rect 2584 64764 2648 64768
rect 2584 64708 2588 64764
rect 2588 64708 2644 64764
rect 2644 64708 2648 64764
rect 2584 64704 2648 64708
rect 2664 64764 2728 64768
rect 2664 64708 2668 64764
rect 2668 64708 2724 64764
rect 2724 64708 2728 64764
rect 2664 64704 2728 64708
rect 2744 64764 2808 64768
rect 2744 64708 2748 64764
rect 2748 64708 2804 64764
rect 2804 64708 2808 64764
rect 2744 64704 2808 64708
rect 2824 64764 2888 64768
rect 2824 64708 2828 64764
rect 2828 64708 2884 64764
rect 2884 64708 2888 64764
rect 2824 64704 2888 64708
rect 5847 64764 5911 64768
rect 5847 64708 5851 64764
rect 5851 64708 5907 64764
rect 5907 64708 5911 64764
rect 5847 64704 5911 64708
rect 5927 64764 5991 64768
rect 5927 64708 5931 64764
rect 5931 64708 5987 64764
rect 5987 64708 5991 64764
rect 5927 64704 5991 64708
rect 6007 64764 6071 64768
rect 6007 64708 6011 64764
rect 6011 64708 6067 64764
rect 6067 64708 6071 64764
rect 6007 64704 6071 64708
rect 6087 64764 6151 64768
rect 6087 64708 6091 64764
rect 6091 64708 6147 64764
rect 6147 64708 6151 64764
rect 6087 64704 6151 64708
rect 9111 64764 9175 64768
rect 9111 64708 9115 64764
rect 9115 64708 9171 64764
rect 9171 64708 9175 64764
rect 9111 64704 9175 64708
rect 9191 64764 9255 64768
rect 9191 64708 9195 64764
rect 9195 64708 9251 64764
rect 9251 64708 9255 64764
rect 9191 64704 9255 64708
rect 9271 64764 9335 64768
rect 9271 64708 9275 64764
rect 9275 64708 9331 64764
rect 9331 64708 9335 64764
rect 9271 64704 9335 64708
rect 9351 64764 9415 64768
rect 9351 64708 9355 64764
rect 9355 64708 9411 64764
rect 9411 64708 9415 64764
rect 9351 64704 9415 64708
rect 4215 64220 4279 64224
rect 4215 64164 4219 64220
rect 4219 64164 4275 64220
rect 4275 64164 4279 64220
rect 4215 64160 4279 64164
rect 4295 64220 4359 64224
rect 4295 64164 4299 64220
rect 4299 64164 4355 64220
rect 4355 64164 4359 64220
rect 4295 64160 4359 64164
rect 4375 64220 4439 64224
rect 4375 64164 4379 64220
rect 4379 64164 4435 64220
rect 4435 64164 4439 64220
rect 4375 64160 4439 64164
rect 4455 64220 4519 64224
rect 4455 64164 4459 64220
rect 4459 64164 4515 64220
rect 4515 64164 4519 64220
rect 4455 64160 4519 64164
rect 7479 64220 7543 64224
rect 7479 64164 7483 64220
rect 7483 64164 7539 64220
rect 7539 64164 7543 64220
rect 7479 64160 7543 64164
rect 7559 64220 7623 64224
rect 7559 64164 7563 64220
rect 7563 64164 7619 64220
rect 7619 64164 7623 64220
rect 7559 64160 7623 64164
rect 7639 64220 7703 64224
rect 7639 64164 7643 64220
rect 7643 64164 7699 64220
rect 7699 64164 7703 64220
rect 7639 64160 7703 64164
rect 7719 64220 7783 64224
rect 7719 64164 7723 64220
rect 7723 64164 7779 64220
rect 7779 64164 7783 64220
rect 7719 64160 7783 64164
rect 2584 63676 2648 63680
rect 2584 63620 2588 63676
rect 2588 63620 2644 63676
rect 2644 63620 2648 63676
rect 2584 63616 2648 63620
rect 2664 63676 2728 63680
rect 2664 63620 2668 63676
rect 2668 63620 2724 63676
rect 2724 63620 2728 63676
rect 2664 63616 2728 63620
rect 2744 63676 2808 63680
rect 2744 63620 2748 63676
rect 2748 63620 2804 63676
rect 2804 63620 2808 63676
rect 2744 63616 2808 63620
rect 2824 63676 2888 63680
rect 2824 63620 2828 63676
rect 2828 63620 2884 63676
rect 2884 63620 2888 63676
rect 2824 63616 2888 63620
rect 5847 63676 5911 63680
rect 5847 63620 5851 63676
rect 5851 63620 5907 63676
rect 5907 63620 5911 63676
rect 5847 63616 5911 63620
rect 5927 63676 5991 63680
rect 5927 63620 5931 63676
rect 5931 63620 5987 63676
rect 5987 63620 5991 63676
rect 5927 63616 5991 63620
rect 6007 63676 6071 63680
rect 6007 63620 6011 63676
rect 6011 63620 6067 63676
rect 6067 63620 6071 63676
rect 6007 63616 6071 63620
rect 6087 63676 6151 63680
rect 6087 63620 6091 63676
rect 6091 63620 6147 63676
rect 6147 63620 6151 63676
rect 6087 63616 6151 63620
rect 9111 63676 9175 63680
rect 9111 63620 9115 63676
rect 9115 63620 9171 63676
rect 9171 63620 9175 63676
rect 9111 63616 9175 63620
rect 9191 63676 9255 63680
rect 9191 63620 9195 63676
rect 9195 63620 9251 63676
rect 9251 63620 9255 63676
rect 9191 63616 9255 63620
rect 9271 63676 9335 63680
rect 9271 63620 9275 63676
rect 9275 63620 9331 63676
rect 9331 63620 9335 63676
rect 9271 63616 9335 63620
rect 9351 63676 9415 63680
rect 9351 63620 9355 63676
rect 9355 63620 9411 63676
rect 9411 63620 9415 63676
rect 9351 63616 9415 63620
rect 4215 63132 4279 63136
rect 4215 63076 4219 63132
rect 4219 63076 4275 63132
rect 4275 63076 4279 63132
rect 4215 63072 4279 63076
rect 4295 63132 4359 63136
rect 4295 63076 4299 63132
rect 4299 63076 4355 63132
rect 4355 63076 4359 63132
rect 4295 63072 4359 63076
rect 4375 63132 4439 63136
rect 4375 63076 4379 63132
rect 4379 63076 4435 63132
rect 4435 63076 4439 63132
rect 4375 63072 4439 63076
rect 4455 63132 4519 63136
rect 4455 63076 4459 63132
rect 4459 63076 4515 63132
rect 4515 63076 4519 63132
rect 4455 63072 4519 63076
rect 7479 63132 7543 63136
rect 7479 63076 7483 63132
rect 7483 63076 7539 63132
rect 7539 63076 7543 63132
rect 7479 63072 7543 63076
rect 7559 63132 7623 63136
rect 7559 63076 7563 63132
rect 7563 63076 7619 63132
rect 7619 63076 7623 63132
rect 7559 63072 7623 63076
rect 7639 63132 7703 63136
rect 7639 63076 7643 63132
rect 7643 63076 7699 63132
rect 7699 63076 7703 63132
rect 7639 63072 7703 63076
rect 7719 63132 7783 63136
rect 7719 63076 7723 63132
rect 7723 63076 7779 63132
rect 7779 63076 7783 63132
rect 7719 63072 7783 63076
rect 3556 62732 3620 62796
rect 2584 62588 2648 62592
rect 2584 62532 2588 62588
rect 2588 62532 2644 62588
rect 2644 62532 2648 62588
rect 2584 62528 2648 62532
rect 2664 62588 2728 62592
rect 2664 62532 2668 62588
rect 2668 62532 2724 62588
rect 2724 62532 2728 62588
rect 2664 62528 2728 62532
rect 2744 62588 2808 62592
rect 2744 62532 2748 62588
rect 2748 62532 2804 62588
rect 2804 62532 2808 62588
rect 2744 62528 2808 62532
rect 2824 62588 2888 62592
rect 2824 62532 2828 62588
rect 2828 62532 2884 62588
rect 2884 62532 2888 62588
rect 2824 62528 2888 62532
rect 5847 62588 5911 62592
rect 5847 62532 5851 62588
rect 5851 62532 5907 62588
rect 5907 62532 5911 62588
rect 5847 62528 5911 62532
rect 5927 62588 5991 62592
rect 5927 62532 5931 62588
rect 5931 62532 5987 62588
rect 5987 62532 5991 62588
rect 5927 62528 5991 62532
rect 6007 62588 6071 62592
rect 6007 62532 6011 62588
rect 6011 62532 6067 62588
rect 6067 62532 6071 62588
rect 6007 62528 6071 62532
rect 6087 62588 6151 62592
rect 6087 62532 6091 62588
rect 6091 62532 6147 62588
rect 6147 62532 6151 62588
rect 6087 62528 6151 62532
rect 9111 62588 9175 62592
rect 9111 62532 9115 62588
rect 9115 62532 9171 62588
rect 9171 62532 9175 62588
rect 9111 62528 9175 62532
rect 9191 62588 9255 62592
rect 9191 62532 9195 62588
rect 9195 62532 9251 62588
rect 9251 62532 9255 62588
rect 9191 62528 9255 62532
rect 9271 62588 9335 62592
rect 9271 62532 9275 62588
rect 9275 62532 9331 62588
rect 9331 62532 9335 62588
rect 9271 62528 9335 62532
rect 9351 62588 9415 62592
rect 9351 62532 9355 62588
rect 9355 62532 9411 62588
rect 9411 62532 9415 62588
rect 9351 62528 9415 62532
rect 4215 62044 4279 62048
rect 4215 61988 4219 62044
rect 4219 61988 4275 62044
rect 4275 61988 4279 62044
rect 4215 61984 4279 61988
rect 4295 62044 4359 62048
rect 4295 61988 4299 62044
rect 4299 61988 4355 62044
rect 4355 61988 4359 62044
rect 4295 61984 4359 61988
rect 4375 62044 4439 62048
rect 4375 61988 4379 62044
rect 4379 61988 4435 62044
rect 4435 61988 4439 62044
rect 4375 61984 4439 61988
rect 4455 62044 4519 62048
rect 4455 61988 4459 62044
rect 4459 61988 4515 62044
rect 4515 61988 4519 62044
rect 4455 61984 4519 61988
rect 7479 62044 7543 62048
rect 7479 61988 7483 62044
rect 7483 61988 7539 62044
rect 7539 61988 7543 62044
rect 7479 61984 7543 61988
rect 7559 62044 7623 62048
rect 7559 61988 7563 62044
rect 7563 61988 7619 62044
rect 7619 61988 7623 62044
rect 7559 61984 7623 61988
rect 7639 62044 7703 62048
rect 7639 61988 7643 62044
rect 7643 61988 7699 62044
rect 7699 61988 7703 62044
rect 7639 61984 7703 61988
rect 7719 62044 7783 62048
rect 7719 61988 7723 62044
rect 7723 61988 7779 62044
rect 7779 61988 7783 62044
rect 7719 61984 7783 61988
rect 2584 61500 2648 61504
rect 2584 61444 2588 61500
rect 2588 61444 2644 61500
rect 2644 61444 2648 61500
rect 2584 61440 2648 61444
rect 2664 61500 2728 61504
rect 2664 61444 2668 61500
rect 2668 61444 2724 61500
rect 2724 61444 2728 61500
rect 2664 61440 2728 61444
rect 2744 61500 2808 61504
rect 2744 61444 2748 61500
rect 2748 61444 2804 61500
rect 2804 61444 2808 61500
rect 2744 61440 2808 61444
rect 2824 61500 2888 61504
rect 2824 61444 2828 61500
rect 2828 61444 2884 61500
rect 2884 61444 2888 61500
rect 2824 61440 2888 61444
rect 5847 61500 5911 61504
rect 5847 61444 5851 61500
rect 5851 61444 5907 61500
rect 5907 61444 5911 61500
rect 5847 61440 5911 61444
rect 5927 61500 5991 61504
rect 5927 61444 5931 61500
rect 5931 61444 5987 61500
rect 5987 61444 5991 61500
rect 5927 61440 5991 61444
rect 6007 61500 6071 61504
rect 6007 61444 6011 61500
rect 6011 61444 6067 61500
rect 6067 61444 6071 61500
rect 6007 61440 6071 61444
rect 6087 61500 6151 61504
rect 6087 61444 6091 61500
rect 6091 61444 6147 61500
rect 6147 61444 6151 61500
rect 6087 61440 6151 61444
rect 9111 61500 9175 61504
rect 9111 61444 9115 61500
rect 9115 61444 9171 61500
rect 9171 61444 9175 61500
rect 9111 61440 9175 61444
rect 9191 61500 9255 61504
rect 9191 61444 9195 61500
rect 9195 61444 9251 61500
rect 9251 61444 9255 61500
rect 9191 61440 9255 61444
rect 9271 61500 9335 61504
rect 9271 61444 9275 61500
rect 9275 61444 9331 61500
rect 9331 61444 9335 61500
rect 9271 61440 9335 61444
rect 9351 61500 9415 61504
rect 9351 61444 9355 61500
rect 9355 61444 9411 61500
rect 9411 61444 9415 61500
rect 9351 61440 9415 61444
rect 8156 61236 8220 61300
rect 9628 61236 9692 61300
rect 4215 60956 4279 60960
rect 4215 60900 4219 60956
rect 4219 60900 4275 60956
rect 4275 60900 4279 60956
rect 4215 60896 4279 60900
rect 4295 60956 4359 60960
rect 4295 60900 4299 60956
rect 4299 60900 4355 60956
rect 4355 60900 4359 60956
rect 4295 60896 4359 60900
rect 4375 60956 4439 60960
rect 4375 60900 4379 60956
rect 4379 60900 4435 60956
rect 4435 60900 4439 60956
rect 4375 60896 4439 60900
rect 4455 60956 4519 60960
rect 4455 60900 4459 60956
rect 4459 60900 4515 60956
rect 4515 60900 4519 60956
rect 4455 60896 4519 60900
rect 7479 60956 7543 60960
rect 7479 60900 7483 60956
rect 7483 60900 7539 60956
rect 7539 60900 7543 60956
rect 7479 60896 7543 60900
rect 7559 60956 7623 60960
rect 7559 60900 7563 60956
rect 7563 60900 7619 60956
rect 7619 60900 7623 60956
rect 7559 60896 7623 60900
rect 7639 60956 7703 60960
rect 7639 60900 7643 60956
rect 7643 60900 7699 60956
rect 7699 60900 7703 60956
rect 7639 60896 7703 60900
rect 7719 60956 7783 60960
rect 7719 60900 7723 60956
rect 7723 60900 7779 60956
rect 7779 60900 7783 60956
rect 7719 60896 7783 60900
rect 8156 60556 8220 60620
rect 9628 60556 9692 60620
rect 10180 60616 10244 60620
rect 10180 60560 10230 60616
rect 10230 60560 10244 60616
rect 10180 60556 10244 60560
rect 2584 60412 2648 60416
rect 2584 60356 2588 60412
rect 2588 60356 2644 60412
rect 2644 60356 2648 60412
rect 2584 60352 2648 60356
rect 2664 60412 2728 60416
rect 2664 60356 2668 60412
rect 2668 60356 2724 60412
rect 2724 60356 2728 60412
rect 2664 60352 2728 60356
rect 2744 60412 2808 60416
rect 2744 60356 2748 60412
rect 2748 60356 2804 60412
rect 2804 60356 2808 60412
rect 2744 60352 2808 60356
rect 2824 60412 2888 60416
rect 2824 60356 2828 60412
rect 2828 60356 2884 60412
rect 2884 60356 2888 60412
rect 2824 60352 2888 60356
rect 5847 60412 5911 60416
rect 5847 60356 5851 60412
rect 5851 60356 5907 60412
rect 5907 60356 5911 60412
rect 5847 60352 5911 60356
rect 5927 60412 5991 60416
rect 5927 60356 5931 60412
rect 5931 60356 5987 60412
rect 5987 60356 5991 60412
rect 5927 60352 5991 60356
rect 6007 60412 6071 60416
rect 6007 60356 6011 60412
rect 6011 60356 6067 60412
rect 6067 60356 6071 60412
rect 6007 60352 6071 60356
rect 6087 60412 6151 60416
rect 6087 60356 6091 60412
rect 6091 60356 6147 60412
rect 6147 60356 6151 60412
rect 6087 60352 6151 60356
rect 9111 60412 9175 60416
rect 9111 60356 9115 60412
rect 9115 60356 9171 60412
rect 9171 60356 9175 60412
rect 9111 60352 9175 60356
rect 9191 60412 9255 60416
rect 9191 60356 9195 60412
rect 9195 60356 9251 60412
rect 9251 60356 9255 60412
rect 9191 60352 9255 60356
rect 9271 60412 9335 60416
rect 9271 60356 9275 60412
rect 9275 60356 9331 60412
rect 9331 60356 9335 60412
rect 9271 60352 9335 60356
rect 9351 60412 9415 60416
rect 9351 60356 9355 60412
rect 9355 60356 9411 60412
rect 9411 60356 9415 60412
rect 9351 60352 9415 60356
rect 4215 59868 4279 59872
rect 4215 59812 4219 59868
rect 4219 59812 4275 59868
rect 4275 59812 4279 59868
rect 4215 59808 4279 59812
rect 4295 59868 4359 59872
rect 4295 59812 4299 59868
rect 4299 59812 4355 59868
rect 4355 59812 4359 59868
rect 4295 59808 4359 59812
rect 4375 59868 4439 59872
rect 4375 59812 4379 59868
rect 4379 59812 4435 59868
rect 4435 59812 4439 59868
rect 4375 59808 4439 59812
rect 4455 59868 4519 59872
rect 4455 59812 4459 59868
rect 4459 59812 4515 59868
rect 4515 59812 4519 59868
rect 4455 59808 4519 59812
rect 7479 59868 7543 59872
rect 7479 59812 7483 59868
rect 7483 59812 7539 59868
rect 7539 59812 7543 59868
rect 7479 59808 7543 59812
rect 7559 59868 7623 59872
rect 7559 59812 7563 59868
rect 7563 59812 7619 59868
rect 7619 59812 7623 59868
rect 7559 59808 7623 59812
rect 7639 59868 7703 59872
rect 7639 59812 7643 59868
rect 7643 59812 7699 59868
rect 7699 59812 7703 59868
rect 7639 59808 7703 59812
rect 7719 59868 7783 59872
rect 7719 59812 7723 59868
rect 7723 59812 7779 59868
rect 7779 59812 7783 59868
rect 7719 59808 7783 59812
rect 3372 59468 3436 59532
rect 2584 59324 2648 59328
rect 2584 59268 2588 59324
rect 2588 59268 2644 59324
rect 2644 59268 2648 59324
rect 2584 59264 2648 59268
rect 2664 59324 2728 59328
rect 2664 59268 2668 59324
rect 2668 59268 2724 59324
rect 2724 59268 2728 59324
rect 2664 59264 2728 59268
rect 2744 59324 2808 59328
rect 2744 59268 2748 59324
rect 2748 59268 2804 59324
rect 2804 59268 2808 59324
rect 2744 59264 2808 59268
rect 2824 59324 2888 59328
rect 2824 59268 2828 59324
rect 2828 59268 2884 59324
rect 2884 59268 2888 59324
rect 2824 59264 2888 59268
rect 5847 59324 5911 59328
rect 5847 59268 5851 59324
rect 5851 59268 5907 59324
rect 5907 59268 5911 59324
rect 5847 59264 5911 59268
rect 5927 59324 5991 59328
rect 5927 59268 5931 59324
rect 5931 59268 5987 59324
rect 5987 59268 5991 59324
rect 5927 59264 5991 59268
rect 6007 59324 6071 59328
rect 6007 59268 6011 59324
rect 6011 59268 6067 59324
rect 6067 59268 6071 59324
rect 6007 59264 6071 59268
rect 6087 59324 6151 59328
rect 6087 59268 6091 59324
rect 6091 59268 6147 59324
rect 6147 59268 6151 59324
rect 6087 59264 6151 59268
rect 9111 59324 9175 59328
rect 9111 59268 9115 59324
rect 9115 59268 9171 59324
rect 9171 59268 9175 59324
rect 9111 59264 9175 59268
rect 9191 59324 9255 59328
rect 9191 59268 9195 59324
rect 9195 59268 9251 59324
rect 9251 59268 9255 59324
rect 9191 59264 9255 59268
rect 9271 59324 9335 59328
rect 9271 59268 9275 59324
rect 9275 59268 9331 59324
rect 9331 59268 9335 59324
rect 9271 59264 9335 59268
rect 9351 59324 9415 59328
rect 9351 59268 9355 59324
rect 9355 59268 9411 59324
rect 9411 59268 9415 59324
rect 9351 59264 9415 59268
rect 4215 58780 4279 58784
rect 4215 58724 4219 58780
rect 4219 58724 4275 58780
rect 4275 58724 4279 58780
rect 4215 58720 4279 58724
rect 4295 58780 4359 58784
rect 4295 58724 4299 58780
rect 4299 58724 4355 58780
rect 4355 58724 4359 58780
rect 4295 58720 4359 58724
rect 4375 58780 4439 58784
rect 4375 58724 4379 58780
rect 4379 58724 4435 58780
rect 4435 58724 4439 58780
rect 4375 58720 4439 58724
rect 4455 58780 4519 58784
rect 4455 58724 4459 58780
rect 4459 58724 4515 58780
rect 4515 58724 4519 58780
rect 4455 58720 4519 58724
rect 7479 58780 7543 58784
rect 7479 58724 7483 58780
rect 7483 58724 7539 58780
rect 7539 58724 7543 58780
rect 7479 58720 7543 58724
rect 7559 58780 7623 58784
rect 7559 58724 7563 58780
rect 7563 58724 7619 58780
rect 7619 58724 7623 58780
rect 7559 58720 7623 58724
rect 7639 58780 7703 58784
rect 7639 58724 7643 58780
rect 7643 58724 7699 58780
rect 7699 58724 7703 58780
rect 7639 58720 7703 58724
rect 7719 58780 7783 58784
rect 7719 58724 7723 58780
rect 7723 58724 7779 58780
rect 7779 58724 7783 58780
rect 7719 58720 7783 58724
rect 2584 58236 2648 58240
rect 2584 58180 2588 58236
rect 2588 58180 2644 58236
rect 2644 58180 2648 58236
rect 2584 58176 2648 58180
rect 2664 58236 2728 58240
rect 2664 58180 2668 58236
rect 2668 58180 2724 58236
rect 2724 58180 2728 58236
rect 2664 58176 2728 58180
rect 2744 58236 2808 58240
rect 2744 58180 2748 58236
rect 2748 58180 2804 58236
rect 2804 58180 2808 58236
rect 2744 58176 2808 58180
rect 2824 58236 2888 58240
rect 2824 58180 2828 58236
rect 2828 58180 2884 58236
rect 2884 58180 2888 58236
rect 2824 58176 2888 58180
rect 5847 58236 5911 58240
rect 5847 58180 5851 58236
rect 5851 58180 5907 58236
rect 5907 58180 5911 58236
rect 5847 58176 5911 58180
rect 5927 58236 5991 58240
rect 5927 58180 5931 58236
rect 5931 58180 5987 58236
rect 5987 58180 5991 58236
rect 5927 58176 5991 58180
rect 6007 58236 6071 58240
rect 6007 58180 6011 58236
rect 6011 58180 6067 58236
rect 6067 58180 6071 58236
rect 6007 58176 6071 58180
rect 6087 58236 6151 58240
rect 6087 58180 6091 58236
rect 6091 58180 6147 58236
rect 6147 58180 6151 58236
rect 6087 58176 6151 58180
rect 9111 58236 9175 58240
rect 9111 58180 9115 58236
rect 9115 58180 9171 58236
rect 9171 58180 9175 58236
rect 9111 58176 9175 58180
rect 9191 58236 9255 58240
rect 9191 58180 9195 58236
rect 9195 58180 9251 58236
rect 9251 58180 9255 58236
rect 9191 58176 9255 58180
rect 9271 58236 9335 58240
rect 9271 58180 9275 58236
rect 9275 58180 9331 58236
rect 9331 58180 9335 58236
rect 9271 58176 9335 58180
rect 9351 58236 9415 58240
rect 9351 58180 9355 58236
rect 9355 58180 9411 58236
rect 9411 58180 9415 58236
rect 9351 58176 9415 58180
rect 4215 57692 4279 57696
rect 4215 57636 4219 57692
rect 4219 57636 4275 57692
rect 4275 57636 4279 57692
rect 4215 57632 4279 57636
rect 4295 57692 4359 57696
rect 4295 57636 4299 57692
rect 4299 57636 4355 57692
rect 4355 57636 4359 57692
rect 4295 57632 4359 57636
rect 4375 57692 4439 57696
rect 4375 57636 4379 57692
rect 4379 57636 4435 57692
rect 4435 57636 4439 57692
rect 4375 57632 4439 57636
rect 4455 57692 4519 57696
rect 4455 57636 4459 57692
rect 4459 57636 4515 57692
rect 4515 57636 4519 57692
rect 4455 57632 4519 57636
rect 7479 57692 7543 57696
rect 7479 57636 7483 57692
rect 7483 57636 7539 57692
rect 7539 57636 7543 57692
rect 7479 57632 7543 57636
rect 7559 57692 7623 57696
rect 7559 57636 7563 57692
rect 7563 57636 7619 57692
rect 7619 57636 7623 57692
rect 7559 57632 7623 57636
rect 7639 57692 7703 57696
rect 7639 57636 7643 57692
rect 7643 57636 7699 57692
rect 7699 57636 7703 57692
rect 7639 57632 7703 57636
rect 7719 57692 7783 57696
rect 7719 57636 7723 57692
rect 7723 57636 7779 57692
rect 7779 57636 7783 57692
rect 7719 57632 7783 57636
rect 2584 57148 2648 57152
rect 2584 57092 2588 57148
rect 2588 57092 2644 57148
rect 2644 57092 2648 57148
rect 2584 57088 2648 57092
rect 2664 57148 2728 57152
rect 2664 57092 2668 57148
rect 2668 57092 2724 57148
rect 2724 57092 2728 57148
rect 2664 57088 2728 57092
rect 2744 57148 2808 57152
rect 2744 57092 2748 57148
rect 2748 57092 2804 57148
rect 2804 57092 2808 57148
rect 2744 57088 2808 57092
rect 2824 57148 2888 57152
rect 2824 57092 2828 57148
rect 2828 57092 2884 57148
rect 2884 57092 2888 57148
rect 2824 57088 2888 57092
rect 5847 57148 5911 57152
rect 5847 57092 5851 57148
rect 5851 57092 5907 57148
rect 5907 57092 5911 57148
rect 5847 57088 5911 57092
rect 5927 57148 5991 57152
rect 5927 57092 5931 57148
rect 5931 57092 5987 57148
rect 5987 57092 5991 57148
rect 5927 57088 5991 57092
rect 6007 57148 6071 57152
rect 6007 57092 6011 57148
rect 6011 57092 6067 57148
rect 6067 57092 6071 57148
rect 6007 57088 6071 57092
rect 6087 57148 6151 57152
rect 6087 57092 6091 57148
rect 6091 57092 6147 57148
rect 6147 57092 6151 57148
rect 6087 57088 6151 57092
rect 9111 57148 9175 57152
rect 9111 57092 9115 57148
rect 9115 57092 9171 57148
rect 9171 57092 9175 57148
rect 9111 57088 9175 57092
rect 9191 57148 9255 57152
rect 9191 57092 9195 57148
rect 9195 57092 9251 57148
rect 9251 57092 9255 57148
rect 9191 57088 9255 57092
rect 9271 57148 9335 57152
rect 9271 57092 9275 57148
rect 9275 57092 9331 57148
rect 9331 57092 9335 57148
rect 9271 57088 9335 57092
rect 9351 57148 9415 57152
rect 9351 57092 9355 57148
rect 9355 57092 9411 57148
rect 9411 57092 9415 57148
rect 9351 57088 9415 57092
rect 4215 56604 4279 56608
rect 4215 56548 4219 56604
rect 4219 56548 4275 56604
rect 4275 56548 4279 56604
rect 4215 56544 4279 56548
rect 4295 56604 4359 56608
rect 4295 56548 4299 56604
rect 4299 56548 4355 56604
rect 4355 56548 4359 56604
rect 4295 56544 4359 56548
rect 4375 56604 4439 56608
rect 4375 56548 4379 56604
rect 4379 56548 4435 56604
rect 4435 56548 4439 56604
rect 4375 56544 4439 56548
rect 4455 56604 4519 56608
rect 4455 56548 4459 56604
rect 4459 56548 4515 56604
rect 4515 56548 4519 56604
rect 4455 56544 4519 56548
rect 7479 56604 7543 56608
rect 7479 56548 7483 56604
rect 7483 56548 7539 56604
rect 7539 56548 7543 56604
rect 7479 56544 7543 56548
rect 7559 56604 7623 56608
rect 7559 56548 7563 56604
rect 7563 56548 7619 56604
rect 7619 56548 7623 56604
rect 7559 56544 7623 56548
rect 7639 56604 7703 56608
rect 7639 56548 7643 56604
rect 7643 56548 7699 56604
rect 7699 56548 7703 56604
rect 7639 56544 7703 56548
rect 7719 56604 7783 56608
rect 7719 56548 7723 56604
rect 7723 56548 7779 56604
rect 7779 56548 7783 56604
rect 7719 56544 7783 56548
rect 10732 56204 10796 56268
rect 2584 56060 2648 56064
rect 2584 56004 2588 56060
rect 2588 56004 2644 56060
rect 2644 56004 2648 56060
rect 2584 56000 2648 56004
rect 2664 56060 2728 56064
rect 2664 56004 2668 56060
rect 2668 56004 2724 56060
rect 2724 56004 2728 56060
rect 2664 56000 2728 56004
rect 2744 56060 2808 56064
rect 2744 56004 2748 56060
rect 2748 56004 2804 56060
rect 2804 56004 2808 56060
rect 2744 56000 2808 56004
rect 2824 56060 2888 56064
rect 2824 56004 2828 56060
rect 2828 56004 2884 56060
rect 2884 56004 2888 56060
rect 2824 56000 2888 56004
rect 5847 56060 5911 56064
rect 5847 56004 5851 56060
rect 5851 56004 5907 56060
rect 5907 56004 5911 56060
rect 5847 56000 5911 56004
rect 5927 56060 5991 56064
rect 5927 56004 5931 56060
rect 5931 56004 5987 56060
rect 5987 56004 5991 56060
rect 5927 56000 5991 56004
rect 6007 56060 6071 56064
rect 6007 56004 6011 56060
rect 6011 56004 6067 56060
rect 6067 56004 6071 56060
rect 6007 56000 6071 56004
rect 6087 56060 6151 56064
rect 6087 56004 6091 56060
rect 6091 56004 6147 56060
rect 6147 56004 6151 56060
rect 6087 56000 6151 56004
rect 9111 56060 9175 56064
rect 9111 56004 9115 56060
rect 9115 56004 9171 56060
rect 9171 56004 9175 56060
rect 9111 56000 9175 56004
rect 9191 56060 9255 56064
rect 9191 56004 9195 56060
rect 9195 56004 9251 56060
rect 9251 56004 9255 56060
rect 9191 56000 9255 56004
rect 9271 56060 9335 56064
rect 9271 56004 9275 56060
rect 9275 56004 9331 56060
rect 9331 56004 9335 56060
rect 9271 56000 9335 56004
rect 9351 56060 9415 56064
rect 9351 56004 9355 56060
rect 9355 56004 9411 56060
rect 9411 56004 9415 56060
rect 9351 56000 9415 56004
rect 7972 55796 8036 55860
rect 4215 55516 4279 55520
rect 4215 55460 4219 55516
rect 4219 55460 4275 55516
rect 4275 55460 4279 55516
rect 4215 55456 4279 55460
rect 4295 55516 4359 55520
rect 4295 55460 4299 55516
rect 4299 55460 4355 55516
rect 4355 55460 4359 55516
rect 4295 55456 4359 55460
rect 4375 55516 4439 55520
rect 4375 55460 4379 55516
rect 4379 55460 4435 55516
rect 4435 55460 4439 55516
rect 4375 55456 4439 55460
rect 4455 55516 4519 55520
rect 4455 55460 4459 55516
rect 4459 55460 4515 55516
rect 4515 55460 4519 55516
rect 4455 55456 4519 55460
rect 7479 55516 7543 55520
rect 7479 55460 7483 55516
rect 7483 55460 7539 55516
rect 7539 55460 7543 55516
rect 7479 55456 7543 55460
rect 7559 55516 7623 55520
rect 7559 55460 7563 55516
rect 7563 55460 7619 55516
rect 7619 55460 7623 55516
rect 7559 55456 7623 55460
rect 7639 55516 7703 55520
rect 7639 55460 7643 55516
rect 7643 55460 7699 55516
rect 7699 55460 7703 55516
rect 7639 55456 7703 55460
rect 7719 55516 7783 55520
rect 7719 55460 7723 55516
rect 7723 55460 7779 55516
rect 7779 55460 7783 55516
rect 7719 55456 7783 55460
rect 2584 54972 2648 54976
rect 2584 54916 2588 54972
rect 2588 54916 2644 54972
rect 2644 54916 2648 54972
rect 2584 54912 2648 54916
rect 2664 54972 2728 54976
rect 2664 54916 2668 54972
rect 2668 54916 2724 54972
rect 2724 54916 2728 54972
rect 2664 54912 2728 54916
rect 2744 54972 2808 54976
rect 2744 54916 2748 54972
rect 2748 54916 2804 54972
rect 2804 54916 2808 54972
rect 2744 54912 2808 54916
rect 2824 54972 2888 54976
rect 2824 54916 2828 54972
rect 2828 54916 2884 54972
rect 2884 54916 2888 54972
rect 2824 54912 2888 54916
rect 5847 54972 5911 54976
rect 5847 54916 5851 54972
rect 5851 54916 5907 54972
rect 5907 54916 5911 54972
rect 5847 54912 5911 54916
rect 5927 54972 5991 54976
rect 5927 54916 5931 54972
rect 5931 54916 5987 54972
rect 5987 54916 5991 54972
rect 5927 54912 5991 54916
rect 6007 54972 6071 54976
rect 6007 54916 6011 54972
rect 6011 54916 6067 54972
rect 6067 54916 6071 54972
rect 6007 54912 6071 54916
rect 6087 54972 6151 54976
rect 6087 54916 6091 54972
rect 6091 54916 6147 54972
rect 6147 54916 6151 54972
rect 6087 54912 6151 54916
rect 9111 54972 9175 54976
rect 9111 54916 9115 54972
rect 9115 54916 9171 54972
rect 9171 54916 9175 54972
rect 9111 54912 9175 54916
rect 9191 54972 9255 54976
rect 9191 54916 9195 54972
rect 9195 54916 9251 54972
rect 9251 54916 9255 54972
rect 9191 54912 9255 54916
rect 9271 54972 9335 54976
rect 9271 54916 9275 54972
rect 9275 54916 9331 54972
rect 9331 54916 9335 54972
rect 9271 54912 9335 54916
rect 9351 54972 9415 54976
rect 9351 54916 9355 54972
rect 9355 54916 9411 54972
rect 9411 54916 9415 54972
rect 9351 54912 9415 54916
rect 4215 54428 4279 54432
rect 4215 54372 4219 54428
rect 4219 54372 4275 54428
rect 4275 54372 4279 54428
rect 4215 54368 4279 54372
rect 4295 54428 4359 54432
rect 4295 54372 4299 54428
rect 4299 54372 4355 54428
rect 4355 54372 4359 54428
rect 4295 54368 4359 54372
rect 4375 54428 4439 54432
rect 4375 54372 4379 54428
rect 4379 54372 4435 54428
rect 4435 54372 4439 54428
rect 4375 54368 4439 54372
rect 4455 54428 4519 54432
rect 4455 54372 4459 54428
rect 4459 54372 4515 54428
rect 4515 54372 4519 54428
rect 4455 54368 4519 54372
rect 7479 54428 7543 54432
rect 7479 54372 7483 54428
rect 7483 54372 7539 54428
rect 7539 54372 7543 54428
rect 7479 54368 7543 54372
rect 7559 54428 7623 54432
rect 7559 54372 7563 54428
rect 7563 54372 7619 54428
rect 7619 54372 7623 54428
rect 7559 54368 7623 54372
rect 7639 54428 7703 54432
rect 7639 54372 7643 54428
rect 7643 54372 7699 54428
rect 7699 54372 7703 54428
rect 7639 54368 7703 54372
rect 7719 54428 7783 54432
rect 7719 54372 7723 54428
rect 7723 54372 7779 54428
rect 7779 54372 7783 54428
rect 7719 54368 7783 54372
rect 11468 54300 11532 54364
rect 2584 53884 2648 53888
rect 2584 53828 2588 53884
rect 2588 53828 2644 53884
rect 2644 53828 2648 53884
rect 2584 53824 2648 53828
rect 2664 53884 2728 53888
rect 2664 53828 2668 53884
rect 2668 53828 2724 53884
rect 2724 53828 2728 53884
rect 2664 53824 2728 53828
rect 2744 53884 2808 53888
rect 2744 53828 2748 53884
rect 2748 53828 2804 53884
rect 2804 53828 2808 53884
rect 2744 53824 2808 53828
rect 2824 53884 2888 53888
rect 2824 53828 2828 53884
rect 2828 53828 2884 53884
rect 2884 53828 2888 53884
rect 2824 53824 2888 53828
rect 5847 53884 5911 53888
rect 5847 53828 5851 53884
rect 5851 53828 5907 53884
rect 5907 53828 5911 53884
rect 5847 53824 5911 53828
rect 5927 53884 5991 53888
rect 5927 53828 5931 53884
rect 5931 53828 5987 53884
rect 5987 53828 5991 53884
rect 5927 53824 5991 53828
rect 6007 53884 6071 53888
rect 6007 53828 6011 53884
rect 6011 53828 6067 53884
rect 6067 53828 6071 53884
rect 6007 53824 6071 53828
rect 6087 53884 6151 53888
rect 6087 53828 6091 53884
rect 6091 53828 6147 53884
rect 6147 53828 6151 53884
rect 6087 53824 6151 53828
rect 9111 53884 9175 53888
rect 9111 53828 9115 53884
rect 9115 53828 9171 53884
rect 9171 53828 9175 53884
rect 9111 53824 9175 53828
rect 9191 53884 9255 53888
rect 9191 53828 9195 53884
rect 9195 53828 9251 53884
rect 9251 53828 9255 53884
rect 9191 53824 9255 53828
rect 9271 53884 9335 53888
rect 9271 53828 9275 53884
rect 9275 53828 9331 53884
rect 9331 53828 9335 53884
rect 9271 53824 9335 53828
rect 9351 53884 9415 53888
rect 9351 53828 9355 53884
rect 9355 53828 9411 53884
rect 9411 53828 9415 53884
rect 9351 53824 9415 53828
rect 8156 53484 8220 53548
rect 4215 53340 4279 53344
rect 4215 53284 4219 53340
rect 4219 53284 4275 53340
rect 4275 53284 4279 53340
rect 4215 53280 4279 53284
rect 4295 53340 4359 53344
rect 4295 53284 4299 53340
rect 4299 53284 4355 53340
rect 4355 53284 4359 53340
rect 4295 53280 4359 53284
rect 4375 53340 4439 53344
rect 4375 53284 4379 53340
rect 4379 53284 4435 53340
rect 4435 53284 4439 53340
rect 4375 53280 4439 53284
rect 4455 53340 4519 53344
rect 4455 53284 4459 53340
rect 4459 53284 4515 53340
rect 4515 53284 4519 53340
rect 4455 53280 4519 53284
rect 7479 53340 7543 53344
rect 7479 53284 7483 53340
rect 7483 53284 7539 53340
rect 7539 53284 7543 53340
rect 7479 53280 7543 53284
rect 7559 53340 7623 53344
rect 7559 53284 7563 53340
rect 7563 53284 7619 53340
rect 7619 53284 7623 53340
rect 7559 53280 7623 53284
rect 7639 53340 7703 53344
rect 7639 53284 7643 53340
rect 7643 53284 7699 53340
rect 7699 53284 7703 53340
rect 7639 53280 7703 53284
rect 7719 53340 7783 53344
rect 7719 53284 7723 53340
rect 7723 53284 7779 53340
rect 7779 53284 7783 53340
rect 7719 53280 7783 53284
rect 10364 53212 10428 53276
rect 2584 52796 2648 52800
rect 2584 52740 2588 52796
rect 2588 52740 2644 52796
rect 2644 52740 2648 52796
rect 2584 52736 2648 52740
rect 2664 52796 2728 52800
rect 2664 52740 2668 52796
rect 2668 52740 2724 52796
rect 2724 52740 2728 52796
rect 2664 52736 2728 52740
rect 2744 52796 2808 52800
rect 2744 52740 2748 52796
rect 2748 52740 2804 52796
rect 2804 52740 2808 52796
rect 2744 52736 2808 52740
rect 2824 52796 2888 52800
rect 2824 52740 2828 52796
rect 2828 52740 2884 52796
rect 2884 52740 2888 52796
rect 2824 52736 2888 52740
rect 5847 52796 5911 52800
rect 5847 52740 5851 52796
rect 5851 52740 5907 52796
rect 5907 52740 5911 52796
rect 5847 52736 5911 52740
rect 5927 52796 5991 52800
rect 5927 52740 5931 52796
rect 5931 52740 5987 52796
rect 5987 52740 5991 52796
rect 5927 52736 5991 52740
rect 6007 52796 6071 52800
rect 6007 52740 6011 52796
rect 6011 52740 6067 52796
rect 6067 52740 6071 52796
rect 6007 52736 6071 52740
rect 6087 52796 6151 52800
rect 6087 52740 6091 52796
rect 6091 52740 6147 52796
rect 6147 52740 6151 52796
rect 6087 52736 6151 52740
rect 9111 52796 9175 52800
rect 9111 52740 9115 52796
rect 9115 52740 9171 52796
rect 9171 52740 9175 52796
rect 9111 52736 9175 52740
rect 9191 52796 9255 52800
rect 9191 52740 9195 52796
rect 9195 52740 9251 52796
rect 9251 52740 9255 52796
rect 9191 52736 9255 52740
rect 9271 52796 9335 52800
rect 9271 52740 9275 52796
rect 9275 52740 9331 52796
rect 9331 52740 9335 52796
rect 9271 52736 9335 52740
rect 9351 52796 9415 52800
rect 9351 52740 9355 52796
rect 9355 52740 9411 52796
rect 9411 52740 9415 52796
rect 9351 52736 9415 52740
rect 10916 52396 10980 52460
rect 4215 52252 4279 52256
rect 4215 52196 4219 52252
rect 4219 52196 4275 52252
rect 4275 52196 4279 52252
rect 4215 52192 4279 52196
rect 4295 52252 4359 52256
rect 4295 52196 4299 52252
rect 4299 52196 4355 52252
rect 4355 52196 4359 52252
rect 4295 52192 4359 52196
rect 4375 52252 4439 52256
rect 4375 52196 4379 52252
rect 4379 52196 4435 52252
rect 4435 52196 4439 52252
rect 4375 52192 4439 52196
rect 4455 52252 4519 52256
rect 4455 52196 4459 52252
rect 4459 52196 4515 52252
rect 4515 52196 4519 52252
rect 4455 52192 4519 52196
rect 7479 52252 7543 52256
rect 7479 52196 7483 52252
rect 7483 52196 7539 52252
rect 7539 52196 7543 52252
rect 7479 52192 7543 52196
rect 7559 52252 7623 52256
rect 7559 52196 7563 52252
rect 7563 52196 7619 52252
rect 7619 52196 7623 52252
rect 7559 52192 7623 52196
rect 7639 52252 7703 52256
rect 7639 52196 7643 52252
rect 7643 52196 7699 52252
rect 7699 52196 7703 52252
rect 7639 52192 7703 52196
rect 7719 52252 7783 52256
rect 7719 52196 7723 52252
rect 7723 52196 7779 52252
rect 7779 52196 7783 52252
rect 7719 52192 7783 52196
rect 2584 51708 2648 51712
rect 2584 51652 2588 51708
rect 2588 51652 2644 51708
rect 2644 51652 2648 51708
rect 2584 51648 2648 51652
rect 2664 51708 2728 51712
rect 2664 51652 2668 51708
rect 2668 51652 2724 51708
rect 2724 51652 2728 51708
rect 2664 51648 2728 51652
rect 2744 51708 2808 51712
rect 2744 51652 2748 51708
rect 2748 51652 2804 51708
rect 2804 51652 2808 51708
rect 2744 51648 2808 51652
rect 2824 51708 2888 51712
rect 2824 51652 2828 51708
rect 2828 51652 2884 51708
rect 2884 51652 2888 51708
rect 2824 51648 2888 51652
rect 5847 51708 5911 51712
rect 5847 51652 5851 51708
rect 5851 51652 5907 51708
rect 5907 51652 5911 51708
rect 5847 51648 5911 51652
rect 5927 51708 5991 51712
rect 5927 51652 5931 51708
rect 5931 51652 5987 51708
rect 5987 51652 5991 51708
rect 5927 51648 5991 51652
rect 6007 51708 6071 51712
rect 6007 51652 6011 51708
rect 6011 51652 6067 51708
rect 6067 51652 6071 51708
rect 6007 51648 6071 51652
rect 6087 51708 6151 51712
rect 6087 51652 6091 51708
rect 6091 51652 6147 51708
rect 6147 51652 6151 51708
rect 6087 51648 6151 51652
rect 9111 51708 9175 51712
rect 9111 51652 9115 51708
rect 9115 51652 9171 51708
rect 9171 51652 9175 51708
rect 9111 51648 9175 51652
rect 9191 51708 9255 51712
rect 9191 51652 9195 51708
rect 9195 51652 9251 51708
rect 9251 51652 9255 51708
rect 9191 51648 9255 51652
rect 9271 51708 9335 51712
rect 9271 51652 9275 51708
rect 9275 51652 9331 51708
rect 9331 51652 9335 51708
rect 9271 51648 9335 51652
rect 9351 51708 9415 51712
rect 9351 51652 9355 51708
rect 9355 51652 9411 51708
rect 9411 51652 9415 51708
rect 9351 51648 9415 51652
rect 7052 51444 7116 51508
rect 3188 51172 3252 51236
rect 6684 51172 6748 51236
rect 4215 51164 4279 51168
rect 4215 51108 4219 51164
rect 4219 51108 4275 51164
rect 4275 51108 4279 51164
rect 4215 51104 4279 51108
rect 4295 51164 4359 51168
rect 4295 51108 4299 51164
rect 4299 51108 4355 51164
rect 4355 51108 4359 51164
rect 4295 51104 4359 51108
rect 4375 51164 4439 51168
rect 4375 51108 4379 51164
rect 4379 51108 4435 51164
rect 4435 51108 4439 51164
rect 4375 51104 4439 51108
rect 4455 51164 4519 51168
rect 4455 51108 4459 51164
rect 4459 51108 4515 51164
rect 4515 51108 4519 51164
rect 4455 51104 4519 51108
rect 8156 51172 8220 51236
rect 7479 51164 7543 51168
rect 7479 51108 7483 51164
rect 7483 51108 7539 51164
rect 7539 51108 7543 51164
rect 7479 51104 7543 51108
rect 7559 51164 7623 51168
rect 7559 51108 7563 51164
rect 7563 51108 7619 51164
rect 7619 51108 7623 51164
rect 7559 51104 7623 51108
rect 7639 51164 7703 51168
rect 7639 51108 7643 51164
rect 7643 51108 7699 51164
rect 7699 51108 7703 51164
rect 7639 51104 7703 51108
rect 7719 51164 7783 51168
rect 7719 51108 7723 51164
rect 7723 51108 7779 51164
rect 7779 51108 7783 51164
rect 7719 51104 7783 51108
rect 3188 50960 3252 50964
rect 3188 50904 3202 50960
rect 3202 50904 3252 50960
rect 3188 50900 3252 50904
rect 3740 50900 3804 50964
rect 6684 50900 6748 50964
rect 2584 50620 2648 50624
rect 2584 50564 2588 50620
rect 2588 50564 2644 50620
rect 2644 50564 2648 50620
rect 2584 50560 2648 50564
rect 2664 50620 2728 50624
rect 2664 50564 2668 50620
rect 2668 50564 2724 50620
rect 2724 50564 2728 50620
rect 2664 50560 2728 50564
rect 2744 50620 2808 50624
rect 2744 50564 2748 50620
rect 2748 50564 2804 50620
rect 2804 50564 2808 50620
rect 2744 50560 2808 50564
rect 2824 50620 2888 50624
rect 2824 50564 2828 50620
rect 2828 50564 2884 50620
rect 2884 50564 2888 50620
rect 2824 50560 2888 50564
rect 5847 50620 5911 50624
rect 5847 50564 5851 50620
rect 5851 50564 5907 50620
rect 5907 50564 5911 50620
rect 5847 50560 5911 50564
rect 5927 50620 5991 50624
rect 5927 50564 5931 50620
rect 5931 50564 5987 50620
rect 5987 50564 5991 50620
rect 5927 50560 5991 50564
rect 6007 50620 6071 50624
rect 6007 50564 6011 50620
rect 6011 50564 6067 50620
rect 6067 50564 6071 50620
rect 6007 50560 6071 50564
rect 6087 50620 6151 50624
rect 6087 50564 6091 50620
rect 6091 50564 6147 50620
rect 6147 50564 6151 50620
rect 6087 50560 6151 50564
rect 8156 50356 8220 50420
rect 9111 50620 9175 50624
rect 9111 50564 9115 50620
rect 9115 50564 9171 50620
rect 9171 50564 9175 50620
rect 9111 50560 9175 50564
rect 9191 50620 9255 50624
rect 9191 50564 9195 50620
rect 9195 50564 9251 50620
rect 9251 50564 9255 50620
rect 9191 50560 9255 50564
rect 9271 50620 9335 50624
rect 9271 50564 9275 50620
rect 9275 50564 9331 50620
rect 9331 50564 9335 50620
rect 9271 50560 9335 50564
rect 9351 50620 9415 50624
rect 9351 50564 9355 50620
rect 9355 50564 9411 50620
rect 9411 50564 9415 50620
rect 9351 50560 9415 50564
rect 11468 50492 11532 50556
rect 10732 50084 10796 50148
rect 4215 50076 4279 50080
rect 4215 50020 4219 50076
rect 4219 50020 4275 50076
rect 4275 50020 4279 50076
rect 4215 50016 4279 50020
rect 4295 50076 4359 50080
rect 4295 50020 4299 50076
rect 4299 50020 4355 50076
rect 4355 50020 4359 50076
rect 4295 50016 4359 50020
rect 4375 50076 4439 50080
rect 4375 50020 4379 50076
rect 4379 50020 4435 50076
rect 4435 50020 4439 50076
rect 4375 50016 4439 50020
rect 4455 50076 4519 50080
rect 4455 50020 4459 50076
rect 4459 50020 4515 50076
rect 4515 50020 4519 50076
rect 4455 50016 4519 50020
rect 7479 50076 7543 50080
rect 7479 50020 7483 50076
rect 7483 50020 7539 50076
rect 7539 50020 7543 50076
rect 7479 50016 7543 50020
rect 7559 50076 7623 50080
rect 7559 50020 7563 50076
rect 7563 50020 7619 50076
rect 7619 50020 7623 50076
rect 7559 50016 7623 50020
rect 7639 50076 7703 50080
rect 7639 50020 7643 50076
rect 7643 50020 7699 50076
rect 7699 50020 7703 50076
rect 7639 50016 7703 50020
rect 7719 50076 7783 50080
rect 7719 50020 7723 50076
rect 7723 50020 7779 50076
rect 7779 50020 7783 50076
rect 7719 50016 7783 50020
rect 2584 49532 2648 49536
rect 2584 49476 2588 49532
rect 2588 49476 2644 49532
rect 2644 49476 2648 49532
rect 2584 49472 2648 49476
rect 2664 49532 2728 49536
rect 2664 49476 2668 49532
rect 2668 49476 2724 49532
rect 2724 49476 2728 49532
rect 2664 49472 2728 49476
rect 2744 49532 2808 49536
rect 2744 49476 2748 49532
rect 2748 49476 2804 49532
rect 2804 49476 2808 49532
rect 2744 49472 2808 49476
rect 2824 49532 2888 49536
rect 2824 49476 2828 49532
rect 2828 49476 2884 49532
rect 2884 49476 2888 49532
rect 2824 49472 2888 49476
rect 7052 49600 7116 49604
rect 7052 49544 7066 49600
rect 7066 49544 7116 49600
rect 7052 49540 7116 49544
rect 5847 49532 5911 49536
rect 5847 49476 5851 49532
rect 5851 49476 5907 49532
rect 5907 49476 5911 49532
rect 5847 49472 5911 49476
rect 5927 49532 5991 49536
rect 5927 49476 5931 49532
rect 5931 49476 5987 49532
rect 5987 49476 5991 49532
rect 5927 49472 5991 49476
rect 6007 49532 6071 49536
rect 6007 49476 6011 49532
rect 6011 49476 6067 49532
rect 6067 49476 6071 49532
rect 6007 49472 6071 49476
rect 6087 49532 6151 49536
rect 6087 49476 6091 49532
rect 6091 49476 6147 49532
rect 6147 49476 6151 49532
rect 6087 49472 6151 49476
rect 9111 49532 9175 49536
rect 9111 49476 9115 49532
rect 9115 49476 9171 49532
rect 9171 49476 9175 49532
rect 9111 49472 9175 49476
rect 9191 49532 9255 49536
rect 9191 49476 9195 49532
rect 9195 49476 9251 49532
rect 9251 49476 9255 49532
rect 9191 49472 9255 49476
rect 9271 49532 9335 49536
rect 9271 49476 9275 49532
rect 9275 49476 9331 49532
rect 9331 49476 9335 49532
rect 9271 49472 9335 49476
rect 9351 49532 9415 49536
rect 9351 49476 9355 49532
rect 9355 49476 9411 49532
rect 9411 49476 9415 49532
rect 9351 49472 9415 49476
rect 4215 48988 4279 48992
rect 4215 48932 4219 48988
rect 4219 48932 4275 48988
rect 4275 48932 4279 48988
rect 4215 48928 4279 48932
rect 4295 48988 4359 48992
rect 4295 48932 4299 48988
rect 4299 48932 4355 48988
rect 4355 48932 4359 48988
rect 4295 48928 4359 48932
rect 4375 48988 4439 48992
rect 4375 48932 4379 48988
rect 4379 48932 4435 48988
rect 4435 48932 4439 48988
rect 4375 48928 4439 48932
rect 4455 48988 4519 48992
rect 4455 48932 4459 48988
rect 4459 48932 4515 48988
rect 4515 48932 4519 48988
rect 4455 48928 4519 48932
rect 7479 48988 7543 48992
rect 7479 48932 7483 48988
rect 7483 48932 7539 48988
rect 7539 48932 7543 48988
rect 7479 48928 7543 48932
rect 7559 48988 7623 48992
rect 7559 48932 7563 48988
rect 7563 48932 7619 48988
rect 7619 48932 7623 48988
rect 7559 48928 7623 48932
rect 7639 48988 7703 48992
rect 7639 48932 7643 48988
rect 7643 48932 7699 48988
rect 7699 48932 7703 48988
rect 7639 48928 7703 48932
rect 7719 48988 7783 48992
rect 7719 48932 7723 48988
rect 7723 48932 7779 48988
rect 7779 48932 7783 48988
rect 7719 48928 7783 48932
rect 8156 48724 8220 48788
rect 7972 48452 8036 48516
rect 2584 48444 2648 48448
rect 2584 48388 2588 48444
rect 2588 48388 2644 48444
rect 2644 48388 2648 48444
rect 2584 48384 2648 48388
rect 2664 48444 2728 48448
rect 2664 48388 2668 48444
rect 2668 48388 2724 48444
rect 2724 48388 2728 48444
rect 2664 48384 2728 48388
rect 2744 48444 2808 48448
rect 2744 48388 2748 48444
rect 2748 48388 2804 48444
rect 2804 48388 2808 48444
rect 2744 48384 2808 48388
rect 2824 48444 2888 48448
rect 2824 48388 2828 48444
rect 2828 48388 2884 48444
rect 2884 48388 2888 48444
rect 2824 48384 2888 48388
rect 5847 48444 5911 48448
rect 5847 48388 5851 48444
rect 5851 48388 5907 48444
rect 5907 48388 5911 48444
rect 5847 48384 5911 48388
rect 5927 48444 5991 48448
rect 5927 48388 5931 48444
rect 5931 48388 5987 48444
rect 5987 48388 5991 48444
rect 5927 48384 5991 48388
rect 6007 48444 6071 48448
rect 6007 48388 6011 48444
rect 6011 48388 6067 48444
rect 6067 48388 6071 48444
rect 6007 48384 6071 48388
rect 6087 48444 6151 48448
rect 6087 48388 6091 48444
rect 6091 48388 6147 48444
rect 6147 48388 6151 48444
rect 6087 48384 6151 48388
rect 9111 48444 9175 48448
rect 9111 48388 9115 48444
rect 9115 48388 9171 48444
rect 9171 48388 9175 48444
rect 9111 48384 9175 48388
rect 9191 48444 9255 48448
rect 9191 48388 9195 48444
rect 9195 48388 9251 48444
rect 9251 48388 9255 48444
rect 9191 48384 9255 48388
rect 9271 48444 9335 48448
rect 9271 48388 9275 48444
rect 9275 48388 9331 48444
rect 9331 48388 9335 48444
rect 9271 48384 9335 48388
rect 9351 48444 9415 48448
rect 9351 48388 9355 48444
rect 9355 48388 9411 48444
rect 9411 48388 9415 48444
rect 9351 48384 9415 48388
rect 7236 48044 7300 48108
rect 4215 47900 4279 47904
rect 4215 47844 4219 47900
rect 4219 47844 4275 47900
rect 4275 47844 4279 47900
rect 4215 47840 4279 47844
rect 4295 47900 4359 47904
rect 4295 47844 4299 47900
rect 4299 47844 4355 47900
rect 4355 47844 4359 47900
rect 4295 47840 4359 47844
rect 4375 47900 4439 47904
rect 4375 47844 4379 47900
rect 4379 47844 4435 47900
rect 4435 47844 4439 47900
rect 4375 47840 4439 47844
rect 4455 47900 4519 47904
rect 4455 47844 4459 47900
rect 4459 47844 4515 47900
rect 4515 47844 4519 47900
rect 4455 47840 4519 47844
rect 7479 47900 7543 47904
rect 7479 47844 7483 47900
rect 7483 47844 7539 47900
rect 7539 47844 7543 47900
rect 7479 47840 7543 47844
rect 7559 47900 7623 47904
rect 7559 47844 7563 47900
rect 7563 47844 7619 47900
rect 7619 47844 7623 47900
rect 7559 47840 7623 47844
rect 7639 47900 7703 47904
rect 7639 47844 7643 47900
rect 7643 47844 7699 47900
rect 7699 47844 7703 47900
rect 7639 47840 7703 47844
rect 7719 47900 7783 47904
rect 7719 47844 7723 47900
rect 7723 47844 7779 47900
rect 7779 47844 7783 47900
rect 7719 47840 7783 47844
rect 8156 47636 8220 47700
rect 2584 47356 2648 47360
rect 2584 47300 2588 47356
rect 2588 47300 2644 47356
rect 2644 47300 2648 47356
rect 2584 47296 2648 47300
rect 2664 47356 2728 47360
rect 2664 47300 2668 47356
rect 2668 47300 2724 47356
rect 2724 47300 2728 47356
rect 2664 47296 2728 47300
rect 2744 47356 2808 47360
rect 2744 47300 2748 47356
rect 2748 47300 2804 47356
rect 2804 47300 2808 47356
rect 2744 47296 2808 47300
rect 2824 47356 2888 47360
rect 2824 47300 2828 47356
rect 2828 47300 2884 47356
rect 2884 47300 2888 47356
rect 2824 47296 2888 47300
rect 5847 47356 5911 47360
rect 5847 47300 5851 47356
rect 5851 47300 5907 47356
rect 5907 47300 5911 47356
rect 5847 47296 5911 47300
rect 5927 47356 5991 47360
rect 5927 47300 5931 47356
rect 5931 47300 5987 47356
rect 5987 47300 5991 47356
rect 5927 47296 5991 47300
rect 6007 47356 6071 47360
rect 6007 47300 6011 47356
rect 6011 47300 6067 47356
rect 6067 47300 6071 47356
rect 6007 47296 6071 47300
rect 6087 47356 6151 47360
rect 6087 47300 6091 47356
rect 6091 47300 6147 47356
rect 6147 47300 6151 47356
rect 6087 47296 6151 47300
rect 9111 47356 9175 47360
rect 9111 47300 9115 47356
rect 9115 47300 9171 47356
rect 9171 47300 9175 47356
rect 9111 47296 9175 47300
rect 9191 47356 9255 47360
rect 9191 47300 9195 47356
rect 9195 47300 9251 47356
rect 9251 47300 9255 47356
rect 9191 47296 9255 47300
rect 9271 47356 9335 47360
rect 9271 47300 9275 47356
rect 9275 47300 9331 47356
rect 9331 47300 9335 47356
rect 9271 47296 9335 47300
rect 9351 47356 9415 47360
rect 9351 47300 9355 47356
rect 9355 47300 9411 47356
rect 9411 47300 9415 47356
rect 9351 47296 9415 47300
rect 4215 46812 4279 46816
rect 4215 46756 4219 46812
rect 4219 46756 4275 46812
rect 4275 46756 4279 46812
rect 4215 46752 4279 46756
rect 4295 46812 4359 46816
rect 4295 46756 4299 46812
rect 4299 46756 4355 46812
rect 4355 46756 4359 46812
rect 4295 46752 4359 46756
rect 4375 46812 4439 46816
rect 4375 46756 4379 46812
rect 4379 46756 4435 46812
rect 4435 46756 4439 46812
rect 4375 46752 4439 46756
rect 4455 46812 4519 46816
rect 4455 46756 4459 46812
rect 4459 46756 4515 46812
rect 4515 46756 4519 46812
rect 4455 46752 4519 46756
rect 7479 46812 7543 46816
rect 7479 46756 7483 46812
rect 7483 46756 7539 46812
rect 7539 46756 7543 46812
rect 7479 46752 7543 46756
rect 7559 46812 7623 46816
rect 7559 46756 7563 46812
rect 7563 46756 7619 46812
rect 7619 46756 7623 46812
rect 7559 46752 7623 46756
rect 7639 46812 7703 46816
rect 7639 46756 7643 46812
rect 7643 46756 7699 46812
rect 7699 46756 7703 46812
rect 7639 46752 7703 46756
rect 7719 46812 7783 46816
rect 7719 46756 7723 46812
rect 7723 46756 7779 46812
rect 7779 46756 7783 46812
rect 7719 46752 7783 46756
rect 2584 46268 2648 46272
rect 2584 46212 2588 46268
rect 2588 46212 2644 46268
rect 2644 46212 2648 46268
rect 2584 46208 2648 46212
rect 2664 46268 2728 46272
rect 2664 46212 2668 46268
rect 2668 46212 2724 46268
rect 2724 46212 2728 46268
rect 2664 46208 2728 46212
rect 2744 46268 2808 46272
rect 2744 46212 2748 46268
rect 2748 46212 2804 46268
rect 2804 46212 2808 46268
rect 2744 46208 2808 46212
rect 2824 46268 2888 46272
rect 2824 46212 2828 46268
rect 2828 46212 2884 46268
rect 2884 46212 2888 46268
rect 2824 46208 2888 46212
rect 5847 46268 5911 46272
rect 5847 46212 5851 46268
rect 5851 46212 5907 46268
rect 5907 46212 5911 46268
rect 5847 46208 5911 46212
rect 5927 46268 5991 46272
rect 5927 46212 5931 46268
rect 5931 46212 5987 46268
rect 5987 46212 5991 46268
rect 5927 46208 5991 46212
rect 6007 46268 6071 46272
rect 6007 46212 6011 46268
rect 6011 46212 6067 46268
rect 6067 46212 6071 46268
rect 6007 46208 6071 46212
rect 6087 46268 6151 46272
rect 6087 46212 6091 46268
rect 6091 46212 6147 46268
rect 6147 46212 6151 46268
rect 6087 46208 6151 46212
rect 9111 46268 9175 46272
rect 9111 46212 9115 46268
rect 9115 46212 9171 46268
rect 9171 46212 9175 46268
rect 9111 46208 9175 46212
rect 9191 46268 9255 46272
rect 9191 46212 9195 46268
rect 9195 46212 9251 46268
rect 9251 46212 9255 46268
rect 9191 46208 9255 46212
rect 9271 46268 9335 46272
rect 9271 46212 9275 46268
rect 9275 46212 9331 46268
rect 9331 46212 9335 46268
rect 9271 46208 9335 46212
rect 9351 46268 9415 46272
rect 9351 46212 9355 46268
rect 9355 46212 9411 46268
rect 9411 46212 9415 46268
rect 9351 46208 9415 46212
rect 9996 46336 10060 46340
rect 9996 46280 10010 46336
rect 10010 46280 10060 46336
rect 9996 46276 10060 46280
rect 4215 45724 4279 45728
rect 4215 45668 4219 45724
rect 4219 45668 4275 45724
rect 4275 45668 4279 45724
rect 4215 45664 4279 45668
rect 4295 45724 4359 45728
rect 4295 45668 4299 45724
rect 4299 45668 4355 45724
rect 4355 45668 4359 45724
rect 4295 45664 4359 45668
rect 4375 45724 4439 45728
rect 4375 45668 4379 45724
rect 4379 45668 4435 45724
rect 4435 45668 4439 45724
rect 4375 45664 4439 45668
rect 4455 45724 4519 45728
rect 4455 45668 4459 45724
rect 4459 45668 4515 45724
rect 4515 45668 4519 45724
rect 4455 45664 4519 45668
rect 7479 45724 7543 45728
rect 7479 45668 7483 45724
rect 7483 45668 7539 45724
rect 7539 45668 7543 45724
rect 7479 45664 7543 45668
rect 7559 45724 7623 45728
rect 7559 45668 7563 45724
rect 7563 45668 7619 45724
rect 7619 45668 7623 45724
rect 7559 45664 7623 45668
rect 7639 45724 7703 45728
rect 7639 45668 7643 45724
rect 7643 45668 7699 45724
rect 7699 45668 7703 45724
rect 7639 45664 7703 45668
rect 7719 45724 7783 45728
rect 7719 45668 7723 45724
rect 7723 45668 7779 45724
rect 7779 45668 7783 45724
rect 7719 45664 7783 45668
rect 3740 45384 3804 45388
rect 3740 45328 3790 45384
rect 3790 45328 3804 45384
rect 3740 45324 3804 45328
rect 2584 45180 2648 45184
rect 2584 45124 2588 45180
rect 2588 45124 2644 45180
rect 2644 45124 2648 45180
rect 2584 45120 2648 45124
rect 2664 45180 2728 45184
rect 2664 45124 2668 45180
rect 2668 45124 2724 45180
rect 2724 45124 2728 45180
rect 2664 45120 2728 45124
rect 2744 45180 2808 45184
rect 2744 45124 2748 45180
rect 2748 45124 2804 45180
rect 2804 45124 2808 45180
rect 2744 45120 2808 45124
rect 2824 45180 2888 45184
rect 2824 45124 2828 45180
rect 2828 45124 2884 45180
rect 2884 45124 2888 45180
rect 2824 45120 2888 45124
rect 5847 45180 5911 45184
rect 5847 45124 5851 45180
rect 5851 45124 5907 45180
rect 5907 45124 5911 45180
rect 5847 45120 5911 45124
rect 5927 45180 5991 45184
rect 5927 45124 5931 45180
rect 5931 45124 5987 45180
rect 5987 45124 5991 45180
rect 5927 45120 5991 45124
rect 6007 45180 6071 45184
rect 6007 45124 6011 45180
rect 6011 45124 6067 45180
rect 6067 45124 6071 45180
rect 6007 45120 6071 45124
rect 6087 45180 6151 45184
rect 6087 45124 6091 45180
rect 6091 45124 6147 45180
rect 6147 45124 6151 45180
rect 6087 45120 6151 45124
rect 9111 45180 9175 45184
rect 9111 45124 9115 45180
rect 9115 45124 9171 45180
rect 9171 45124 9175 45180
rect 9111 45120 9175 45124
rect 9191 45180 9255 45184
rect 9191 45124 9195 45180
rect 9195 45124 9251 45180
rect 9251 45124 9255 45180
rect 9191 45120 9255 45124
rect 9271 45180 9335 45184
rect 9271 45124 9275 45180
rect 9275 45124 9331 45180
rect 9331 45124 9335 45180
rect 9271 45120 9335 45124
rect 9351 45180 9415 45184
rect 9351 45124 9355 45180
rect 9355 45124 9411 45180
rect 9411 45124 9415 45180
rect 9351 45120 9415 45124
rect 7972 44780 8036 44844
rect 4215 44636 4279 44640
rect 4215 44580 4219 44636
rect 4219 44580 4275 44636
rect 4275 44580 4279 44636
rect 4215 44576 4279 44580
rect 4295 44636 4359 44640
rect 4295 44580 4299 44636
rect 4299 44580 4355 44636
rect 4355 44580 4359 44636
rect 4295 44576 4359 44580
rect 4375 44636 4439 44640
rect 4375 44580 4379 44636
rect 4379 44580 4435 44636
rect 4435 44580 4439 44636
rect 4375 44576 4439 44580
rect 4455 44636 4519 44640
rect 4455 44580 4459 44636
rect 4459 44580 4515 44636
rect 4515 44580 4519 44636
rect 4455 44576 4519 44580
rect 7479 44636 7543 44640
rect 7479 44580 7483 44636
rect 7483 44580 7539 44636
rect 7539 44580 7543 44636
rect 7479 44576 7543 44580
rect 7559 44636 7623 44640
rect 7559 44580 7563 44636
rect 7563 44580 7619 44636
rect 7619 44580 7623 44636
rect 7559 44576 7623 44580
rect 7639 44636 7703 44640
rect 7639 44580 7643 44636
rect 7643 44580 7699 44636
rect 7699 44580 7703 44636
rect 7639 44576 7703 44580
rect 7719 44636 7783 44640
rect 7719 44580 7723 44636
rect 7723 44580 7779 44636
rect 7779 44580 7783 44636
rect 7719 44576 7783 44580
rect 3556 44372 3620 44436
rect 11100 44372 11164 44436
rect 7236 44236 7300 44300
rect 2584 44092 2648 44096
rect 2584 44036 2588 44092
rect 2588 44036 2644 44092
rect 2644 44036 2648 44092
rect 2584 44032 2648 44036
rect 2664 44092 2728 44096
rect 2664 44036 2668 44092
rect 2668 44036 2724 44092
rect 2724 44036 2728 44092
rect 2664 44032 2728 44036
rect 2744 44092 2808 44096
rect 2744 44036 2748 44092
rect 2748 44036 2804 44092
rect 2804 44036 2808 44092
rect 2744 44032 2808 44036
rect 2824 44092 2888 44096
rect 2824 44036 2828 44092
rect 2828 44036 2884 44092
rect 2884 44036 2888 44092
rect 2824 44032 2888 44036
rect 5847 44092 5911 44096
rect 5847 44036 5851 44092
rect 5851 44036 5907 44092
rect 5907 44036 5911 44092
rect 5847 44032 5911 44036
rect 5927 44092 5991 44096
rect 5927 44036 5931 44092
rect 5931 44036 5987 44092
rect 5987 44036 5991 44092
rect 5927 44032 5991 44036
rect 6007 44092 6071 44096
rect 6007 44036 6011 44092
rect 6011 44036 6067 44092
rect 6067 44036 6071 44092
rect 6007 44032 6071 44036
rect 6087 44092 6151 44096
rect 6087 44036 6091 44092
rect 6091 44036 6147 44092
rect 6147 44036 6151 44092
rect 6087 44032 6151 44036
rect 9111 44092 9175 44096
rect 9111 44036 9115 44092
rect 9115 44036 9171 44092
rect 9171 44036 9175 44092
rect 9111 44032 9175 44036
rect 9191 44092 9255 44096
rect 9191 44036 9195 44092
rect 9195 44036 9251 44092
rect 9251 44036 9255 44092
rect 9191 44032 9255 44036
rect 9271 44092 9335 44096
rect 9271 44036 9275 44092
rect 9275 44036 9331 44092
rect 9331 44036 9335 44092
rect 9271 44032 9335 44036
rect 9351 44092 9415 44096
rect 9351 44036 9355 44092
rect 9355 44036 9411 44092
rect 9411 44036 9415 44092
rect 9351 44032 9415 44036
rect 4215 43548 4279 43552
rect 4215 43492 4219 43548
rect 4219 43492 4275 43548
rect 4275 43492 4279 43548
rect 4215 43488 4279 43492
rect 4295 43548 4359 43552
rect 4295 43492 4299 43548
rect 4299 43492 4355 43548
rect 4355 43492 4359 43548
rect 4295 43488 4359 43492
rect 4375 43548 4439 43552
rect 4375 43492 4379 43548
rect 4379 43492 4435 43548
rect 4435 43492 4439 43548
rect 4375 43488 4439 43492
rect 4455 43548 4519 43552
rect 4455 43492 4459 43548
rect 4459 43492 4515 43548
rect 4515 43492 4519 43548
rect 4455 43488 4519 43492
rect 7479 43548 7543 43552
rect 7479 43492 7483 43548
rect 7483 43492 7539 43548
rect 7539 43492 7543 43548
rect 7479 43488 7543 43492
rect 7559 43548 7623 43552
rect 7559 43492 7563 43548
rect 7563 43492 7619 43548
rect 7619 43492 7623 43548
rect 7559 43488 7623 43492
rect 7639 43548 7703 43552
rect 7639 43492 7643 43548
rect 7643 43492 7699 43548
rect 7699 43492 7703 43548
rect 7639 43488 7703 43492
rect 7719 43548 7783 43552
rect 7719 43492 7723 43548
rect 7723 43492 7779 43548
rect 7779 43492 7783 43548
rect 7719 43488 7783 43492
rect 11468 43480 11532 43484
rect 11468 43424 11482 43480
rect 11482 43424 11532 43480
rect 11468 43420 11532 43424
rect 8156 43012 8220 43076
rect 2584 43004 2648 43008
rect 2584 42948 2588 43004
rect 2588 42948 2644 43004
rect 2644 42948 2648 43004
rect 2584 42944 2648 42948
rect 2664 43004 2728 43008
rect 2664 42948 2668 43004
rect 2668 42948 2724 43004
rect 2724 42948 2728 43004
rect 2664 42944 2728 42948
rect 2744 43004 2808 43008
rect 2744 42948 2748 43004
rect 2748 42948 2804 43004
rect 2804 42948 2808 43004
rect 2744 42944 2808 42948
rect 2824 43004 2888 43008
rect 2824 42948 2828 43004
rect 2828 42948 2884 43004
rect 2884 42948 2888 43004
rect 2824 42944 2888 42948
rect 5847 43004 5911 43008
rect 5847 42948 5851 43004
rect 5851 42948 5907 43004
rect 5907 42948 5911 43004
rect 5847 42944 5911 42948
rect 5927 43004 5991 43008
rect 5927 42948 5931 43004
rect 5931 42948 5987 43004
rect 5987 42948 5991 43004
rect 5927 42944 5991 42948
rect 6007 43004 6071 43008
rect 6007 42948 6011 43004
rect 6011 42948 6067 43004
rect 6067 42948 6071 43004
rect 6007 42944 6071 42948
rect 6087 43004 6151 43008
rect 6087 42948 6091 43004
rect 6091 42948 6147 43004
rect 6147 42948 6151 43004
rect 6087 42944 6151 42948
rect 9111 43004 9175 43008
rect 9111 42948 9115 43004
rect 9115 42948 9171 43004
rect 9171 42948 9175 43004
rect 9111 42944 9175 42948
rect 9191 43004 9255 43008
rect 9191 42948 9195 43004
rect 9195 42948 9251 43004
rect 9251 42948 9255 43004
rect 9191 42944 9255 42948
rect 9271 43004 9335 43008
rect 9271 42948 9275 43004
rect 9275 42948 9331 43004
rect 9331 42948 9335 43004
rect 9271 42944 9335 42948
rect 9351 43004 9415 43008
rect 9351 42948 9355 43004
rect 9355 42948 9411 43004
rect 9411 42948 9415 43004
rect 9351 42944 9415 42948
rect 8340 42740 8404 42804
rect 10732 42604 10796 42668
rect 10548 42468 10612 42532
rect 4215 42460 4279 42464
rect 4215 42404 4219 42460
rect 4219 42404 4275 42460
rect 4275 42404 4279 42460
rect 4215 42400 4279 42404
rect 4295 42460 4359 42464
rect 4295 42404 4299 42460
rect 4299 42404 4355 42460
rect 4355 42404 4359 42460
rect 4295 42400 4359 42404
rect 4375 42460 4439 42464
rect 4375 42404 4379 42460
rect 4379 42404 4435 42460
rect 4435 42404 4439 42460
rect 4375 42400 4439 42404
rect 4455 42460 4519 42464
rect 4455 42404 4459 42460
rect 4459 42404 4515 42460
rect 4515 42404 4519 42460
rect 4455 42400 4519 42404
rect 7479 42460 7543 42464
rect 7479 42404 7483 42460
rect 7483 42404 7539 42460
rect 7539 42404 7543 42460
rect 7479 42400 7543 42404
rect 7559 42460 7623 42464
rect 7559 42404 7563 42460
rect 7563 42404 7619 42460
rect 7619 42404 7623 42460
rect 7559 42400 7623 42404
rect 7639 42460 7703 42464
rect 7639 42404 7643 42460
rect 7643 42404 7699 42460
rect 7699 42404 7703 42460
rect 7639 42400 7703 42404
rect 7719 42460 7783 42464
rect 7719 42404 7723 42460
rect 7723 42404 7779 42460
rect 7779 42404 7783 42460
rect 7719 42400 7783 42404
rect 10364 42332 10428 42396
rect 10916 42060 10980 42124
rect 2584 41916 2648 41920
rect 2584 41860 2588 41916
rect 2588 41860 2644 41916
rect 2644 41860 2648 41916
rect 2584 41856 2648 41860
rect 2664 41916 2728 41920
rect 2664 41860 2668 41916
rect 2668 41860 2724 41916
rect 2724 41860 2728 41916
rect 2664 41856 2728 41860
rect 2744 41916 2808 41920
rect 2744 41860 2748 41916
rect 2748 41860 2804 41916
rect 2804 41860 2808 41916
rect 2744 41856 2808 41860
rect 2824 41916 2888 41920
rect 2824 41860 2828 41916
rect 2828 41860 2884 41916
rect 2884 41860 2888 41916
rect 2824 41856 2888 41860
rect 5847 41916 5911 41920
rect 5847 41860 5851 41916
rect 5851 41860 5907 41916
rect 5907 41860 5911 41916
rect 5847 41856 5911 41860
rect 5927 41916 5991 41920
rect 5927 41860 5931 41916
rect 5931 41860 5987 41916
rect 5987 41860 5991 41916
rect 5927 41856 5991 41860
rect 6007 41916 6071 41920
rect 6007 41860 6011 41916
rect 6011 41860 6067 41916
rect 6067 41860 6071 41916
rect 6007 41856 6071 41860
rect 6087 41916 6151 41920
rect 6087 41860 6091 41916
rect 6091 41860 6147 41916
rect 6147 41860 6151 41916
rect 6087 41856 6151 41860
rect 9111 41916 9175 41920
rect 9111 41860 9115 41916
rect 9115 41860 9171 41916
rect 9171 41860 9175 41916
rect 9111 41856 9175 41860
rect 9191 41916 9255 41920
rect 9191 41860 9195 41916
rect 9195 41860 9251 41916
rect 9251 41860 9255 41916
rect 9191 41856 9255 41860
rect 9271 41916 9335 41920
rect 9271 41860 9275 41916
rect 9275 41860 9331 41916
rect 9331 41860 9335 41916
rect 9271 41856 9335 41860
rect 9351 41916 9415 41920
rect 9351 41860 9355 41916
rect 9355 41860 9411 41916
rect 9411 41860 9415 41916
rect 9351 41856 9415 41860
rect 8156 41516 8220 41580
rect 4215 41372 4279 41376
rect 4215 41316 4219 41372
rect 4219 41316 4275 41372
rect 4275 41316 4279 41372
rect 4215 41312 4279 41316
rect 4295 41372 4359 41376
rect 4295 41316 4299 41372
rect 4299 41316 4355 41372
rect 4355 41316 4359 41372
rect 4295 41312 4359 41316
rect 4375 41372 4439 41376
rect 4375 41316 4379 41372
rect 4379 41316 4435 41372
rect 4435 41316 4439 41372
rect 4375 41312 4439 41316
rect 4455 41372 4519 41376
rect 4455 41316 4459 41372
rect 4459 41316 4515 41372
rect 4515 41316 4519 41372
rect 4455 41312 4519 41316
rect 7479 41372 7543 41376
rect 7479 41316 7483 41372
rect 7483 41316 7539 41372
rect 7539 41316 7543 41372
rect 7479 41312 7543 41316
rect 7559 41372 7623 41376
rect 7559 41316 7563 41372
rect 7563 41316 7619 41372
rect 7619 41316 7623 41372
rect 7559 41312 7623 41316
rect 7639 41372 7703 41376
rect 7639 41316 7643 41372
rect 7643 41316 7699 41372
rect 7699 41316 7703 41372
rect 7639 41312 7703 41316
rect 7719 41372 7783 41376
rect 7719 41316 7723 41372
rect 7723 41316 7779 41372
rect 7779 41316 7783 41372
rect 7719 41312 7783 41316
rect 8156 41244 8220 41308
rect 2584 40828 2648 40832
rect 2584 40772 2588 40828
rect 2588 40772 2644 40828
rect 2644 40772 2648 40828
rect 2584 40768 2648 40772
rect 2664 40828 2728 40832
rect 2664 40772 2668 40828
rect 2668 40772 2724 40828
rect 2724 40772 2728 40828
rect 2664 40768 2728 40772
rect 2744 40828 2808 40832
rect 2744 40772 2748 40828
rect 2748 40772 2804 40828
rect 2804 40772 2808 40828
rect 2744 40768 2808 40772
rect 2824 40828 2888 40832
rect 2824 40772 2828 40828
rect 2828 40772 2884 40828
rect 2884 40772 2888 40828
rect 2824 40768 2888 40772
rect 5847 40828 5911 40832
rect 5847 40772 5851 40828
rect 5851 40772 5907 40828
rect 5907 40772 5911 40828
rect 5847 40768 5911 40772
rect 5927 40828 5991 40832
rect 5927 40772 5931 40828
rect 5931 40772 5987 40828
rect 5987 40772 5991 40828
rect 5927 40768 5991 40772
rect 6007 40828 6071 40832
rect 6007 40772 6011 40828
rect 6011 40772 6067 40828
rect 6067 40772 6071 40828
rect 6007 40768 6071 40772
rect 6087 40828 6151 40832
rect 6087 40772 6091 40828
rect 6091 40772 6147 40828
rect 6147 40772 6151 40828
rect 6087 40768 6151 40772
rect 9111 40828 9175 40832
rect 9111 40772 9115 40828
rect 9115 40772 9171 40828
rect 9171 40772 9175 40828
rect 9111 40768 9175 40772
rect 9191 40828 9255 40832
rect 9191 40772 9195 40828
rect 9195 40772 9251 40828
rect 9251 40772 9255 40828
rect 9191 40768 9255 40772
rect 9271 40828 9335 40832
rect 9271 40772 9275 40828
rect 9275 40772 9331 40828
rect 9331 40772 9335 40828
rect 9271 40768 9335 40772
rect 9351 40828 9415 40832
rect 9351 40772 9355 40828
rect 9355 40772 9411 40828
rect 9411 40772 9415 40828
rect 9351 40768 9415 40772
rect 8524 40760 8588 40764
rect 8524 40704 8574 40760
rect 8574 40704 8588 40760
rect 8524 40700 8588 40704
rect 7972 40428 8036 40492
rect 10180 40488 10244 40492
rect 10180 40432 10194 40488
rect 10194 40432 10244 40488
rect 10180 40428 10244 40432
rect 4215 40284 4279 40288
rect 4215 40228 4219 40284
rect 4219 40228 4275 40284
rect 4275 40228 4279 40284
rect 4215 40224 4279 40228
rect 4295 40284 4359 40288
rect 4295 40228 4299 40284
rect 4299 40228 4355 40284
rect 4355 40228 4359 40284
rect 4295 40224 4359 40228
rect 4375 40284 4439 40288
rect 4375 40228 4379 40284
rect 4379 40228 4435 40284
rect 4435 40228 4439 40284
rect 4375 40224 4439 40228
rect 4455 40284 4519 40288
rect 4455 40228 4459 40284
rect 4459 40228 4515 40284
rect 4515 40228 4519 40284
rect 4455 40224 4519 40228
rect 7479 40284 7543 40288
rect 7479 40228 7483 40284
rect 7483 40228 7539 40284
rect 7539 40228 7543 40284
rect 7479 40224 7543 40228
rect 7559 40284 7623 40288
rect 7559 40228 7563 40284
rect 7563 40228 7619 40284
rect 7619 40228 7623 40284
rect 7559 40224 7623 40228
rect 7639 40284 7703 40288
rect 7639 40228 7643 40284
rect 7643 40228 7699 40284
rect 7699 40228 7703 40284
rect 7639 40224 7703 40228
rect 7719 40284 7783 40288
rect 7719 40228 7723 40284
rect 7723 40228 7779 40284
rect 7779 40228 7783 40284
rect 7719 40224 7783 40228
rect 10548 40156 10612 40220
rect 2584 39740 2648 39744
rect 2584 39684 2588 39740
rect 2588 39684 2644 39740
rect 2644 39684 2648 39740
rect 2584 39680 2648 39684
rect 2664 39740 2728 39744
rect 2664 39684 2668 39740
rect 2668 39684 2724 39740
rect 2724 39684 2728 39740
rect 2664 39680 2728 39684
rect 2744 39740 2808 39744
rect 2744 39684 2748 39740
rect 2748 39684 2804 39740
rect 2804 39684 2808 39740
rect 2744 39680 2808 39684
rect 2824 39740 2888 39744
rect 2824 39684 2828 39740
rect 2828 39684 2884 39740
rect 2884 39684 2888 39740
rect 2824 39680 2888 39684
rect 5847 39740 5911 39744
rect 5847 39684 5851 39740
rect 5851 39684 5907 39740
rect 5907 39684 5911 39740
rect 5847 39680 5911 39684
rect 5927 39740 5991 39744
rect 5927 39684 5931 39740
rect 5931 39684 5987 39740
rect 5987 39684 5991 39740
rect 5927 39680 5991 39684
rect 6007 39740 6071 39744
rect 6007 39684 6011 39740
rect 6011 39684 6067 39740
rect 6067 39684 6071 39740
rect 6007 39680 6071 39684
rect 6087 39740 6151 39744
rect 6087 39684 6091 39740
rect 6091 39684 6147 39740
rect 6147 39684 6151 39740
rect 6087 39680 6151 39684
rect 9111 39740 9175 39744
rect 9111 39684 9115 39740
rect 9115 39684 9171 39740
rect 9171 39684 9175 39740
rect 9111 39680 9175 39684
rect 9191 39740 9255 39744
rect 9191 39684 9195 39740
rect 9195 39684 9251 39740
rect 9251 39684 9255 39740
rect 9191 39680 9255 39684
rect 9271 39740 9335 39744
rect 9271 39684 9275 39740
rect 9275 39684 9331 39740
rect 9331 39684 9335 39740
rect 9271 39680 9335 39684
rect 9351 39740 9415 39744
rect 9351 39684 9355 39740
rect 9355 39684 9411 39740
rect 9411 39684 9415 39740
rect 9351 39680 9415 39684
rect 10364 39612 10428 39676
rect 10916 39612 10980 39676
rect 8524 39476 8588 39540
rect 4215 39196 4279 39200
rect 4215 39140 4219 39196
rect 4219 39140 4275 39196
rect 4275 39140 4279 39196
rect 4215 39136 4279 39140
rect 4295 39196 4359 39200
rect 4295 39140 4299 39196
rect 4299 39140 4355 39196
rect 4355 39140 4359 39196
rect 4295 39136 4359 39140
rect 4375 39196 4439 39200
rect 4375 39140 4379 39196
rect 4379 39140 4435 39196
rect 4435 39140 4439 39196
rect 4375 39136 4439 39140
rect 4455 39196 4519 39200
rect 4455 39140 4459 39196
rect 4459 39140 4515 39196
rect 4515 39140 4519 39196
rect 4455 39136 4519 39140
rect 7479 39196 7543 39200
rect 7479 39140 7483 39196
rect 7483 39140 7539 39196
rect 7539 39140 7543 39196
rect 7479 39136 7543 39140
rect 7559 39196 7623 39200
rect 7559 39140 7563 39196
rect 7563 39140 7619 39196
rect 7619 39140 7623 39196
rect 7559 39136 7623 39140
rect 7639 39196 7703 39200
rect 7639 39140 7643 39196
rect 7643 39140 7699 39196
rect 7699 39140 7703 39196
rect 7639 39136 7703 39140
rect 7719 39196 7783 39200
rect 7719 39140 7723 39196
rect 7723 39140 7779 39196
rect 7779 39140 7783 39196
rect 7719 39136 7783 39140
rect 8892 38796 8956 38860
rect 11468 38660 11532 38724
rect 2584 38652 2648 38656
rect 2584 38596 2588 38652
rect 2588 38596 2644 38652
rect 2644 38596 2648 38652
rect 2584 38592 2648 38596
rect 2664 38652 2728 38656
rect 2664 38596 2668 38652
rect 2668 38596 2724 38652
rect 2724 38596 2728 38652
rect 2664 38592 2728 38596
rect 2744 38652 2808 38656
rect 2744 38596 2748 38652
rect 2748 38596 2804 38652
rect 2804 38596 2808 38652
rect 2744 38592 2808 38596
rect 2824 38652 2888 38656
rect 2824 38596 2828 38652
rect 2828 38596 2884 38652
rect 2884 38596 2888 38652
rect 2824 38592 2888 38596
rect 5847 38652 5911 38656
rect 5847 38596 5851 38652
rect 5851 38596 5907 38652
rect 5907 38596 5911 38652
rect 5847 38592 5911 38596
rect 5927 38652 5991 38656
rect 5927 38596 5931 38652
rect 5931 38596 5987 38652
rect 5987 38596 5991 38652
rect 5927 38592 5991 38596
rect 6007 38652 6071 38656
rect 6007 38596 6011 38652
rect 6011 38596 6067 38652
rect 6067 38596 6071 38652
rect 6007 38592 6071 38596
rect 6087 38652 6151 38656
rect 6087 38596 6091 38652
rect 6091 38596 6147 38652
rect 6147 38596 6151 38652
rect 6087 38592 6151 38596
rect 9111 38652 9175 38656
rect 9111 38596 9115 38652
rect 9115 38596 9171 38652
rect 9171 38596 9175 38652
rect 9111 38592 9175 38596
rect 9191 38652 9255 38656
rect 9191 38596 9195 38652
rect 9195 38596 9251 38652
rect 9251 38596 9255 38652
rect 9191 38592 9255 38596
rect 9271 38652 9335 38656
rect 9271 38596 9275 38652
rect 9275 38596 9331 38652
rect 9331 38596 9335 38652
rect 9271 38592 9335 38596
rect 9351 38652 9415 38656
rect 9351 38596 9355 38652
rect 9355 38596 9411 38652
rect 9411 38596 9415 38652
rect 9351 38592 9415 38596
rect 9812 38584 9876 38588
rect 9812 38528 9826 38584
rect 9826 38528 9876 38584
rect 9812 38524 9876 38528
rect 8340 38252 8404 38316
rect 8524 38252 8588 38316
rect 8892 38116 8956 38180
rect 4215 38108 4279 38112
rect 4215 38052 4219 38108
rect 4219 38052 4275 38108
rect 4275 38052 4279 38108
rect 4215 38048 4279 38052
rect 4295 38108 4359 38112
rect 4295 38052 4299 38108
rect 4299 38052 4355 38108
rect 4355 38052 4359 38108
rect 4295 38048 4359 38052
rect 4375 38108 4439 38112
rect 4375 38052 4379 38108
rect 4379 38052 4435 38108
rect 4435 38052 4439 38108
rect 4375 38048 4439 38052
rect 4455 38108 4519 38112
rect 4455 38052 4459 38108
rect 4459 38052 4515 38108
rect 4515 38052 4519 38108
rect 4455 38048 4519 38052
rect 7479 38108 7543 38112
rect 7479 38052 7483 38108
rect 7483 38052 7539 38108
rect 7539 38052 7543 38108
rect 7479 38048 7543 38052
rect 7559 38108 7623 38112
rect 7559 38052 7563 38108
rect 7563 38052 7619 38108
rect 7619 38052 7623 38108
rect 7559 38048 7623 38052
rect 7639 38108 7703 38112
rect 7639 38052 7643 38108
rect 7643 38052 7699 38108
rect 7699 38052 7703 38108
rect 7639 38048 7703 38052
rect 7719 38108 7783 38112
rect 7719 38052 7723 38108
rect 7723 38052 7779 38108
rect 7779 38052 7783 38108
rect 7719 38048 7783 38052
rect 8524 37844 8588 37908
rect 9628 37708 9692 37772
rect 2584 37564 2648 37568
rect 2584 37508 2588 37564
rect 2588 37508 2644 37564
rect 2644 37508 2648 37564
rect 2584 37504 2648 37508
rect 2664 37564 2728 37568
rect 2664 37508 2668 37564
rect 2668 37508 2724 37564
rect 2724 37508 2728 37564
rect 2664 37504 2728 37508
rect 2744 37564 2808 37568
rect 2744 37508 2748 37564
rect 2748 37508 2804 37564
rect 2804 37508 2808 37564
rect 2744 37504 2808 37508
rect 2824 37564 2888 37568
rect 2824 37508 2828 37564
rect 2828 37508 2884 37564
rect 2884 37508 2888 37564
rect 2824 37504 2888 37508
rect 5847 37564 5911 37568
rect 5847 37508 5851 37564
rect 5851 37508 5907 37564
rect 5907 37508 5911 37564
rect 5847 37504 5911 37508
rect 5927 37564 5991 37568
rect 5927 37508 5931 37564
rect 5931 37508 5987 37564
rect 5987 37508 5991 37564
rect 5927 37504 5991 37508
rect 6007 37564 6071 37568
rect 6007 37508 6011 37564
rect 6011 37508 6067 37564
rect 6067 37508 6071 37564
rect 6007 37504 6071 37508
rect 6087 37564 6151 37568
rect 6087 37508 6091 37564
rect 6091 37508 6147 37564
rect 6147 37508 6151 37564
rect 6087 37504 6151 37508
rect 9111 37564 9175 37568
rect 9111 37508 9115 37564
rect 9115 37508 9171 37564
rect 9171 37508 9175 37564
rect 9111 37504 9175 37508
rect 9191 37564 9255 37568
rect 9191 37508 9195 37564
rect 9195 37508 9251 37564
rect 9251 37508 9255 37564
rect 9191 37504 9255 37508
rect 9271 37564 9335 37568
rect 9271 37508 9275 37564
rect 9275 37508 9331 37564
rect 9331 37508 9335 37564
rect 9271 37504 9335 37508
rect 9351 37564 9415 37568
rect 9351 37508 9355 37564
rect 9355 37508 9411 37564
rect 9411 37508 9415 37564
rect 9351 37504 9415 37508
rect 3372 37164 3436 37228
rect 4215 37020 4279 37024
rect 4215 36964 4219 37020
rect 4219 36964 4275 37020
rect 4275 36964 4279 37020
rect 4215 36960 4279 36964
rect 4295 37020 4359 37024
rect 4295 36964 4299 37020
rect 4299 36964 4355 37020
rect 4355 36964 4359 37020
rect 4295 36960 4359 36964
rect 4375 37020 4439 37024
rect 4375 36964 4379 37020
rect 4379 36964 4435 37020
rect 4435 36964 4439 37020
rect 4375 36960 4439 36964
rect 4455 37020 4519 37024
rect 4455 36964 4459 37020
rect 4459 36964 4515 37020
rect 4515 36964 4519 37020
rect 4455 36960 4519 36964
rect 7479 37020 7543 37024
rect 7479 36964 7483 37020
rect 7483 36964 7539 37020
rect 7539 36964 7543 37020
rect 7479 36960 7543 36964
rect 7559 37020 7623 37024
rect 7559 36964 7563 37020
rect 7563 36964 7619 37020
rect 7619 36964 7623 37020
rect 7559 36960 7623 36964
rect 7639 37020 7703 37024
rect 7639 36964 7643 37020
rect 7643 36964 7699 37020
rect 7699 36964 7703 37020
rect 7639 36960 7703 36964
rect 7719 37020 7783 37024
rect 7719 36964 7723 37020
rect 7723 36964 7779 37020
rect 7779 36964 7783 37020
rect 7719 36960 7783 36964
rect 10548 36816 10612 36820
rect 10548 36760 10598 36816
rect 10598 36760 10612 36816
rect 10548 36756 10612 36760
rect 11652 36816 11716 36820
rect 11652 36760 11666 36816
rect 11666 36760 11716 36816
rect 11652 36756 11716 36760
rect 10180 36620 10244 36684
rect 2584 36476 2648 36480
rect 2584 36420 2588 36476
rect 2588 36420 2644 36476
rect 2644 36420 2648 36476
rect 2584 36416 2648 36420
rect 2664 36476 2728 36480
rect 2664 36420 2668 36476
rect 2668 36420 2724 36476
rect 2724 36420 2728 36476
rect 2664 36416 2728 36420
rect 2744 36476 2808 36480
rect 2744 36420 2748 36476
rect 2748 36420 2804 36476
rect 2804 36420 2808 36476
rect 2744 36416 2808 36420
rect 2824 36476 2888 36480
rect 2824 36420 2828 36476
rect 2828 36420 2884 36476
rect 2884 36420 2888 36476
rect 2824 36416 2888 36420
rect 5847 36476 5911 36480
rect 5847 36420 5851 36476
rect 5851 36420 5907 36476
rect 5907 36420 5911 36476
rect 5847 36416 5911 36420
rect 5927 36476 5991 36480
rect 5927 36420 5931 36476
rect 5931 36420 5987 36476
rect 5987 36420 5991 36476
rect 5927 36416 5991 36420
rect 6007 36476 6071 36480
rect 6007 36420 6011 36476
rect 6011 36420 6067 36476
rect 6067 36420 6071 36476
rect 6007 36416 6071 36420
rect 6087 36476 6151 36480
rect 6087 36420 6091 36476
rect 6091 36420 6147 36476
rect 6147 36420 6151 36476
rect 6087 36416 6151 36420
rect 9111 36476 9175 36480
rect 9111 36420 9115 36476
rect 9115 36420 9171 36476
rect 9171 36420 9175 36476
rect 9111 36416 9175 36420
rect 9191 36476 9255 36480
rect 9191 36420 9195 36476
rect 9195 36420 9251 36476
rect 9251 36420 9255 36476
rect 9191 36416 9255 36420
rect 9271 36476 9335 36480
rect 9271 36420 9275 36476
rect 9275 36420 9331 36476
rect 9331 36420 9335 36476
rect 9271 36416 9335 36420
rect 9351 36476 9415 36480
rect 9351 36420 9355 36476
rect 9355 36420 9411 36476
rect 9411 36420 9415 36476
rect 9351 36416 9415 36420
rect 8340 36212 8404 36276
rect 8892 36000 8956 36004
rect 8892 35944 8906 36000
rect 8906 35944 8956 36000
rect 8892 35940 8956 35944
rect 4215 35932 4279 35936
rect 4215 35876 4219 35932
rect 4219 35876 4275 35932
rect 4275 35876 4279 35932
rect 4215 35872 4279 35876
rect 4295 35932 4359 35936
rect 4295 35876 4299 35932
rect 4299 35876 4355 35932
rect 4355 35876 4359 35932
rect 4295 35872 4359 35876
rect 4375 35932 4439 35936
rect 4375 35876 4379 35932
rect 4379 35876 4435 35932
rect 4435 35876 4439 35932
rect 4375 35872 4439 35876
rect 4455 35932 4519 35936
rect 4455 35876 4459 35932
rect 4459 35876 4515 35932
rect 4515 35876 4519 35932
rect 4455 35872 4519 35876
rect 7479 35932 7543 35936
rect 7479 35876 7483 35932
rect 7483 35876 7539 35932
rect 7539 35876 7543 35932
rect 7479 35872 7543 35876
rect 7559 35932 7623 35936
rect 7559 35876 7563 35932
rect 7563 35876 7619 35932
rect 7619 35876 7623 35932
rect 7559 35872 7623 35876
rect 7639 35932 7703 35936
rect 7639 35876 7643 35932
rect 7643 35876 7699 35932
rect 7699 35876 7703 35932
rect 7639 35872 7703 35876
rect 7719 35932 7783 35936
rect 7719 35876 7723 35932
rect 7723 35876 7779 35932
rect 7779 35876 7783 35932
rect 7719 35872 7783 35876
rect 2584 35388 2648 35392
rect 2584 35332 2588 35388
rect 2588 35332 2644 35388
rect 2644 35332 2648 35388
rect 2584 35328 2648 35332
rect 2664 35388 2728 35392
rect 2664 35332 2668 35388
rect 2668 35332 2724 35388
rect 2724 35332 2728 35388
rect 2664 35328 2728 35332
rect 2744 35388 2808 35392
rect 2744 35332 2748 35388
rect 2748 35332 2804 35388
rect 2804 35332 2808 35388
rect 2744 35328 2808 35332
rect 2824 35388 2888 35392
rect 2824 35332 2828 35388
rect 2828 35332 2884 35388
rect 2884 35332 2888 35388
rect 2824 35328 2888 35332
rect 5847 35388 5911 35392
rect 5847 35332 5851 35388
rect 5851 35332 5907 35388
rect 5907 35332 5911 35388
rect 5847 35328 5911 35332
rect 5927 35388 5991 35392
rect 5927 35332 5931 35388
rect 5931 35332 5987 35388
rect 5987 35332 5991 35388
rect 5927 35328 5991 35332
rect 6007 35388 6071 35392
rect 6007 35332 6011 35388
rect 6011 35332 6067 35388
rect 6067 35332 6071 35388
rect 6007 35328 6071 35332
rect 6087 35388 6151 35392
rect 6087 35332 6091 35388
rect 6091 35332 6147 35388
rect 6147 35332 6151 35388
rect 6087 35328 6151 35332
rect 9111 35388 9175 35392
rect 9111 35332 9115 35388
rect 9115 35332 9171 35388
rect 9171 35332 9175 35388
rect 9111 35328 9175 35332
rect 9191 35388 9255 35392
rect 9191 35332 9195 35388
rect 9195 35332 9251 35388
rect 9251 35332 9255 35388
rect 9191 35328 9255 35332
rect 9271 35388 9335 35392
rect 9271 35332 9275 35388
rect 9275 35332 9331 35388
rect 9331 35332 9335 35388
rect 9271 35328 9335 35332
rect 9351 35388 9415 35392
rect 9351 35332 9355 35388
rect 9355 35332 9411 35388
rect 9411 35332 9415 35388
rect 9351 35328 9415 35332
rect 4215 34844 4279 34848
rect 4215 34788 4219 34844
rect 4219 34788 4275 34844
rect 4275 34788 4279 34844
rect 4215 34784 4279 34788
rect 4295 34844 4359 34848
rect 4295 34788 4299 34844
rect 4299 34788 4355 34844
rect 4355 34788 4359 34844
rect 4295 34784 4359 34788
rect 4375 34844 4439 34848
rect 4375 34788 4379 34844
rect 4379 34788 4435 34844
rect 4435 34788 4439 34844
rect 4375 34784 4439 34788
rect 4455 34844 4519 34848
rect 4455 34788 4459 34844
rect 4459 34788 4515 34844
rect 4515 34788 4519 34844
rect 4455 34784 4519 34788
rect 7479 34844 7543 34848
rect 7479 34788 7483 34844
rect 7483 34788 7539 34844
rect 7539 34788 7543 34844
rect 7479 34784 7543 34788
rect 7559 34844 7623 34848
rect 7559 34788 7563 34844
rect 7563 34788 7619 34844
rect 7619 34788 7623 34844
rect 7559 34784 7623 34788
rect 7639 34844 7703 34848
rect 7639 34788 7643 34844
rect 7643 34788 7699 34844
rect 7699 34788 7703 34844
rect 7639 34784 7703 34788
rect 7719 34844 7783 34848
rect 7719 34788 7723 34844
rect 7723 34788 7779 34844
rect 7779 34788 7783 34844
rect 7719 34784 7783 34788
rect 8708 34504 8772 34508
rect 8708 34448 8722 34504
rect 8722 34448 8772 34504
rect 8708 34444 8772 34448
rect 2584 34300 2648 34304
rect 2584 34244 2588 34300
rect 2588 34244 2644 34300
rect 2644 34244 2648 34300
rect 2584 34240 2648 34244
rect 2664 34300 2728 34304
rect 2664 34244 2668 34300
rect 2668 34244 2724 34300
rect 2724 34244 2728 34300
rect 2664 34240 2728 34244
rect 2744 34300 2808 34304
rect 2744 34244 2748 34300
rect 2748 34244 2804 34300
rect 2804 34244 2808 34300
rect 2744 34240 2808 34244
rect 2824 34300 2888 34304
rect 2824 34244 2828 34300
rect 2828 34244 2884 34300
rect 2884 34244 2888 34300
rect 2824 34240 2888 34244
rect 5847 34300 5911 34304
rect 5847 34244 5851 34300
rect 5851 34244 5907 34300
rect 5907 34244 5911 34300
rect 5847 34240 5911 34244
rect 5927 34300 5991 34304
rect 5927 34244 5931 34300
rect 5931 34244 5987 34300
rect 5987 34244 5991 34300
rect 5927 34240 5991 34244
rect 6007 34300 6071 34304
rect 6007 34244 6011 34300
rect 6011 34244 6067 34300
rect 6067 34244 6071 34300
rect 6007 34240 6071 34244
rect 6087 34300 6151 34304
rect 6087 34244 6091 34300
rect 6091 34244 6147 34300
rect 6147 34244 6151 34300
rect 6087 34240 6151 34244
rect 9111 34300 9175 34304
rect 9111 34244 9115 34300
rect 9115 34244 9171 34300
rect 9171 34244 9175 34300
rect 9111 34240 9175 34244
rect 9191 34300 9255 34304
rect 9191 34244 9195 34300
rect 9195 34244 9251 34300
rect 9251 34244 9255 34300
rect 9191 34240 9255 34244
rect 9271 34300 9335 34304
rect 9271 34244 9275 34300
rect 9275 34244 9331 34300
rect 9331 34244 9335 34300
rect 9271 34240 9335 34244
rect 9351 34300 9415 34304
rect 9351 34244 9355 34300
rect 9355 34244 9411 34300
rect 9411 34244 9415 34300
rect 9351 34240 9415 34244
rect 4215 33756 4279 33760
rect 4215 33700 4219 33756
rect 4219 33700 4275 33756
rect 4275 33700 4279 33756
rect 4215 33696 4279 33700
rect 4295 33756 4359 33760
rect 4295 33700 4299 33756
rect 4299 33700 4355 33756
rect 4355 33700 4359 33756
rect 4295 33696 4359 33700
rect 4375 33756 4439 33760
rect 4375 33700 4379 33756
rect 4379 33700 4435 33756
rect 4435 33700 4439 33756
rect 4375 33696 4439 33700
rect 4455 33756 4519 33760
rect 4455 33700 4459 33756
rect 4459 33700 4515 33756
rect 4515 33700 4519 33756
rect 4455 33696 4519 33700
rect 7479 33756 7543 33760
rect 7479 33700 7483 33756
rect 7483 33700 7539 33756
rect 7539 33700 7543 33756
rect 7479 33696 7543 33700
rect 7559 33756 7623 33760
rect 7559 33700 7563 33756
rect 7563 33700 7619 33756
rect 7619 33700 7623 33756
rect 7559 33696 7623 33700
rect 7639 33756 7703 33760
rect 7639 33700 7643 33756
rect 7643 33700 7699 33756
rect 7699 33700 7703 33756
rect 7639 33696 7703 33700
rect 7719 33756 7783 33760
rect 7719 33700 7723 33756
rect 7723 33700 7779 33756
rect 7779 33700 7783 33756
rect 7719 33696 7783 33700
rect 8524 33492 8588 33556
rect 10548 33356 10612 33420
rect 2584 33212 2648 33216
rect 2584 33156 2588 33212
rect 2588 33156 2644 33212
rect 2644 33156 2648 33212
rect 2584 33152 2648 33156
rect 2664 33212 2728 33216
rect 2664 33156 2668 33212
rect 2668 33156 2724 33212
rect 2724 33156 2728 33212
rect 2664 33152 2728 33156
rect 2744 33212 2808 33216
rect 2744 33156 2748 33212
rect 2748 33156 2804 33212
rect 2804 33156 2808 33212
rect 2744 33152 2808 33156
rect 2824 33212 2888 33216
rect 2824 33156 2828 33212
rect 2828 33156 2884 33212
rect 2884 33156 2888 33212
rect 2824 33152 2888 33156
rect 5847 33212 5911 33216
rect 5847 33156 5851 33212
rect 5851 33156 5907 33212
rect 5907 33156 5911 33212
rect 5847 33152 5911 33156
rect 5927 33212 5991 33216
rect 5927 33156 5931 33212
rect 5931 33156 5987 33212
rect 5987 33156 5991 33212
rect 5927 33152 5991 33156
rect 6007 33212 6071 33216
rect 6007 33156 6011 33212
rect 6011 33156 6067 33212
rect 6067 33156 6071 33212
rect 6007 33152 6071 33156
rect 6087 33212 6151 33216
rect 6087 33156 6091 33212
rect 6091 33156 6147 33212
rect 6147 33156 6151 33212
rect 6087 33152 6151 33156
rect 9111 33212 9175 33216
rect 9111 33156 9115 33212
rect 9115 33156 9171 33212
rect 9171 33156 9175 33212
rect 9111 33152 9175 33156
rect 9191 33212 9255 33216
rect 9191 33156 9195 33212
rect 9195 33156 9251 33212
rect 9251 33156 9255 33212
rect 9191 33152 9255 33156
rect 9271 33212 9335 33216
rect 9271 33156 9275 33212
rect 9275 33156 9331 33212
rect 9331 33156 9335 33212
rect 9271 33152 9335 33156
rect 9351 33212 9415 33216
rect 9351 33156 9355 33212
rect 9355 33156 9411 33212
rect 9411 33156 9415 33212
rect 9351 33152 9415 33156
rect 10548 33144 10612 33148
rect 10548 33088 10598 33144
rect 10598 33088 10612 33144
rect 10548 33084 10612 33088
rect 4215 32668 4279 32672
rect 4215 32612 4219 32668
rect 4219 32612 4275 32668
rect 4275 32612 4279 32668
rect 4215 32608 4279 32612
rect 4295 32668 4359 32672
rect 4295 32612 4299 32668
rect 4299 32612 4355 32668
rect 4355 32612 4359 32668
rect 4295 32608 4359 32612
rect 4375 32668 4439 32672
rect 4375 32612 4379 32668
rect 4379 32612 4435 32668
rect 4435 32612 4439 32668
rect 4375 32608 4439 32612
rect 4455 32668 4519 32672
rect 4455 32612 4459 32668
rect 4459 32612 4515 32668
rect 4515 32612 4519 32668
rect 4455 32608 4519 32612
rect 7479 32668 7543 32672
rect 7479 32612 7483 32668
rect 7483 32612 7539 32668
rect 7539 32612 7543 32668
rect 7479 32608 7543 32612
rect 7559 32668 7623 32672
rect 7559 32612 7563 32668
rect 7563 32612 7619 32668
rect 7619 32612 7623 32668
rect 7559 32608 7623 32612
rect 7639 32668 7703 32672
rect 7639 32612 7643 32668
rect 7643 32612 7699 32668
rect 7699 32612 7703 32668
rect 7639 32608 7703 32612
rect 7719 32668 7783 32672
rect 7719 32612 7723 32668
rect 7723 32612 7779 32668
rect 7779 32612 7783 32668
rect 7719 32608 7783 32612
rect 10732 32540 10796 32604
rect 2584 32124 2648 32128
rect 2584 32068 2588 32124
rect 2588 32068 2644 32124
rect 2644 32068 2648 32124
rect 2584 32064 2648 32068
rect 2664 32124 2728 32128
rect 2664 32068 2668 32124
rect 2668 32068 2724 32124
rect 2724 32068 2728 32124
rect 2664 32064 2728 32068
rect 2744 32124 2808 32128
rect 2744 32068 2748 32124
rect 2748 32068 2804 32124
rect 2804 32068 2808 32124
rect 2744 32064 2808 32068
rect 2824 32124 2888 32128
rect 2824 32068 2828 32124
rect 2828 32068 2884 32124
rect 2884 32068 2888 32124
rect 2824 32064 2888 32068
rect 5847 32124 5911 32128
rect 5847 32068 5851 32124
rect 5851 32068 5907 32124
rect 5907 32068 5911 32124
rect 5847 32064 5911 32068
rect 5927 32124 5991 32128
rect 5927 32068 5931 32124
rect 5931 32068 5987 32124
rect 5987 32068 5991 32124
rect 5927 32064 5991 32068
rect 6007 32124 6071 32128
rect 6007 32068 6011 32124
rect 6011 32068 6067 32124
rect 6067 32068 6071 32124
rect 6007 32064 6071 32068
rect 6087 32124 6151 32128
rect 6087 32068 6091 32124
rect 6091 32068 6147 32124
rect 6147 32068 6151 32124
rect 6087 32064 6151 32068
rect 9111 32124 9175 32128
rect 9111 32068 9115 32124
rect 9115 32068 9171 32124
rect 9171 32068 9175 32124
rect 9111 32064 9175 32068
rect 9191 32124 9255 32128
rect 9191 32068 9195 32124
rect 9195 32068 9251 32124
rect 9251 32068 9255 32124
rect 9191 32064 9255 32068
rect 9271 32124 9335 32128
rect 9271 32068 9275 32124
rect 9275 32068 9331 32124
rect 9331 32068 9335 32124
rect 9271 32064 9335 32068
rect 9351 32124 9415 32128
rect 9351 32068 9355 32124
rect 9355 32068 9411 32124
rect 9411 32068 9415 32124
rect 9351 32064 9415 32068
rect 10732 31996 10796 32060
rect 10548 31724 10612 31788
rect 4215 31580 4279 31584
rect 4215 31524 4219 31580
rect 4219 31524 4275 31580
rect 4275 31524 4279 31580
rect 4215 31520 4279 31524
rect 4295 31580 4359 31584
rect 4295 31524 4299 31580
rect 4299 31524 4355 31580
rect 4355 31524 4359 31580
rect 4295 31520 4359 31524
rect 4375 31580 4439 31584
rect 4375 31524 4379 31580
rect 4379 31524 4435 31580
rect 4435 31524 4439 31580
rect 4375 31520 4439 31524
rect 4455 31580 4519 31584
rect 4455 31524 4459 31580
rect 4459 31524 4515 31580
rect 4515 31524 4519 31580
rect 4455 31520 4519 31524
rect 7479 31580 7543 31584
rect 7479 31524 7483 31580
rect 7483 31524 7539 31580
rect 7539 31524 7543 31580
rect 7479 31520 7543 31524
rect 7559 31580 7623 31584
rect 7559 31524 7563 31580
rect 7563 31524 7619 31580
rect 7619 31524 7623 31580
rect 7559 31520 7623 31524
rect 7639 31580 7703 31584
rect 7639 31524 7643 31580
rect 7643 31524 7699 31580
rect 7699 31524 7703 31580
rect 7639 31520 7703 31524
rect 7719 31580 7783 31584
rect 7719 31524 7723 31580
rect 7723 31524 7779 31580
rect 7779 31524 7783 31580
rect 7719 31520 7783 31524
rect 2584 31036 2648 31040
rect 2584 30980 2588 31036
rect 2588 30980 2644 31036
rect 2644 30980 2648 31036
rect 2584 30976 2648 30980
rect 2664 31036 2728 31040
rect 2664 30980 2668 31036
rect 2668 30980 2724 31036
rect 2724 30980 2728 31036
rect 2664 30976 2728 30980
rect 2744 31036 2808 31040
rect 2744 30980 2748 31036
rect 2748 30980 2804 31036
rect 2804 30980 2808 31036
rect 2744 30976 2808 30980
rect 2824 31036 2888 31040
rect 2824 30980 2828 31036
rect 2828 30980 2884 31036
rect 2884 30980 2888 31036
rect 2824 30976 2888 30980
rect 5847 31036 5911 31040
rect 5847 30980 5851 31036
rect 5851 30980 5907 31036
rect 5907 30980 5911 31036
rect 5847 30976 5911 30980
rect 5927 31036 5991 31040
rect 5927 30980 5931 31036
rect 5931 30980 5987 31036
rect 5987 30980 5991 31036
rect 5927 30976 5991 30980
rect 6007 31036 6071 31040
rect 6007 30980 6011 31036
rect 6011 30980 6067 31036
rect 6067 30980 6071 31036
rect 6007 30976 6071 30980
rect 6087 31036 6151 31040
rect 6087 30980 6091 31036
rect 6091 30980 6147 31036
rect 6147 30980 6151 31036
rect 6087 30976 6151 30980
rect 9111 31036 9175 31040
rect 9111 30980 9115 31036
rect 9115 30980 9171 31036
rect 9171 30980 9175 31036
rect 9111 30976 9175 30980
rect 9191 31036 9255 31040
rect 9191 30980 9195 31036
rect 9195 30980 9251 31036
rect 9251 30980 9255 31036
rect 9191 30976 9255 30980
rect 9271 31036 9335 31040
rect 9271 30980 9275 31036
rect 9275 30980 9331 31036
rect 9331 30980 9335 31036
rect 9271 30976 9335 30980
rect 9351 31036 9415 31040
rect 9351 30980 9355 31036
rect 9355 30980 9411 31036
rect 9411 30980 9415 31036
rect 9351 30976 9415 30980
rect 9996 30772 10060 30836
rect 10732 30500 10796 30564
rect 4215 30492 4279 30496
rect 4215 30436 4219 30492
rect 4219 30436 4275 30492
rect 4275 30436 4279 30492
rect 4215 30432 4279 30436
rect 4295 30492 4359 30496
rect 4295 30436 4299 30492
rect 4299 30436 4355 30492
rect 4355 30436 4359 30492
rect 4295 30432 4359 30436
rect 4375 30492 4439 30496
rect 4375 30436 4379 30492
rect 4379 30436 4435 30492
rect 4435 30436 4439 30492
rect 4375 30432 4439 30436
rect 4455 30492 4519 30496
rect 4455 30436 4459 30492
rect 4459 30436 4515 30492
rect 4515 30436 4519 30492
rect 4455 30432 4519 30436
rect 7479 30492 7543 30496
rect 7479 30436 7483 30492
rect 7483 30436 7539 30492
rect 7539 30436 7543 30492
rect 7479 30432 7543 30436
rect 7559 30492 7623 30496
rect 7559 30436 7563 30492
rect 7563 30436 7619 30492
rect 7619 30436 7623 30492
rect 7559 30432 7623 30436
rect 7639 30492 7703 30496
rect 7639 30436 7643 30492
rect 7643 30436 7699 30492
rect 7699 30436 7703 30492
rect 7639 30432 7703 30436
rect 7719 30492 7783 30496
rect 7719 30436 7723 30492
rect 7723 30436 7779 30492
rect 7779 30436 7783 30492
rect 7719 30432 7783 30436
rect 2584 29948 2648 29952
rect 2584 29892 2588 29948
rect 2588 29892 2644 29948
rect 2644 29892 2648 29948
rect 2584 29888 2648 29892
rect 2664 29948 2728 29952
rect 2664 29892 2668 29948
rect 2668 29892 2724 29948
rect 2724 29892 2728 29948
rect 2664 29888 2728 29892
rect 2744 29948 2808 29952
rect 2744 29892 2748 29948
rect 2748 29892 2804 29948
rect 2804 29892 2808 29948
rect 2744 29888 2808 29892
rect 2824 29948 2888 29952
rect 2824 29892 2828 29948
rect 2828 29892 2884 29948
rect 2884 29892 2888 29948
rect 2824 29888 2888 29892
rect 5847 29948 5911 29952
rect 5847 29892 5851 29948
rect 5851 29892 5907 29948
rect 5907 29892 5911 29948
rect 5847 29888 5911 29892
rect 5927 29948 5991 29952
rect 5927 29892 5931 29948
rect 5931 29892 5987 29948
rect 5987 29892 5991 29948
rect 5927 29888 5991 29892
rect 6007 29948 6071 29952
rect 6007 29892 6011 29948
rect 6011 29892 6067 29948
rect 6067 29892 6071 29948
rect 6007 29888 6071 29892
rect 6087 29948 6151 29952
rect 6087 29892 6091 29948
rect 6091 29892 6147 29948
rect 6147 29892 6151 29948
rect 6087 29888 6151 29892
rect 9111 29948 9175 29952
rect 9111 29892 9115 29948
rect 9115 29892 9171 29948
rect 9171 29892 9175 29948
rect 9111 29888 9175 29892
rect 9191 29948 9255 29952
rect 9191 29892 9195 29948
rect 9195 29892 9251 29948
rect 9251 29892 9255 29948
rect 9191 29888 9255 29892
rect 9271 29948 9335 29952
rect 9271 29892 9275 29948
rect 9275 29892 9331 29948
rect 9331 29892 9335 29948
rect 9271 29888 9335 29892
rect 9351 29948 9415 29952
rect 9351 29892 9355 29948
rect 9355 29892 9411 29948
rect 9411 29892 9415 29948
rect 9351 29888 9415 29892
rect 9812 29684 9876 29748
rect 11652 29684 11716 29748
rect 10180 29608 10244 29612
rect 10180 29552 10194 29608
rect 10194 29552 10244 29608
rect 10180 29548 10244 29552
rect 4215 29404 4279 29408
rect 4215 29348 4219 29404
rect 4219 29348 4275 29404
rect 4275 29348 4279 29404
rect 4215 29344 4279 29348
rect 4295 29404 4359 29408
rect 4295 29348 4299 29404
rect 4299 29348 4355 29404
rect 4355 29348 4359 29404
rect 4295 29344 4359 29348
rect 4375 29404 4439 29408
rect 4375 29348 4379 29404
rect 4379 29348 4435 29404
rect 4435 29348 4439 29404
rect 4375 29344 4439 29348
rect 4455 29404 4519 29408
rect 4455 29348 4459 29404
rect 4459 29348 4515 29404
rect 4515 29348 4519 29404
rect 4455 29344 4519 29348
rect 7479 29404 7543 29408
rect 7479 29348 7483 29404
rect 7483 29348 7539 29404
rect 7539 29348 7543 29404
rect 7479 29344 7543 29348
rect 7559 29404 7623 29408
rect 7559 29348 7563 29404
rect 7563 29348 7619 29404
rect 7619 29348 7623 29404
rect 7559 29344 7623 29348
rect 7639 29404 7703 29408
rect 7639 29348 7643 29404
rect 7643 29348 7699 29404
rect 7699 29348 7703 29404
rect 7639 29344 7703 29348
rect 7719 29404 7783 29408
rect 7719 29348 7723 29404
rect 7723 29348 7779 29404
rect 7779 29348 7783 29404
rect 7719 29344 7783 29348
rect 10916 29276 10980 29340
rect 2584 28860 2648 28864
rect 2584 28804 2588 28860
rect 2588 28804 2644 28860
rect 2644 28804 2648 28860
rect 2584 28800 2648 28804
rect 2664 28860 2728 28864
rect 2664 28804 2668 28860
rect 2668 28804 2724 28860
rect 2724 28804 2728 28860
rect 2664 28800 2728 28804
rect 2744 28860 2808 28864
rect 2744 28804 2748 28860
rect 2748 28804 2804 28860
rect 2804 28804 2808 28860
rect 2744 28800 2808 28804
rect 2824 28860 2888 28864
rect 2824 28804 2828 28860
rect 2828 28804 2884 28860
rect 2884 28804 2888 28860
rect 2824 28800 2888 28804
rect 5847 28860 5911 28864
rect 5847 28804 5851 28860
rect 5851 28804 5907 28860
rect 5907 28804 5911 28860
rect 5847 28800 5911 28804
rect 5927 28860 5991 28864
rect 5927 28804 5931 28860
rect 5931 28804 5987 28860
rect 5987 28804 5991 28860
rect 5927 28800 5991 28804
rect 6007 28860 6071 28864
rect 6007 28804 6011 28860
rect 6011 28804 6067 28860
rect 6067 28804 6071 28860
rect 6007 28800 6071 28804
rect 6087 28860 6151 28864
rect 6087 28804 6091 28860
rect 6091 28804 6147 28860
rect 6147 28804 6151 28860
rect 6087 28800 6151 28804
rect 9111 28860 9175 28864
rect 9111 28804 9115 28860
rect 9115 28804 9171 28860
rect 9171 28804 9175 28860
rect 9111 28800 9175 28804
rect 9191 28860 9255 28864
rect 9191 28804 9195 28860
rect 9195 28804 9251 28860
rect 9251 28804 9255 28860
rect 9191 28800 9255 28804
rect 9271 28860 9335 28864
rect 9271 28804 9275 28860
rect 9275 28804 9331 28860
rect 9331 28804 9335 28860
rect 9271 28800 9335 28804
rect 9351 28860 9415 28864
rect 9351 28804 9355 28860
rect 9355 28804 9411 28860
rect 9411 28804 9415 28860
rect 9351 28800 9415 28804
rect 4215 28316 4279 28320
rect 4215 28260 4219 28316
rect 4219 28260 4275 28316
rect 4275 28260 4279 28316
rect 4215 28256 4279 28260
rect 4295 28316 4359 28320
rect 4295 28260 4299 28316
rect 4299 28260 4355 28316
rect 4355 28260 4359 28316
rect 4295 28256 4359 28260
rect 4375 28316 4439 28320
rect 4375 28260 4379 28316
rect 4379 28260 4435 28316
rect 4435 28260 4439 28316
rect 4375 28256 4439 28260
rect 4455 28316 4519 28320
rect 4455 28260 4459 28316
rect 4459 28260 4515 28316
rect 4515 28260 4519 28316
rect 4455 28256 4519 28260
rect 7479 28316 7543 28320
rect 7479 28260 7483 28316
rect 7483 28260 7539 28316
rect 7539 28260 7543 28316
rect 7479 28256 7543 28260
rect 7559 28316 7623 28320
rect 7559 28260 7563 28316
rect 7563 28260 7619 28316
rect 7619 28260 7623 28316
rect 7559 28256 7623 28260
rect 7639 28316 7703 28320
rect 7639 28260 7643 28316
rect 7643 28260 7699 28316
rect 7699 28260 7703 28316
rect 7639 28256 7703 28260
rect 7719 28316 7783 28320
rect 7719 28260 7723 28316
rect 7723 28260 7779 28316
rect 7779 28260 7783 28316
rect 7719 28256 7783 28260
rect 10364 28188 10428 28252
rect 2584 27772 2648 27776
rect 2584 27716 2588 27772
rect 2588 27716 2644 27772
rect 2644 27716 2648 27772
rect 2584 27712 2648 27716
rect 2664 27772 2728 27776
rect 2664 27716 2668 27772
rect 2668 27716 2724 27772
rect 2724 27716 2728 27772
rect 2664 27712 2728 27716
rect 2744 27772 2808 27776
rect 2744 27716 2748 27772
rect 2748 27716 2804 27772
rect 2804 27716 2808 27772
rect 2744 27712 2808 27716
rect 2824 27772 2888 27776
rect 2824 27716 2828 27772
rect 2828 27716 2884 27772
rect 2884 27716 2888 27772
rect 2824 27712 2888 27716
rect 5847 27772 5911 27776
rect 5847 27716 5851 27772
rect 5851 27716 5907 27772
rect 5907 27716 5911 27772
rect 5847 27712 5911 27716
rect 5927 27772 5991 27776
rect 5927 27716 5931 27772
rect 5931 27716 5987 27772
rect 5987 27716 5991 27772
rect 5927 27712 5991 27716
rect 6007 27772 6071 27776
rect 6007 27716 6011 27772
rect 6011 27716 6067 27772
rect 6067 27716 6071 27772
rect 6007 27712 6071 27716
rect 6087 27772 6151 27776
rect 6087 27716 6091 27772
rect 6091 27716 6147 27772
rect 6147 27716 6151 27772
rect 6087 27712 6151 27716
rect 9111 27772 9175 27776
rect 9111 27716 9115 27772
rect 9115 27716 9171 27772
rect 9171 27716 9175 27772
rect 9111 27712 9175 27716
rect 9191 27772 9255 27776
rect 9191 27716 9195 27772
rect 9195 27716 9251 27772
rect 9251 27716 9255 27772
rect 9191 27712 9255 27716
rect 9271 27772 9335 27776
rect 9271 27716 9275 27772
rect 9275 27716 9331 27772
rect 9331 27716 9335 27772
rect 9271 27712 9335 27716
rect 9351 27772 9415 27776
rect 9351 27716 9355 27772
rect 9355 27716 9411 27772
rect 9411 27716 9415 27772
rect 9351 27712 9415 27716
rect 4215 27228 4279 27232
rect 4215 27172 4219 27228
rect 4219 27172 4275 27228
rect 4275 27172 4279 27228
rect 4215 27168 4279 27172
rect 4295 27228 4359 27232
rect 4295 27172 4299 27228
rect 4299 27172 4355 27228
rect 4355 27172 4359 27228
rect 4295 27168 4359 27172
rect 4375 27228 4439 27232
rect 4375 27172 4379 27228
rect 4379 27172 4435 27228
rect 4435 27172 4439 27228
rect 4375 27168 4439 27172
rect 4455 27228 4519 27232
rect 4455 27172 4459 27228
rect 4459 27172 4515 27228
rect 4515 27172 4519 27228
rect 4455 27168 4519 27172
rect 7479 27228 7543 27232
rect 7479 27172 7483 27228
rect 7483 27172 7539 27228
rect 7539 27172 7543 27228
rect 7479 27168 7543 27172
rect 7559 27228 7623 27232
rect 7559 27172 7563 27228
rect 7563 27172 7619 27228
rect 7619 27172 7623 27228
rect 7559 27168 7623 27172
rect 7639 27228 7703 27232
rect 7639 27172 7643 27228
rect 7643 27172 7699 27228
rect 7699 27172 7703 27228
rect 7639 27168 7703 27172
rect 7719 27228 7783 27232
rect 7719 27172 7723 27228
rect 7723 27172 7779 27228
rect 7779 27172 7783 27228
rect 7719 27168 7783 27172
rect 2584 26684 2648 26688
rect 2584 26628 2588 26684
rect 2588 26628 2644 26684
rect 2644 26628 2648 26684
rect 2584 26624 2648 26628
rect 2664 26684 2728 26688
rect 2664 26628 2668 26684
rect 2668 26628 2724 26684
rect 2724 26628 2728 26684
rect 2664 26624 2728 26628
rect 2744 26684 2808 26688
rect 2744 26628 2748 26684
rect 2748 26628 2804 26684
rect 2804 26628 2808 26684
rect 2744 26624 2808 26628
rect 2824 26684 2888 26688
rect 2824 26628 2828 26684
rect 2828 26628 2884 26684
rect 2884 26628 2888 26684
rect 2824 26624 2888 26628
rect 5847 26684 5911 26688
rect 5847 26628 5851 26684
rect 5851 26628 5907 26684
rect 5907 26628 5911 26684
rect 5847 26624 5911 26628
rect 5927 26684 5991 26688
rect 5927 26628 5931 26684
rect 5931 26628 5987 26684
rect 5987 26628 5991 26684
rect 5927 26624 5991 26628
rect 6007 26684 6071 26688
rect 6007 26628 6011 26684
rect 6011 26628 6067 26684
rect 6067 26628 6071 26684
rect 6007 26624 6071 26628
rect 6087 26684 6151 26688
rect 6087 26628 6091 26684
rect 6091 26628 6147 26684
rect 6147 26628 6151 26684
rect 6087 26624 6151 26628
rect 9111 26684 9175 26688
rect 9111 26628 9115 26684
rect 9115 26628 9171 26684
rect 9171 26628 9175 26684
rect 9111 26624 9175 26628
rect 9191 26684 9255 26688
rect 9191 26628 9195 26684
rect 9195 26628 9251 26684
rect 9251 26628 9255 26684
rect 9191 26624 9255 26628
rect 9271 26684 9335 26688
rect 9271 26628 9275 26684
rect 9275 26628 9331 26684
rect 9331 26628 9335 26684
rect 9271 26624 9335 26628
rect 9351 26684 9415 26688
rect 9351 26628 9355 26684
rect 9355 26628 9411 26684
rect 9411 26628 9415 26684
rect 9351 26624 9415 26628
rect 4215 26140 4279 26144
rect 4215 26084 4219 26140
rect 4219 26084 4275 26140
rect 4275 26084 4279 26140
rect 4215 26080 4279 26084
rect 4295 26140 4359 26144
rect 4295 26084 4299 26140
rect 4299 26084 4355 26140
rect 4355 26084 4359 26140
rect 4295 26080 4359 26084
rect 4375 26140 4439 26144
rect 4375 26084 4379 26140
rect 4379 26084 4435 26140
rect 4435 26084 4439 26140
rect 4375 26080 4439 26084
rect 4455 26140 4519 26144
rect 4455 26084 4459 26140
rect 4459 26084 4515 26140
rect 4515 26084 4519 26140
rect 4455 26080 4519 26084
rect 7479 26140 7543 26144
rect 7479 26084 7483 26140
rect 7483 26084 7539 26140
rect 7539 26084 7543 26140
rect 7479 26080 7543 26084
rect 7559 26140 7623 26144
rect 7559 26084 7563 26140
rect 7563 26084 7619 26140
rect 7619 26084 7623 26140
rect 7559 26080 7623 26084
rect 7639 26140 7703 26144
rect 7639 26084 7643 26140
rect 7643 26084 7699 26140
rect 7699 26084 7703 26140
rect 7639 26080 7703 26084
rect 7719 26140 7783 26144
rect 7719 26084 7723 26140
rect 7723 26084 7779 26140
rect 7779 26084 7783 26140
rect 7719 26080 7783 26084
rect 2584 25596 2648 25600
rect 2584 25540 2588 25596
rect 2588 25540 2644 25596
rect 2644 25540 2648 25596
rect 2584 25536 2648 25540
rect 2664 25596 2728 25600
rect 2664 25540 2668 25596
rect 2668 25540 2724 25596
rect 2724 25540 2728 25596
rect 2664 25536 2728 25540
rect 2744 25596 2808 25600
rect 2744 25540 2748 25596
rect 2748 25540 2804 25596
rect 2804 25540 2808 25596
rect 2744 25536 2808 25540
rect 2824 25596 2888 25600
rect 2824 25540 2828 25596
rect 2828 25540 2884 25596
rect 2884 25540 2888 25596
rect 2824 25536 2888 25540
rect 5847 25596 5911 25600
rect 5847 25540 5851 25596
rect 5851 25540 5907 25596
rect 5907 25540 5911 25596
rect 5847 25536 5911 25540
rect 5927 25596 5991 25600
rect 5927 25540 5931 25596
rect 5931 25540 5987 25596
rect 5987 25540 5991 25596
rect 5927 25536 5991 25540
rect 6007 25596 6071 25600
rect 6007 25540 6011 25596
rect 6011 25540 6067 25596
rect 6067 25540 6071 25596
rect 6007 25536 6071 25540
rect 6087 25596 6151 25600
rect 6087 25540 6091 25596
rect 6091 25540 6147 25596
rect 6147 25540 6151 25596
rect 6087 25536 6151 25540
rect 9111 25596 9175 25600
rect 9111 25540 9115 25596
rect 9115 25540 9171 25596
rect 9171 25540 9175 25596
rect 9111 25536 9175 25540
rect 9191 25596 9255 25600
rect 9191 25540 9195 25596
rect 9195 25540 9251 25596
rect 9251 25540 9255 25596
rect 9191 25536 9255 25540
rect 9271 25596 9335 25600
rect 9271 25540 9275 25596
rect 9275 25540 9331 25596
rect 9331 25540 9335 25596
rect 9271 25536 9335 25540
rect 9351 25596 9415 25600
rect 9351 25540 9355 25596
rect 9355 25540 9411 25596
rect 9411 25540 9415 25596
rect 9351 25536 9415 25540
rect 4215 25052 4279 25056
rect 4215 24996 4219 25052
rect 4219 24996 4275 25052
rect 4275 24996 4279 25052
rect 4215 24992 4279 24996
rect 4295 25052 4359 25056
rect 4295 24996 4299 25052
rect 4299 24996 4355 25052
rect 4355 24996 4359 25052
rect 4295 24992 4359 24996
rect 4375 25052 4439 25056
rect 4375 24996 4379 25052
rect 4379 24996 4435 25052
rect 4435 24996 4439 25052
rect 4375 24992 4439 24996
rect 4455 25052 4519 25056
rect 4455 24996 4459 25052
rect 4459 24996 4515 25052
rect 4515 24996 4519 25052
rect 4455 24992 4519 24996
rect 7479 25052 7543 25056
rect 7479 24996 7483 25052
rect 7483 24996 7539 25052
rect 7539 24996 7543 25052
rect 7479 24992 7543 24996
rect 7559 25052 7623 25056
rect 7559 24996 7563 25052
rect 7563 24996 7619 25052
rect 7619 24996 7623 25052
rect 7559 24992 7623 24996
rect 7639 25052 7703 25056
rect 7639 24996 7643 25052
rect 7643 24996 7699 25052
rect 7699 24996 7703 25052
rect 7639 24992 7703 24996
rect 7719 25052 7783 25056
rect 7719 24996 7723 25052
rect 7723 24996 7779 25052
rect 7779 24996 7783 25052
rect 7719 24992 7783 24996
rect 2584 24508 2648 24512
rect 2584 24452 2588 24508
rect 2588 24452 2644 24508
rect 2644 24452 2648 24508
rect 2584 24448 2648 24452
rect 2664 24508 2728 24512
rect 2664 24452 2668 24508
rect 2668 24452 2724 24508
rect 2724 24452 2728 24508
rect 2664 24448 2728 24452
rect 2744 24508 2808 24512
rect 2744 24452 2748 24508
rect 2748 24452 2804 24508
rect 2804 24452 2808 24508
rect 2744 24448 2808 24452
rect 2824 24508 2888 24512
rect 2824 24452 2828 24508
rect 2828 24452 2884 24508
rect 2884 24452 2888 24508
rect 2824 24448 2888 24452
rect 5847 24508 5911 24512
rect 5847 24452 5851 24508
rect 5851 24452 5907 24508
rect 5907 24452 5911 24508
rect 5847 24448 5911 24452
rect 5927 24508 5991 24512
rect 5927 24452 5931 24508
rect 5931 24452 5987 24508
rect 5987 24452 5991 24508
rect 5927 24448 5991 24452
rect 6007 24508 6071 24512
rect 6007 24452 6011 24508
rect 6011 24452 6067 24508
rect 6067 24452 6071 24508
rect 6007 24448 6071 24452
rect 6087 24508 6151 24512
rect 6087 24452 6091 24508
rect 6091 24452 6147 24508
rect 6147 24452 6151 24508
rect 6087 24448 6151 24452
rect 9111 24508 9175 24512
rect 9111 24452 9115 24508
rect 9115 24452 9171 24508
rect 9171 24452 9175 24508
rect 9111 24448 9175 24452
rect 9191 24508 9255 24512
rect 9191 24452 9195 24508
rect 9195 24452 9251 24508
rect 9251 24452 9255 24508
rect 9191 24448 9255 24452
rect 9271 24508 9335 24512
rect 9271 24452 9275 24508
rect 9275 24452 9331 24508
rect 9331 24452 9335 24508
rect 9271 24448 9335 24452
rect 9351 24508 9415 24512
rect 9351 24452 9355 24508
rect 9355 24452 9411 24508
rect 9411 24452 9415 24508
rect 9351 24448 9415 24452
rect 4215 23964 4279 23968
rect 4215 23908 4219 23964
rect 4219 23908 4275 23964
rect 4275 23908 4279 23964
rect 4215 23904 4279 23908
rect 4295 23964 4359 23968
rect 4295 23908 4299 23964
rect 4299 23908 4355 23964
rect 4355 23908 4359 23964
rect 4295 23904 4359 23908
rect 4375 23964 4439 23968
rect 4375 23908 4379 23964
rect 4379 23908 4435 23964
rect 4435 23908 4439 23964
rect 4375 23904 4439 23908
rect 4455 23964 4519 23968
rect 4455 23908 4459 23964
rect 4459 23908 4515 23964
rect 4515 23908 4519 23964
rect 4455 23904 4519 23908
rect 7479 23964 7543 23968
rect 7479 23908 7483 23964
rect 7483 23908 7539 23964
rect 7539 23908 7543 23964
rect 7479 23904 7543 23908
rect 7559 23964 7623 23968
rect 7559 23908 7563 23964
rect 7563 23908 7619 23964
rect 7619 23908 7623 23964
rect 7559 23904 7623 23908
rect 7639 23964 7703 23968
rect 7639 23908 7643 23964
rect 7643 23908 7699 23964
rect 7699 23908 7703 23964
rect 7639 23904 7703 23908
rect 7719 23964 7783 23968
rect 7719 23908 7723 23964
rect 7723 23908 7779 23964
rect 7779 23908 7783 23964
rect 7719 23904 7783 23908
rect 2584 23420 2648 23424
rect 2584 23364 2588 23420
rect 2588 23364 2644 23420
rect 2644 23364 2648 23420
rect 2584 23360 2648 23364
rect 2664 23420 2728 23424
rect 2664 23364 2668 23420
rect 2668 23364 2724 23420
rect 2724 23364 2728 23420
rect 2664 23360 2728 23364
rect 2744 23420 2808 23424
rect 2744 23364 2748 23420
rect 2748 23364 2804 23420
rect 2804 23364 2808 23420
rect 2744 23360 2808 23364
rect 2824 23420 2888 23424
rect 2824 23364 2828 23420
rect 2828 23364 2884 23420
rect 2884 23364 2888 23420
rect 2824 23360 2888 23364
rect 5847 23420 5911 23424
rect 5847 23364 5851 23420
rect 5851 23364 5907 23420
rect 5907 23364 5911 23420
rect 5847 23360 5911 23364
rect 5927 23420 5991 23424
rect 5927 23364 5931 23420
rect 5931 23364 5987 23420
rect 5987 23364 5991 23420
rect 5927 23360 5991 23364
rect 6007 23420 6071 23424
rect 6007 23364 6011 23420
rect 6011 23364 6067 23420
rect 6067 23364 6071 23420
rect 6007 23360 6071 23364
rect 6087 23420 6151 23424
rect 6087 23364 6091 23420
rect 6091 23364 6147 23420
rect 6147 23364 6151 23420
rect 6087 23360 6151 23364
rect 9111 23420 9175 23424
rect 9111 23364 9115 23420
rect 9115 23364 9171 23420
rect 9171 23364 9175 23420
rect 9111 23360 9175 23364
rect 9191 23420 9255 23424
rect 9191 23364 9195 23420
rect 9195 23364 9251 23420
rect 9251 23364 9255 23420
rect 9191 23360 9255 23364
rect 9271 23420 9335 23424
rect 9271 23364 9275 23420
rect 9275 23364 9331 23420
rect 9331 23364 9335 23420
rect 9271 23360 9335 23364
rect 9351 23420 9415 23424
rect 9351 23364 9355 23420
rect 9355 23364 9411 23420
rect 9411 23364 9415 23420
rect 9351 23360 9415 23364
rect 4215 22876 4279 22880
rect 4215 22820 4219 22876
rect 4219 22820 4275 22876
rect 4275 22820 4279 22876
rect 4215 22816 4279 22820
rect 4295 22876 4359 22880
rect 4295 22820 4299 22876
rect 4299 22820 4355 22876
rect 4355 22820 4359 22876
rect 4295 22816 4359 22820
rect 4375 22876 4439 22880
rect 4375 22820 4379 22876
rect 4379 22820 4435 22876
rect 4435 22820 4439 22876
rect 4375 22816 4439 22820
rect 4455 22876 4519 22880
rect 4455 22820 4459 22876
rect 4459 22820 4515 22876
rect 4515 22820 4519 22876
rect 4455 22816 4519 22820
rect 7479 22876 7543 22880
rect 7479 22820 7483 22876
rect 7483 22820 7539 22876
rect 7539 22820 7543 22876
rect 7479 22816 7543 22820
rect 7559 22876 7623 22880
rect 7559 22820 7563 22876
rect 7563 22820 7619 22876
rect 7619 22820 7623 22876
rect 7559 22816 7623 22820
rect 7639 22876 7703 22880
rect 7639 22820 7643 22876
rect 7643 22820 7699 22876
rect 7699 22820 7703 22876
rect 7639 22816 7703 22820
rect 7719 22876 7783 22880
rect 7719 22820 7723 22876
rect 7723 22820 7779 22876
rect 7779 22820 7783 22876
rect 7719 22816 7783 22820
rect 2584 22332 2648 22336
rect 2584 22276 2588 22332
rect 2588 22276 2644 22332
rect 2644 22276 2648 22332
rect 2584 22272 2648 22276
rect 2664 22332 2728 22336
rect 2664 22276 2668 22332
rect 2668 22276 2724 22332
rect 2724 22276 2728 22332
rect 2664 22272 2728 22276
rect 2744 22332 2808 22336
rect 2744 22276 2748 22332
rect 2748 22276 2804 22332
rect 2804 22276 2808 22332
rect 2744 22272 2808 22276
rect 2824 22332 2888 22336
rect 2824 22276 2828 22332
rect 2828 22276 2884 22332
rect 2884 22276 2888 22332
rect 2824 22272 2888 22276
rect 5847 22332 5911 22336
rect 5847 22276 5851 22332
rect 5851 22276 5907 22332
rect 5907 22276 5911 22332
rect 5847 22272 5911 22276
rect 5927 22332 5991 22336
rect 5927 22276 5931 22332
rect 5931 22276 5987 22332
rect 5987 22276 5991 22332
rect 5927 22272 5991 22276
rect 6007 22332 6071 22336
rect 6007 22276 6011 22332
rect 6011 22276 6067 22332
rect 6067 22276 6071 22332
rect 6007 22272 6071 22276
rect 6087 22332 6151 22336
rect 6087 22276 6091 22332
rect 6091 22276 6147 22332
rect 6147 22276 6151 22332
rect 6087 22272 6151 22276
rect 9111 22332 9175 22336
rect 9111 22276 9115 22332
rect 9115 22276 9171 22332
rect 9171 22276 9175 22332
rect 9111 22272 9175 22276
rect 9191 22332 9255 22336
rect 9191 22276 9195 22332
rect 9195 22276 9251 22332
rect 9251 22276 9255 22332
rect 9191 22272 9255 22276
rect 9271 22332 9335 22336
rect 9271 22276 9275 22332
rect 9275 22276 9331 22332
rect 9331 22276 9335 22332
rect 9271 22272 9335 22276
rect 9351 22332 9415 22336
rect 9351 22276 9355 22332
rect 9355 22276 9411 22332
rect 9411 22276 9415 22332
rect 9351 22272 9415 22276
rect 10916 22264 10980 22268
rect 10916 22208 10966 22264
rect 10966 22208 10980 22264
rect 10916 22204 10980 22208
rect 4215 21788 4279 21792
rect 4215 21732 4219 21788
rect 4219 21732 4275 21788
rect 4275 21732 4279 21788
rect 4215 21728 4279 21732
rect 4295 21788 4359 21792
rect 4295 21732 4299 21788
rect 4299 21732 4355 21788
rect 4355 21732 4359 21788
rect 4295 21728 4359 21732
rect 4375 21788 4439 21792
rect 4375 21732 4379 21788
rect 4379 21732 4435 21788
rect 4435 21732 4439 21788
rect 4375 21728 4439 21732
rect 4455 21788 4519 21792
rect 4455 21732 4459 21788
rect 4459 21732 4515 21788
rect 4515 21732 4519 21788
rect 4455 21728 4519 21732
rect 7479 21788 7543 21792
rect 7479 21732 7483 21788
rect 7483 21732 7539 21788
rect 7539 21732 7543 21788
rect 7479 21728 7543 21732
rect 7559 21788 7623 21792
rect 7559 21732 7563 21788
rect 7563 21732 7619 21788
rect 7619 21732 7623 21788
rect 7559 21728 7623 21732
rect 7639 21788 7703 21792
rect 7639 21732 7643 21788
rect 7643 21732 7699 21788
rect 7699 21732 7703 21788
rect 7639 21728 7703 21732
rect 7719 21788 7783 21792
rect 7719 21732 7723 21788
rect 7723 21732 7779 21788
rect 7779 21732 7783 21788
rect 7719 21728 7783 21732
rect 2584 21244 2648 21248
rect 2584 21188 2588 21244
rect 2588 21188 2644 21244
rect 2644 21188 2648 21244
rect 2584 21184 2648 21188
rect 2664 21244 2728 21248
rect 2664 21188 2668 21244
rect 2668 21188 2724 21244
rect 2724 21188 2728 21244
rect 2664 21184 2728 21188
rect 2744 21244 2808 21248
rect 2744 21188 2748 21244
rect 2748 21188 2804 21244
rect 2804 21188 2808 21244
rect 2744 21184 2808 21188
rect 2824 21244 2888 21248
rect 2824 21188 2828 21244
rect 2828 21188 2884 21244
rect 2884 21188 2888 21244
rect 2824 21184 2888 21188
rect 5847 21244 5911 21248
rect 5847 21188 5851 21244
rect 5851 21188 5907 21244
rect 5907 21188 5911 21244
rect 5847 21184 5911 21188
rect 5927 21244 5991 21248
rect 5927 21188 5931 21244
rect 5931 21188 5987 21244
rect 5987 21188 5991 21244
rect 5927 21184 5991 21188
rect 6007 21244 6071 21248
rect 6007 21188 6011 21244
rect 6011 21188 6067 21244
rect 6067 21188 6071 21244
rect 6007 21184 6071 21188
rect 6087 21244 6151 21248
rect 6087 21188 6091 21244
rect 6091 21188 6147 21244
rect 6147 21188 6151 21244
rect 6087 21184 6151 21188
rect 9111 21244 9175 21248
rect 9111 21188 9115 21244
rect 9115 21188 9171 21244
rect 9171 21188 9175 21244
rect 9111 21184 9175 21188
rect 9191 21244 9255 21248
rect 9191 21188 9195 21244
rect 9195 21188 9251 21244
rect 9251 21188 9255 21244
rect 9191 21184 9255 21188
rect 9271 21244 9335 21248
rect 9271 21188 9275 21244
rect 9275 21188 9331 21244
rect 9331 21188 9335 21244
rect 9271 21184 9335 21188
rect 9351 21244 9415 21248
rect 9351 21188 9355 21244
rect 9355 21188 9411 21244
rect 9411 21188 9415 21244
rect 9351 21184 9415 21188
rect 4215 20700 4279 20704
rect 4215 20644 4219 20700
rect 4219 20644 4275 20700
rect 4275 20644 4279 20700
rect 4215 20640 4279 20644
rect 4295 20700 4359 20704
rect 4295 20644 4299 20700
rect 4299 20644 4355 20700
rect 4355 20644 4359 20700
rect 4295 20640 4359 20644
rect 4375 20700 4439 20704
rect 4375 20644 4379 20700
rect 4379 20644 4435 20700
rect 4435 20644 4439 20700
rect 4375 20640 4439 20644
rect 4455 20700 4519 20704
rect 4455 20644 4459 20700
rect 4459 20644 4515 20700
rect 4515 20644 4519 20700
rect 4455 20640 4519 20644
rect 7479 20700 7543 20704
rect 7479 20644 7483 20700
rect 7483 20644 7539 20700
rect 7539 20644 7543 20700
rect 7479 20640 7543 20644
rect 7559 20700 7623 20704
rect 7559 20644 7563 20700
rect 7563 20644 7619 20700
rect 7619 20644 7623 20700
rect 7559 20640 7623 20644
rect 7639 20700 7703 20704
rect 7639 20644 7643 20700
rect 7643 20644 7699 20700
rect 7699 20644 7703 20700
rect 7639 20640 7703 20644
rect 7719 20700 7783 20704
rect 7719 20644 7723 20700
rect 7723 20644 7779 20700
rect 7779 20644 7783 20700
rect 7719 20640 7783 20644
rect 2584 20156 2648 20160
rect 2584 20100 2588 20156
rect 2588 20100 2644 20156
rect 2644 20100 2648 20156
rect 2584 20096 2648 20100
rect 2664 20156 2728 20160
rect 2664 20100 2668 20156
rect 2668 20100 2724 20156
rect 2724 20100 2728 20156
rect 2664 20096 2728 20100
rect 2744 20156 2808 20160
rect 2744 20100 2748 20156
rect 2748 20100 2804 20156
rect 2804 20100 2808 20156
rect 2744 20096 2808 20100
rect 2824 20156 2888 20160
rect 2824 20100 2828 20156
rect 2828 20100 2884 20156
rect 2884 20100 2888 20156
rect 2824 20096 2888 20100
rect 5847 20156 5911 20160
rect 5847 20100 5851 20156
rect 5851 20100 5907 20156
rect 5907 20100 5911 20156
rect 5847 20096 5911 20100
rect 5927 20156 5991 20160
rect 5927 20100 5931 20156
rect 5931 20100 5987 20156
rect 5987 20100 5991 20156
rect 5927 20096 5991 20100
rect 6007 20156 6071 20160
rect 6007 20100 6011 20156
rect 6011 20100 6067 20156
rect 6067 20100 6071 20156
rect 6007 20096 6071 20100
rect 6087 20156 6151 20160
rect 6087 20100 6091 20156
rect 6091 20100 6147 20156
rect 6147 20100 6151 20156
rect 6087 20096 6151 20100
rect 9111 20156 9175 20160
rect 9111 20100 9115 20156
rect 9115 20100 9171 20156
rect 9171 20100 9175 20156
rect 9111 20096 9175 20100
rect 9191 20156 9255 20160
rect 9191 20100 9195 20156
rect 9195 20100 9251 20156
rect 9251 20100 9255 20156
rect 9191 20096 9255 20100
rect 9271 20156 9335 20160
rect 9271 20100 9275 20156
rect 9275 20100 9331 20156
rect 9331 20100 9335 20156
rect 9271 20096 9335 20100
rect 9351 20156 9415 20160
rect 9351 20100 9355 20156
rect 9355 20100 9411 20156
rect 9411 20100 9415 20156
rect 9351 20096 9415 20100
rect 4215 19612 4279 19616
rect 4215 19556 4219 19612
rect 4219 19556 4275 19612
rect 4275 19556 4279 19612
rect 4215 19552 4279 19556
rect 4295 19612 4359 19616
rect 4295 19556 4299 19612
rect 4299 19556 4355 19612
rect 4355 19556 4359 19612
rect 4295 19552 4359 19556
rect 4375 19612 4439 19616
rect 4375 19556 4379 19612
rect 4379 19556 4435 19612
rect 4435 19556 4439 19612
rect 4375 19552 4439 19556
rect 4455 19612 4519 19616
rect 4455 19556 4459 19612
rect 4459 19556 4515 19612
rect 4515 19556 4519 19612
rect 4455 19552 4519 19556
rect 7479 19612 7543 19616
rect 7479 19556 7483 19612
rect 7483 19556 7539 19612
rect 7539 19556 7543 19612
rect 7479 19552 7543 19556
rect 7559 19612 7623 19616
rect 7559 19556 7563 19612
rect 7563 19556 7619 19612
rect 7619 19556 7623 19612
rect 7559 19552 7623 19556
rect 7639 19612 7703 19616
rect 7639 19556 7643 19612
rect 7643 19556 7699 19612
rect 7699 19556 7703 19612
rect 7639 19552 7703 19556
rect 7719 19612 7783 19616
rect 7719 19556 7723 19612
rect 7723 19556 7779 19612
rect 7779 19556 7783 19612
rect 7719 19552 7783 19556
rect 2584 19068 2648 19072
rect 2584 19012 2588 19068
rect 2588 19012 2644 19068
rect 2644 19012 2648 19068
rect 2584 19008 2648 19012
rect 2664 19068 2728 19072
rect 2664 19012 2668 19068
rect 2668 19012 2724 19068
rect 2724 19012 2728 19068
rect 2664 19008 2728 19012
rect 2744 19068 2808 19072
rect 2744 19012 2748 19068
rect 2748 19012 2804 19068
rect 2804 19012 2808 19068
rect 2744 19008 2808 19012
rect 2824 19068 2888 19072
rect 2824 19012 2828 19068
rect 2828 19012 2884 19068
rect 2884 19012 2888 19068
rect 2824 19008 2888 19012
rect 5847 19068 5911 19072
rect 5847 19012 5851 19068
rect 5851 19012 5907 19068
rect 5907 19012 5911 19068
rect 5847 19008 5911 19012
rect 5927 19068 5991 19072
rect 5927 19012 5931 19068
rect 5931 19012 5987 19068
rect 5987 19012 5991 19068
rect 5927 19008 5991 19012
rect 6007 19068 6071 19072
rect 6007 19012 6011 19068
rect 6011 19012 6067 19068
rect 6067 19012 6071 19068
rect 6007 19008 6071 19012
rect 6087 19068 6151 19072
rect 6087 19012 6091 19068
rect 6091 19012 6147 19068
rect 6147 19012 6151 19068
rect 6087 19008 6151 19012
rect 9111 19068 9175 19072
rect 9111 19012 9115 19068
rect 9115 19012 9171 19068
rect 9171 19012 9175 19068
rect 9111 19008 9175 19012
rect 9191 19068 9255 19072
rect 9191 19012 9195 19068
rect 9195 19012 9251 19068
rect 9251 19012 9255 19068
rect 9191 19008 9255 19012
rect 9271 19068 9335 19072
rect 9271 19012 9275 19068
rect 9275 19012 9331 19068
rect 9331 19012 9335 19068
rect 9271 19008 9335 19012
rect 9351 19068 9415 19072
rect 9351 19012 9355 19068
rect 9355 19012 9411 19068
rect 9411 19012 9415 19068
rect 9351 19008 9415 19012
rect 4215 18524 4279 18528
rect 4215 18468 4219 18524
rect 4219 18468 4275 18524
rect 4275 18468 4279 18524
rect 4215 18464 4279 18468
rect 4295 18524 4359 18528
rect 4295 18468 4299 18524
rect 4299 18468 4355 18524
rect 4355 18468 4359 18524
rect 4295 18464 4359 18468
rect 4375 18524 4439 18528
rect 4375 18468 4379 18524
rect 4379 18468 4435 18524
rect 4435 18468 4439 18524
rect 4375 18464 4439 18468
rect 4455 18524 4519 18528
rect 4455 18468 4459 18524
rect 4459 18468 4515 18524
rect 4515 18468 4519 18524
rect 4455 18464 4519 18468
rect 7479 18524 7543 18528
rect 7479 18468 7483 18524
rect 7483 18468 7539 18524
rect 7539 18468 7543 18524
rect 7479 18464 7543 18468
rect 7559 18524 7623 18528
rect 7559 18468 7563 18524
rect 7563 18468 7619 18524
rect 7619 18468 7623 18524
rect 7559 18464 7623 18468
rect 7639 18524 7703 18528
rect 7639 18468 7643 18524
rect 7643 18468 7699 18524
rect 7699 18468 7703 18524
rect 7639 18464 7703 18468
rect 7719 18524 7783 18528
rect 7719 18468 7723 18524
rect 7723 18468 7779 18524
rect 7779 18468 7783 18524
rect 7719 18464 7783 18468
rect 8892 18396 8956 18460
rect 2584 17980 2648 17984
rect 2584 17924 2588 17980
rect 2588 17924 2644 17980
rect 2644 17924 2648 17980
rect 2584 17920 2648 17924
rect 2664 17980 2728 17984
rect 2664 17924 2668 17980
rect 2668 17924 2724 17980
rect 2724 17924 2728 17980
rect 2664 17920 2728 17924
rect 2744 17980 2808 17984
rect 2744 17924 2748 17980
rect 2748 17924 2804 17980
rect 2804 17924 2808 17980
rect 2744 17920 2808 17924
rect 2824 17980 2888 17984
rect 2824 17924 2828 17980
rect 2828 17924 2884 17980
rect 2884 17924 2888 17980
rect 2824 17920 2888 17924
rect 5847 17980 5911 17984
rect 5847 17924 5851 17980
rect 5851 17924 5907 17980
rect 5907 17924 5911 17980
rect 5847 17920 5911 17924
rect 5927 17980 5991 17984
rect 5927 17924 5931 17980
rect 5931 17924 5987 17980
rect 5987 17924 5991 17980
rect 5927 17920 5991 17924
rect 6007 17980 6071 17984
rect 6007 17924 6011 17980
rect 6011 17924 6067 17980
rect 6067 17924 6071 17980
rect 6007 17920 6071 17924
rect 6087 17980 6151 17984
rect 6087 17924 6091 17980
rect 6091 17924 6147 17980
rect 6147 17924 6151 17980
rect 6087 17920 6151 17924
rect 9111 17980 9175 17984
rect 9111 17924 9115 17980
rect 9115 17924 9171 17980
rect 9171 17924 9175 17980
rect 9111 17920 9175 17924
rect 9191 17980 9255 17984
rect 9191 17924 9195 17980
rect 9195 17924 9251 17980
rect 9251 17924 9255 17980
rect 9191 17920 9255 17924
rect 9271 17980 9335 17984
rect 9271 17924 9275 17980
rect 9275 17924 9331 17980
rect 9331 17924 9335 17980
rect 9271 17920 9335 17924
rect 9351 17980 9415 17984
rect 9351 17924 9355 17980
rect 9355 17924 9411 17980
rect 9411 17924 9415 17980
rect 9351 17920 9415 17924
rect 4215 17436 4279 17440
rect 4215 17380 4219 17436
rect 4219 17380 4275 17436
rect 4275 17380 4279 17436
rect 4215 17376 4279 17380
rect 4295 17436 4359 17440
rect 4295 17380 4299 17436
rect 4299 17380 4355 17436
rect 4355 17380 4359 17436
rect 4295 17376 4359 17380
rect 4375 17436 4439 17440
rect 4375 17380 4379 17436
rect 4379 17380 4435 17436
rect 4435 17380 4439 17436
rect 4375 17376 4439 17380
rect 4455 17436 4519 17440
rect 4455 17380 4459 17436
rect 4459 17380 4515 17436
rect 4515 17380 4519 17436
rect 4455 17376 4519 17380
rect 7479 17436 7543 17440
rect 7479 17380 7483 17436
rect 7483 17380 7539 17436
rect 7539 17380 7543 17436
rect 7479 17376 7543 17380
rect 7559 17436 7623 17440
rect 7559 17380 7563 17436
rect 7563 17380 7619 17436
rect 7619 17380 7623 17436
rect 7559 17376 7623 17380
rect 7639 17436 7703 17440
rect 7639 17380 7643 17436
rect 7643 17380 7699 17436
rect 7699 17380 7703 17436
rect 7639 17376 7703 17380
rect 7719 17436 7783 17440
rect 7719 17380 7723 17436
rect 7723 17380 7779 17436
rect 7779 17380 7783 17436
rect 7719 17376 7783 17380
rect 2584 16892 2648 16896
rect 2584 16836 2588 16892
rect 2588 16836 2644 16892
rect 2644 16836 2648 16892
rect 2584 16832 2648 16836
rect 2664 16892 2728 16896
rect 2664 16836 2668 16892
rect 2668 16836 2724 16892
rect 2724 16836 2728 16892
rect 2664 16832 2728 16836
rect 2744 16892 2808 16896
rect 2744 16836 2748 16892
rect 2748 16836 2804 16892
rect 2804 16836 2808 16892
rect 2744 16832 2808 16836
rect 2824 16892 2888 16896
rect 2824 16836 2828 16892
rect 2828 16836 2884 16892
rect 2884 16836 2888 16892
rect 2824 16832 2888 16836
rect 5847 16892 5911 16896
rect 5847 16836 5851 16892
rect 5851 16836 5907 16892
rect 5907 16836 5911 16892
rect 5847 16832 5911 16836
rect 5927 16892 5991 16896
rect 5927 16836 5931 16892
rect 5931 16836 5987 16892
rect 5987 16836 5991 16892
rect 5927 16832 5991 16836
rect 6007 16892 6071 16896
rect 6007 16836 6011 16892
rect 6011 16836 6067 16892
rect 6067 16836 6071 16892
rect 6007 16832 6071 16836
rect 6087 16892 6151 16896
rect 6087 16836 6091 16892
rect 6091 16836 6147 16892
rect 6147 16836 6151 16892
rect 6087 16832 6151 16836
rect 9111 16892 9175 16896
rect 9111 16836 9115 16892
rect 9115 16836 9171 16892
rect 9171 16836 9175 16892
rect 9111 16832 9175 16836
rect 9191 16892 9255 16896
rect 9191 16836 9195 16892
rect 9195 16836 9251 16892
rect 9251 16836 9255 16892
rect 9191 16832 9255 16836
rect 9271 16892 9335 16896
rect 9271 16836 9275 16892
rect 9275 16836 9331 16892
rect 9331 16836 9335 16892
rect 9271 16832 9335 16836
rect 9351 16892 9415 16896
rect 9351 16836 9355 16892
rect 9355 16836 9411 16892
rect 9411 16836 9415 16892
rect 9351 16832 9415 16836
rect 4215 16348 4279 16352
rect 4215 16292 4219 16348
rect 4219 16292 4275 16348
rect 4275 16292 4279 16348
rect 4215 16288 4279 16292
rect 4295 16348 4359 16352
rect 4295 16292 4299 16348
rect 4299 16292 4355 16348
rect 4355 16292 4359 16348
rect 4295 16288 4359 16292
rect 4375 16348 4439 16352
rect 4375 16292 4379 16348
rect 4379 16292 4435 16348
rect 4435 16292 4439 16348
rect 4375 16288 4439 16292
rect 4455 16348 4519 16352
rect 4455 16292 4459 16348
rect 4459 16292 4515 16348
rect 4515 16292 4519 16348
rect 4455 16288 4519 16292
rect 7479 16348 7543 16352
rect 7479 16292 7483 16348
rect 7483 16292 7539 16348
rect 7539 16292 7543 16348
rect 7479 16288 7543 16292
rect 7559 16348 7623 16352
rect 7559 16292 7563 16348
rect 7563 16292 7619 16348
rect 7619 16292 7623 16348
rect 7559 16288 7623 16292
rect 7639 16348 7703 16352
rect 7639 16292 7643 16348
rect 7643 16292 7699 16348
rect 7699 16292 7703 16348
rect 7639 16288 7703 16292
rect 7719 16348 7783 16352
rect 7719 16292 7723 16348
rect 7723 16292 7779 16348
rect 7779 16292 7783 16348
rect 7719 16288 7783 16292
rect 2584 15804 2648 15808
rect 2584 15748 2588 15804
rect 2588 15748 2644 15804
rect 2644 15748 2648 15804
rect 2584 15744 2648 15748
rect 2664 15804 2728 15808
rect 2664 15748 2668 15804
rect 2668 15748 2724 15804
rect 2724 15748 2728 15804
rect 2664 15744 2728 15748
rect 2744 15804 2808 15808
rect 2744 15748 2748 15804
rect 2748 15748 2804 15804
rect 2804 15748 2808 15804
rect 2744 15744 2808 15748
rect 2824 15804 2888 15808
rect 2824 15748 2828 15804
rect 2828 15748 2884 15804
rect 2884 15748 2888 15804
rect 2824 15744 2888 15748
rect 5847 15804 5911 15808
rect 5847 15748 5851 15804
rect 5851 15748 5907 15804
rect 5907 15748 5911 15804
rect 5847 15744 5911 15748
rect 5927 15804 5991 15808
rect 5927 15748 5931 15804
rect 5931 15748 5987 15804
rect 5987 15748 5991 15804
rect 5927 15744 5991 15748
rect 6007 15804 6071 15808
rect 6007 15748 6011 15804
rect 6011 15748 6067 15804
rect 6067 15748 6071 15804
rect 6007 15744 6071 15748
rect 6087 15804 6151 15808
rect 6087 15748 6091 15804
rect 6091 15748 6147 15804
rect 6147 15748 6151 15804
rect 6087 15744 6151 15748
rect 9111 15804 9175 15808
rect 9111 15748 9115 15804
rect 9115 15748 9171 15804
rect 9171 15748 9175 15804
rect 9111 15744 9175 15748
rect 9191 15804 9255 15808
rect 9191 15748 9195 15804
rect 9195 15748 9251 15804
rect 9251 15748 9255 15804
rect 9191 15744 9255 15748
rect 9271 15804 9335 15808
rect 9271 15748 9275 15804
rect 9275 15748 9331 15804
rect 9331 15748 9335 15804
rect 9271 15744 9335 15748
rect 9351 15804 9415 15808
rect 9351 15748 9355 15804
rect 9355 15748 9411 15804
rect 9411 15748 9415 15804
rect 9351 15744 9415 15748
rect 4215 15260 4279 15264
rect 4215 15204 4219 15260
rect 4219 15204 4275 15260
rect 4275 15204 4279 15260
rect 4215 15200 4279 15204
rect 4295 15260 4359 15264
rect 4295 15204 4299 15260
rect 4299 15204 4355 15260
rect 4355 15204 4359 15260
rect 4295 15200 4359 15204
rect 4375 15260 4439 15264
rect 4375 15204 4379 15260
rect 4379 15204 4435 15260
rect 4435 15204 4439 15260
rect 4375 15200 4439 15204
rect 4455 15260 4519 15264
rect 4455 15204 4459 15260
rect 4459 15204 4515 15260
rect 4515 15204 4519 15260
rect 4455 15200 4519 15204
rect 7479 15260 7543 15264
rect 7479 15204 7483 15260
rect 7483 15204 7539 15260
rect 7539 15204 7543 15260
rect 7479 15200 7543 15204
rect 7559 15260 7623 15264
rect 7559 15204 7563 15260
rect 7563 15204 7619 15260
rect 7619 15204 7623 15260
rect 7559 15200 7623 15204
rect 7639 15260 7703 15264
rect 7639 15204 7643 15260
rect 7643 15204 7699 15260
rect 7699 15204 7703 15260
rect 7639 15200 7703 15204
rect 7719 15260 7783 15264
rect 7719 15204 7723 15260
rect 7723 15204 7779 15260
rect 7779 15204 7783 15260
rect 7719 15200 7783 15204
rect 2584 14716 2648 14720
rect 2584 14660 2588 14716
rect 2588 14660 2644 14716
rect 2644 14660 2648 14716
rect 2584 14656 2648 14660
rect 2664 14716 2728 14720
rect 2664 14660 2668 14716
rect 2668 14660 2724 14716
rect 2724 14660 2728 14716
rect 2664 14656 2728 14660
rect 2744 14716 2808 14720
rect 2744 14660 2748 14716
rect 2748 14660 2804 14716
rect 2804 14660 2808 14716
rect 2744 14656 2808 14660
rect 2824 14716 2888 14720
rect 2824 14660 2828 14716
rect 2828 14660 2884 14716
rect 2884 14660 2888 14716
rect 2824 14656 2888 14660
rect 5847 14716 5911 14720
rect 5847 14660 5851 14716
rect 5851 14660 5907 14716
rect 5907 14660 5911 14716
rect 5847 14656 5911 14660
rect 5927 14716 5991 14720
rect 5927 14660 5931 14716
rect 5931 14660 5987 14716
rect 5987 14660 5991 14716
rect 5927 14656 5991 14660
rect 6007 14716 6071 14720
rect 6007 14660 6011 14716
rect 6011 14660 6067 14716
rect 6067 14660 6071 14716
rect 6007 14656 6071 14660
rect 6087 14716 6151 14720
rect 6087 14660 6091 14716
rect 6091 14660 6147 14716
rect 6147 14660 6151 14716
rect 6087 14656 6151 14660
rect 9111 14716 9175 14720
rect 9111 14660 9115 14716
rect 9115 14660 9171 14716
rect 9171 14660 9175 14716
rect 9111 14656 9175 14660
rect 9191 14716 9255 14720
rect 9191 14660 9195 14716
rect 9195 14660 9251 14716
rect 9251 14660 9255 14716
rect 9191 14656 9255 14660
rect 9271 14716 9335 14720
rect 9271 14660 9275 14716
rect 9275 14660 9331 14716
rect 9331 14660 9335 14716
rect 9271 14656 9335 14660
rect 9351 14716 9415 14720
rect 9351 14660 9355 14716
rect 9355 14660 9411 14716
rect 9411 14660 9415 14716
rect 9351 14656 9415 14660
rect 7236 14648 7300 14652
rect 7236 14592 7286 14648
rect 7286 14592 7300 14648
rect 7236 14588 7300 14592
rect 4215 14172 4279 14176
rect 4215 14116 4219 14172
rect 4219 14116 4275 14172
rect 4275 14116 4279 14172
rect 4215 14112 4279 14116
rect 4295 14172 4359 14176
rect 4295 14116 4299 14172
rect 4299 14116 4355 14172
rect 4355 14116 4359 14172
rect 4295 14112 4359 14116
rect 4375 14172 4439 14176
rect 4375 14116 4379 14172
rect 4379 14116 4435 14172
rect 4435 14116 4439 14172
rect 4375 14112 4439 14116
rect 4455 14172 4519 14176
rect 4455 14116 4459 14172
rect 4459 14116 4515 14172
rect 4515 14116 4519 14172
rect 4455 14112 4519 14116
rect 7479 14172 7543 14176
rect 7479 14116 7483 14172
rect 7483 14116 7539 14172
rect 7539 14116 7543 14172
rect 7479 14112 7543 14116
rect 7559 14172 7623 14176
rect 7559 14116 7563 14172
rect 7563 14116 7619 14172
rect 7619 14116 7623 14172
rect 7559 14112 7623 14116
rect 7639 14172 7703 14176
rect 7639 14116 7643 14172
rect 7643 14116 7699 14172
rect 7699 14116 7703 14172
rect 7639 14112 7703 14116
rect 7719 14172 7783 14176
rect 7719 14116 7723 14172
rect 7723 14116 7779 14172
rect 7779 14116 7783 14172
rect 7719 14112 7783 14116
rect 2584 13628 2648 13632
rect 2584 13572 2588 13628
rect 2588 13572 2644 13628
rect 2644 13572 2648 13628
rect 2584 13568 2648 13572
rect 2664 13628 2728 13632
rect 2664 13572 2668 13628
rect 2668 13572 2724 13628
rect 2724 13572 2728 13628
rect 2664 13568 2728 13572
rect 2744 13628 2808 13632
rect 2744 13572 2748 13628
rect 2748 13572 2804 13628
rect 2804 13572 2808 13628
rect 2744 13568 2808 13572
rect 2824 13628 2888 13632
rect 2824 13572 2828 13628
rect 2828 13572 2884 13628
rect 2884 13572 2888 13628
rect 2824 13568 2888 13572
rect 5847 13628 5911 13632
rect 5847 13572 5851 13628
rect 5851 13572 5907 13628
rect 5907 13572 5911 13628
rect 5847 13568 5911 13572
rect 5927 13628 5991 13632
rect 5927 13572 5931 13628
rect 5931 13572 5987 13628
rect 5987 13572 5991 13628
rect 5927 13568 5991 13572
rect 6007 13628 6071 13632
rect 6007 13572 6011 13628
rect 6011 13572 6067 13628
rect 6067 13572 6071 13628
rect 6007 13568 6071 13572
rect 6087 13628 6151 13632
rect 6087 13572 6091 13628
rect 6091 13572 6147 13628
rect 6147 13572 6151 13628
rect 6087 13568 6151 13572
rect 9111 13628 9175 13632
rect 9111 13572 9115 13628
rect 9115 13572 9171 13628
rect 9171 13572 9175 13628
rect 9111 13568 9175 13572
rect 9191 13628 9255 13632
rect 9191 13572 9195 13628
rect 9195 13572 9251 13628
rect 9251 13572 9255 13628
rect 9191 13568 9255 13572
rect 9271 13628 9335 13632
rect 9271 13572 9275 13628
rect 9275 13572 9331 13628
rect 9331 13572 9335 13628
rect 9271 13568 9335 13572
rect 9351 13628 9415 13632
rect 9351 13572 9355 13628
rect 9355 13572 9411 13628
rect 9411 13572 9415 13628
rect 9351 13568 9415 13572
rect 7236 13500 7300 13564
rect 4215 13084 4279 13088
rect 4215 13028 4219 13084
rect 4219 13028 4275 13084
rect 4275 13028 4279 13084
rect 4215 13024 4279 13028
rect 4295 13084 4359 13088
rect 4295 13028 4299 13084
rect 4299 13028 4355 13084
rect 4355 13028 4359 13084
rect 4295 13024 4359 13028
rect 4375 13084 4439 13088
rect 4375 13028 4379 13084
rect 4379 13028 4435 13084
rect 4435 13028 4439 13084
rect 4375 13024 4439 13028
rect 4455 13084 4519 13088
rect 4455 13028 4459 13084
rect 4459 13028 4515 13084
rect 4515 13028 4519 13084
rect 4455 13024 4519 13028
rect 7479 13084 7543 13088
rect 7479 13028 7483 13084
rect 7483 13028 7539 13084
rect 7539 13028 7543 13084
rect 7479 13024 7543 13028
rect 7559 13084 7623 13088
rect 7559 13028 7563 13084
rect 7563 13028 7619 13084
rect 7619 13028 7623 13084
rect 7559 13024 7623 13028
rect 7639 13084 7703 13088
rect 7639 13028 7643 13084
rect 7643 13028 7699 13084
rect 7699 13028 7703 13084
rect 7639 13024 7703 13028
rect 7719 13084 7783 13088
rect 7719 13028 7723 13084
rect 7723 13028 7779 13084
rect 7779 13028 7783 13084
rect 7719 13024 7783 13028
rect 2584 12540 2648 12544
rect 2584 12484 2588 12540
rect 2588 12484 2644 12540
rect 2644 12484 2648 12540
rect 2584 12480 2648 12484
rect 2664 12540 2728 12544
rect 2664 12484 2668 12540
rect 2668 12484 2724 12540
rect 2724 12484 2728 12540
rect 2664 12480 2728 12484
rect 2744 12540 2808 12544
rect 2744 12484 2748 12540
rect 2748 12484 2804 12540
rect 2804 12484 2808 12540
rect 2744 12480 2808 12484
rect 2824 12540 2888 12544
rect 2824 12484 2828 12540
rect 2828 12484 2884 12540
rect 2884 12484 2888 12540
rect 2824 12480 2888 12484
rect 5847 12540 5911 12544
rect 5847 12484 5851 12540
rect 5851 12484 5907 12540
rect 5907 12484 5911 12540
rect 5847 12480 5911 12484
rect 5927 12540 5991 12544
rect 5927 12484 5931 12540
rect 5931 12484 5987 12540
rect 5987 12484 5991 12540
rect 5927 12480 5991 12484
rect 6007 12540 6071 12544
rect 6007 12484 6011 12540
rect 6011 12484 6067 12540
rect 6067 12484 6071 12540
rect 6007 12480 6071 12484
rect 6087 12540 6151 12544
rect 6087 12484 6091 12540
rect 6091 12484 6147 12540
rect 6147 12484 6151 12540
rect 6087 12480 6151 12484
rect 9111 12540 9175 12544
rect 9111 12484 9115 12540
rect 9115 12484 9171 12540
rect 9171 12484 9175 12540
rect 9111 12480 9175 12484
rect 9191 12540 9255 12544
rect 9191 12484 9195 12540
rect 9195 12484 9251 12540
rect 9251 12484 9255 12540
rect 9191 12480 9255 12484
rect 9271 12540 9335 12544
rect 9271 12484 9275 12540
rect 9275 12484 9331 12540
rect 9331 12484 9335 12540
rect 9271 12480 9335 12484
rect 9351 12540 9415 12544
rect 9351 12484 9355 12540
rect 9355 12484 9411 12540
rect 9411 12484 9415 12540
rect 9351 12480 9415 12484
rect 4215 11996 4279 12000
rect 4215 11940 4219 11996
rect 4219 11940 4275 11996
rect 4275 11940 4279 11996
rect 4215 11936 4279 11940
rect 4295 11996 4359 12000
rect 4295 11940 4299 11996
rect 4299 11940 4355 11996
rect 4355 11940 4359 11996
rect 4295 11936 4359 11940
rect 4375 11996 4439 12000
rect 4375 11940 4379 11996
rect 4379 11940 4435 11996
rect 4435 11940 4439 11996
rect 4375 11936 4439 11940
rect 4455 11996 4519 12000
rect 4455 11940 4459 11996
rect 4459 11940 4515 11996
rect 4515 11940 4519 11996
rect 4455 11936 4519 11940
rect 7479 11996 7543 12000
rect 7479 11940 7483 11996
rect 7483 11940 7539 11996
rect 7539 11940 7543 11996
rect 7479 11936 7543 11940
rect 7559 11996 7623 12000
rect 7559 11940 7563 11996
rect 7563 11940 7619 11996
rect 7619 11940 7623 11996
rect 7559 11936 7623 11940
rect 7639 11996 7703 12000
rect 7639 11940 7643 11996
rect 7643 11940 7699 11996
rect 7699 11940 7703 11996
rect 7639 11936 7703 11940
rect 7719 11996 7783 12000
rect 7719 11940 7723 11996
rect 7723 11940 7779 11996
rect 7779 11940 7783 11996
rect 7719 11936 7783 11940
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5847 11452 5911 11456
rect 5847 11396 5851 11452
rect 5851 11396 5907 11452
rect 5907 11396 5911 11452
rect 5847 11392 5911 11396
rect 5927 11452 5991 11456
rect 5927 11396 5931 11452
rect 5931 11396 5987 11452
rect 5987 11396 5991 11452
rect 5927 11392 5991 11396
rect 6007 11452 6071 11456
rect 6007 11396 6011 11452
rect 6011 11396 6067 11452
rect 6067 11396 6071 11452
rect 6007 11392 6071 11396
rect 6087 11452 6151 11456
rect 6087 11396 6091 11452
rect 6091 11396 6147 11452
rect 6147 11396 6151 11452
rect 6087 11392 6151 11396
rect 9111 11452 9175 11456
rect 9111 11396 9115 11452
rect 9115 11396 9171 11452
rect 9171 11396 9175 11452
rect 9111 11392 9175 11396
rect 9191 11452 9255 11456
rect 9191 11396 9195 11452
rect 9195 11396 9251 11452
rect 9251 11396 9255 11452
rect 9191 11392 9255 11396
rect 9271 11452 9335 11456
rect 9271 11396 9275 11452
rect 9275 11396 9331 11452
rect 9331 11396 9335 11452
rect 9271 11392 9335 11396
rect 9351 11452 9415 11456
rect 9351 11396 9355 11452
rect 9355 11396 9411 11452
rect 9411 11396 9415 11452
rect 9351 11392 9415 11396
rect 4215 10908 4279 10912
rect 4215 10852 4219 10908
rect 4219 10852 4275 10908
rect 4275 10852 4279 10908
rect 4215 10848 4279 10852
rect 4295 10908 4359 10912
rect 4295 10852 4299 10908
rect 4299 10852 4355 10908
rect 4355 10852 4359 10908
rect 4295 10848 4359 10852
rect 4375 10908 4439 10912
rect 4375 10852 4379 10908
rect 4379 10852 4435 10908
rect 4435 10852 4439 10908
rect 4375 10848 4439 10852
rect 4455 10908 4519 10912
rect 4455 10852 4459 10908
rect 4459 10852 4515 10908
rect 4515 10852 4519 10908
rect 4455 10848 4519 10852
rect 7479 10908 7543 10912
rect 7479 10852 7483 10908
rect 7483 10852 7539 10908
rect 7539 10852 7543 10908
rect 7479 10848 7543 10852
rect 7559 10908 7623 10912
rect 7559 10852 7563 10908
rect 7563 10852 7619 10908
rect 7619 10852 7623 10908
rect 7559 10848 7623 10852
rect 7639 10908 7703 10912
rect 7639 10852 7643 10908
rect 7643 10852 7699 10908
rect 7699 10852 7703 10908
rect 7639 10848 7703 10852
rect 7719 10908 7783 10912
rect 7719 10852 7723 10908
rect 7723 10852 7779 10908
rect 7779 10852 7783 10908
rect 7719 10848 7783 10852
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5847 10364 5911 10368
rect 5847 10308 5851 10364
rect 5851 10308 5907 10364
rect 5907 10308 5911 10364
rect 5847 10304 5911 10308
rect 5927 10364 5991 10368
rect 5927 10308 5931 10364
rect 5931 10308 5987 10364
rect 5987 10308 5991 10364
rect 5927 10304 5991 10308
rect 6007 10364 6071 10368
rect 6007 10308 6011 10364
rect 6011 10308 6067 10364
rect 6067 10308 6071 10364
rect 6007 10304 6071 10308
rect 6087 10364 6151 10368
rect 6087 10308 6091 10364
rect 6091 10308 6147 10364
rect 6147 10308 6151 10364
rect 6087 10304 6151 10308
rect 9111 10364 9175 10368
rect 9111 10308 9115 10364
rect 9115 10308 9171 10364
rect 9171 10308 9175 10364
rect 9111 10304 9175 10308
rect 9191 10364 9255 10368
rect 9191 10308 9195 10364
rect 9195 10308 9251 10364
rect 9251 10308 9255 10364
rect 9191 10304 9255 10308
rect 9271 10364 9335 10368
rect 9271 10308 9275 10364
rect 9275 10308 9331 10364
rect 9331 10308 9335 10364
rect 9271 10304 9335 10308
rect 9351 10364 9415 10368
rect 9351 10308 9355 10364
rect 9355 10308 9411 10364
rect 9411 10308 9415 10364
rect 9351 10304 9415 10308
rect 8892 10100 8956 10164
rect 4215 9820 4279 9824
rect 4215 9764 4219 9820
rect 4219 9764 4275 9820
rect 4275 9764 4279 9820
rect 4215 9760 4279 9764
rect 4295 9820 4359 9824
rect 4295 9764 4299 9820
rect 4299 9764 4355 9820
rect 4355 9764 4359 9820
rect 4295 9760 4359 9764
rect 4375 9820 4439 9824
rect 4375 9764 4379 9820
rect 4379 9764 4435 9820
rect 4435 9764 4439 9820
rect 4375 9760 4439 9764
rect 4455 9820 4519 9824
rect 4455 9764 4459 9820
rect 4459 9764 4515 9820
rect 4515 9764 4519 9820
rect 4455 9760 4519 9764
rect 7479 9820 7543 9824
rect 7479 9764 7483 9820
rect 7483 9764 7539 9820
rect 7539 9764 7543 9820
rect 7479 9760 7543 9764
rect 7559 9820 7623 9824
rect 7559 9764 7563 9820
rect 7563 9764 7619 9820
rect 7619 9764 7623 9820
rect 7559 9760 7623 9764
rect 7639 9820 7703 9824
rect 7639 9764 7643 9820
rect 7643 9764 7699 9820
rect 7699 9764 7703 9820
rect 7639 9760 7703 9764
rect 7719 9820 7783 9824
rect 7719 9764 7723 9820
rect 7723 9764 7779 9820
rect 7779 9764 7783 9820
rect 7719 9760 7783 9764
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5847 9276 5911 9280
rect 5847 9220 5851 9276
rect 5851 9220 5907 9276
rect 5907 9220 5911 9276
rect 5847 9216 5911 9220
rect 5927 9276 5991 9280
rect 5927 9220 5931 9276
rect 5931 9220 5987 9276
rect 5987 9220 5991 9276
rect 5927 9216 5991 9220
rect 6007 9276 6071 9280
rect 6007 9220 6011 9276
rect 6011 9220 6067 9276
rect 6067 9220 6071 9276
rect 6007 9216 6071 9220
rect 6087 9276 6151 9280
rect 6087 9220 6091 9276
rect 6091 9220 6147 9276
rect 6147 9220 6151 9276
rect 6087 9216 6151 9220
rect 9111 9276 9175 9280
rect 9111 9220 9115 9276
rect 9115 9220 9171 9276
rect 9171 9220 9175 9276
rect 9111 9216 9175 9220
rect 9191 9276 9255 9280
rect 9191 9220 9195 9276
rect 9195 9220 9251 9276
rect 9251 9220 9255 9276
rect 9191 9216 9255 9220
rect 9271 9276 9335 9280
rect 9271 9220 9275 9276
rect 9275 9220 9331 9276
rect 9331 9220 9335 9276
rect 9271 9216 9335 9220
rect 9351 9276 9415 9280
rect 9351 9220 9355 9276
rect 9355 9220 9411 9276
rect 9411 9220 9415 9276
rect 9351 9216 9415 9220
rect 4215 8732 4279 8736
rect 4215 8676 4219 8732
rect 4219 8676 4275 8732
rect 4275 8676 4279 8732
rect 4215 8672 4279 8676
rect 4295 8732 4359 8736
rect 4295 8676 4299 8732
rect 4299 8676 4355 8732
rect 4355 8676 4359 8732
rect 4295 8672 4359 8676
rect 4375 8732 4439 8736
rect 4375 8676 4379 8732
rect 4379 8676 4435 8732
rect 4435 8676 4439 8732
rect 4375 8672 4439 8676
rect 4455 8732 4519 8736
rect 4455 8676 4459 8732
rect 4459 8676 4515 8732
rect 4515 8676 4519 8732
rect 4455 8672 4519 8676
rect 7479 8732 7543 8736
rect 7479 8676 7483 8732
rect 7483 8676 7539 8732
rect 7539 8676 7543 8732
rect 7479 8672 7543 8676
rect 7559 8732 7623 8736
rect 7559 8676 7563 8732
rect 7563 8676 7619 8732
rect 7619 8676 7623 8732
rect 7559 8672 7623 8676
rect 7639 8732 7703 8736
rect 7639 8676 7643 8732
rect 7643 8676 7699 8732
rect 7699 8676 7703 8732
rect 7639 8672 7703 8676
rect 7719 8732 7783 8736
rect 7719 8676 7723 8732
rect 7723 8676 7779 8732
rect 7779 8676 7783 8732
rect 7719 8672 7783 8676
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5847 8188 5911 8192
rect 5847 8132 5851 8188
rect 5851 8132 5907 8188
rect 5907 8132 5911 8188
rect 5847 8128 5911 8132
rect 5927 8188 5991 8192
rect 5927 8132 5931 8188
rect 5931 8132 5987 8188
rect 5987 8132 5991 8188
rect 5927 8128 5991 8132
rect 6007 8188 6071 8192
rect 6007 8132 6011 8188
rect 6011 8132 6067 8188
rect 6067 8132 6071 8188
rect 6007 8128 6071 8132
rect 6087 8188 6151 8192
rect 6087 8132 6091 8188
rect 6091 8132 6147 8188
rect 6147 8132 6151 8188
rect 6087 8128 6151 8132
rect 9111 8188 9175 8192
rect 9111 8132 9115 8188
rect 9115 8132 9171 8188
rect 9171 8132 9175 8188
rect 9111 8128 9175 8132
rect 9191 8188 9255 8192
rect 9191 8132 9195 8188
rect 9195 8132 9251 8188
rect 9251 8132 9255 8188
rect 9191 8128 9255 8132
rect 9271 8188 9335 8192
rect 9271 8132 9275 8188
rect 9275 8132 9331 8188
rect 9331 8132 9335 8188
rect 9271 8128 9335 8132
rect 9351 8188 9415 8192
rect 9351 8132 9355 8188
rect 9355 8132 9411 8188
rect 9411 8132 9415 8188
rect 9351 8128 9415 8132
rect 4215 7644 4279 7648
rect 4215 7588 4219 7644
rect 4219 7588 4275 7644
rect 4275 7588 4279 7644
rect 4215 7584 4279 7588
rect 4295 7644 4359 7648
rect 4295 7588 4299 7644
rect 4299 7588 4355 7644
rect 4355 7588 4359 7644
rect 4295 7584 4359 7588
rect 4375 7644 4439 7648
rect 4375 7588 4379 7644
rect 4379 7588 4435 7644
rect 4435 7588 4439 7644
rect 4375 7584 4439 7588
rect 4455 7644 4519 7648
rect 4455 7588 4459 7644
rect 4459 7588 4515 7644
rect 4515 7588 4519 7644
rect 4455 7584 4519 7588
rect 7479 7644 7543 7648
rect 7479 7588 7483 7644
rect 7483 7588 7539 7644
rect 7539 7588 7543 7644
rect 7479 7584 7543 7588
rect 7559 7644 7623 7648
rect 7559 7588 7563 7644
rect 7563 7588 7619 7644
rect 7619 7588 7623 7644
rect 7559 7584 7623 7588
rect 7639 7644 7703 7648
rect 7639 7588 7643 7644
rect 7643 7588 7699 7644
rect 7699 7588 7703 7644
rect 7639 7584 7703 7588
rect 7719 7644 7783 7648
rect 7719 7588 7723 7644
rect 7723 7588 7779 7644
rect 7779 7588 7783 7644
rect 7719 7584 7783 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5847 7100 5911 7104
rect 5847 7044 5851 7100
rect 5851 7044 5907 7100
rect 5907 7044 5911 7100
rect 5847 7040 5911 7044
rect 5927 7100 5991 7104
rect 5927 7044 5931 7100
rect 5931 7044 5987 7100
rect 5987 7044 5991 7100
rect 5927 7040 5991 7044
rect 6007 7100 6071 7104
rect 6007 7044 6011 7100
rect 6011 7044 6067 7100
rect 6067 7044 6071 7100
rect 6007 7040 6071 7044
rect 6087 7100 6151 7104
rect 6087 7044 6091 7100
rect 6091 7044 6147 7100
rect 6147 7044 6151 7100
rect 6087 7040 6151 7044
rect 9111 7100 9175 7104
rect 9111 7044 9115 7100
rect 9115 7044 9171 7100
rect 9171 7044 9175 7100
rect 9111 7040 9175 7044
rect 9191 7100 9255 7104
rect 9191 7044 9195 7100
rect 9195 7044 9251 7100
rect 9251 7044 9255 7100
rect 9191 7040 9255 7044
rect 9271 7100 9335 7104
rect 9271 7044 9275 7100
rect 9275 7044 9331 7100
rect 9331 7044 9335 7100
rect 9271 7040 9335 7044
rect 9351 7100 9415 7104
rect 9351 7044 9355 7100
rect 9355 7044 9411 7100
rect 9411 7044 9415 7100
rect 9351 7040 9415 7044
rect 4215 6556 4279 6560
rect 4215 6500 4219 6556
rect 4219 6500 4275 6556
rect 4275 6500 4279 6556
rect 4215 6496 4279 6500
rect 4295 6556 4359 6560
rect 4295 6500 4299 6556
rect 4299 6500 4355 6556
rect 4355 6500 4359 6556
rect 4295 6496 4359 6500
rect 4375 6556 4439 6560
rect 4375 6500 4379 6556
rect 4379 6500 4435 6556
rect 4435 6500 4439 6556
rect 4375 6496 4439 6500
rect 4455 6556 4519 6560
rect 4455 6500 4459 6556
rect 4459 6500 4515 6556
rect 4515 6500 4519 6556
rect 4455 6496 4519 6500
rect 7479 6556 7543 6560
rect 7479 6500 7483 6556
rect 7483 6500 7539 6556
rect 7539 6500 7543 6556
rect 7479 6496 7543 6500
rect 7559 6556 7623 6560
rect 7559 6500 7563 6556
rect 7563 6500 7619 6556
rect 7619 6500 7623 6556
rect 7559 6496 7623 6500
rect 7639 6556 7703 6560
rect 7639 6500 7643 6556
rect 7643 6500 7699 6556
rect 7699 6500 7703 6556
rect 7639 6496 7703 6500
rect 7719 6556 7783 6560
rect 7719 6500 7723 6556
rect 7723 6500 7779 6556
rect 7779 6500 7783 6556
rect 7719 6496 7783 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5847 6012 5911 6016
rect 5847 5956 5851 6012
rect 5851 5956 5907 6012
rect 5907 5956 5911 6012
rect 5847 5952 5911 5956
rect 5927 6012 5991 6016
rect 5927 5956 5931 6012
rect 5931 5956 5987 6012
rect 5987 5956 5991 6012
rect 5927 5952 5991 5956
rect 6007 6012 6071 6016
rect 6007 5956 6011 6012
rect 6011 5956 6067 6012
rect 6067 5956 6071 6012
rect 6007 5952 6071 5956
rect 6087 6012 6151 6016
rect 6087 5956 6091 6012
rect 6091 5956 6147 6012
rect 6147 5956 6151 6012
rect 6087 5952 6151 5956
rect 9111 6012 9175 6016
rect 9111 5956 9115 6012
rect 9115 5956 9171 6012
rect 9171 5956 9175 6012
rect 9111 5952 9175 5956
rect 9191 6012 9255 6016
rect 9191 5956 9195 6012
rect 9195 5956 9251 6012
rect 9251 5956 9255 6012
rect 9191 5952 9255 5956
rect 9271 6012 9335 6016
rect 9271 5956 9275 6012
rect 9275 5956 9331 6012
rect 9331 5956 9335 6012
rect 9271 5952 9335 5956
rect 9351 6012 9415 6016
rect 9351 5956 9355 6012
rect 9355 5956 9411 6012
rect 9411 5956 9415 6012
rect 9351 5952 9415 5956
rect 4215 5468 4279 5472
rect 4215 5412 4219 5468
rect 4219 5412 4275 5468
rect 4275 5412 4279 5468
rect 4215 5408 4279 5412
rect 4295 5468 4359 5472
rect 4295 5412 4299 5468
rect 4299 5412 4355 5468
rect 4355 5412 4359 5468
rect 4295 5408 4359 5412
rect 4375 5468 4439 5472
rect 4375 5412 4379 5468
rect 4379 5412 4435 5468
rect 4435 5412 4439 5468
rect 4375 5408 4439 5412
rect 4455 5468 4519 5472
rect 4455 5412 4459 5468
rect 4459 5412 4515 5468
rect 4515 5412 4519 5468
rect 4455 5408 4519 5412
rect 7479 5468 7543 5472
rect 7479 5412 7483 5468
rect 7483 5412 7539 5468
rect 7539 5412 7543 5468
rect 7479 5408 7543 5412
rect 7559 5468 7623 5472
rect 7559 5412 7563 5468
rect 7563 5412 7619 5468
rect 7619 5412 7623 5468
rect 7559 5408 7623 5412
rect 7639 5468 7703 5472
rect 7639 5412 7643 5468
rect 7643 5412 7699 5468
rect 7699 5412 7703 5468
rect 7639 5408 7703 5412
rect 7719 5468 7783 5472
rect 7719 5412 7723 5468
rect 7723 5412 7779 5468
rect 7779 5412 7783 5468
rect 7719 5408 7783 5412
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5847 4924 5911 4928
rect 5847 4868 5851 4924
rect 5851 4868 5907 4924
rect 5907 4868 5911 4924
rect 5847 4864 5911 4868
rect 5927 4924 5991 4928
rect 5927 4868 5931 4924
rect 5931 4868 5987 4924
rect 5987 4868 5991 4924
rect 5927 4864 5991 4868
rect 6007 4924 6071 4928
rect 6007 4868 6011 4924
rect 6011 4868 6067 4924
rect 6067 4868 6071 4924
rect 6007 4864 6071 4868
rect 6087 4924 6151 4928
rect 6087 4868 6091 4924
rect 6091 4868 6147 4924
rect 6147 4868 6151 4924
rect 6087 4864 6151 4868
rect 9111 4924 9175 4928
rect 9111 4868 9115 4924
rect 9115 4868 9171 4924
rect 9171 4868 9175 4924
rect 9111 4864 9175 4868
rect 9191 4924 9255 4928
rect 9191 4868 9195 4924
rect 9195 4868 9251 4924
rect 9251 4868 9255 4924
rect 9191 4864 9255 4868
rect 9271 4924 9335 4928
rect 9271 4868 9275 4924
rect 9275 4868 9331 4924
rect 9331 4868 9335 4924
rect 9271 4864 9335 4868
rect 9351 4924 9415 4928
rect 9351 4868 9355 4924
rect 9355 4868 9411 4924
rect 9411 4868 9415 4924
rect 9351 4864 9415 4868
rect 4215 4380 4279 4384
rect 4215 4324 4219 4380
rect 4219 4324 4275 4380
rect 4275 4324 4279 4380
rect 4215 4320 4279 4324
rect 4295 4380 4359 4384
rect 4295 4324 4299 4380
rect 4299 4324 4355 4380
rect 4355 4324 4359 4380
rect 4295 4320 4359 4324
rect 4375 4380 4439 4384
rect 4375 4324 4379 4380
rect 4379 4324 4435 4380
rect 4435 4324 4439 4380
rect 4375 4320 4439 4324
rect 4455 4380 4519 4384
rect 4455 4324 4459 4380
rect 4459 4324 4515 4380
rect 4515 4324 4519 4380
rect 4455 4320 4519 4324
rect 7479 4380 7543 4384
rect 7479 4324 7483 4380
rect 7483 4324 7539 4380
rect 7539 4324 7543 4380
rect 7479 4320 7543 4324
rect 7559 4380 7623 4384
rect 7559 4324 7563 4380
rect 7563 4324 7619 4380
rect 7619 4324 7623 4380
rect 7559 4320 7623 4324
rect 7639 4380 7703 4384
rect 7639 4324 7643 4380
rect 7643 4324 7699 4380
rect 7699 4324 7703 4380
rect 7639 4320 7703 4324
rect 7719 4380 7783 4384
rect 7719 4324 7723 4380
rect 7723 4324 7779 4380
rect 7779 4324 7783 4380
rect 7719 4320 7783 4324
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5847 3836 5911 3840
rect 5847 3780 5851 3836
rect 5851 3780 5907 3836
rect 5907 3780 5911 3836
rect 5847 3776 5911 3780
rect 5927 3836 5991 3840
rect 5927 3780 5931 3836
rect 5931 3780 5987 3836
rect 5987 3780 5991 3836
rect 5927 3776 5991 3780
rect 6007 3836 6071 3840
rect 6007 3780 6011 3836
rect 6011 3780 6067 3836
rect 6067 3780 6071 3836
rect 6007 3776 6071 3780
rect 6087 3836 6151 3840
rect 6087 3780 6091 3836
rect 6091 3780 6147 3836
rect 6147 3780 6151 3836
rect 6087 3776 6151 3780
rect 9111 3836 9175 3840
rect 9111 3780 9115 3836
rect 9115 3780 9171 3836
rect 9171 3780 9175 3836
rect 9111 3776 9175 3780
rect 9191 3836 9255 3840
rect 9191 3780 9195 3836
rect 9195 3780 9251 3836
rect 9251 3780 9255 3836
rect 9191 3776 9255 3780
rect 9271 3836 9335 3840
rect 9271 3780 9275 3836
rect 9275 3780 9331 3836
rect 9331 3780 9335 3836
rect 9271 3776 9335 3780
rect 9351 3836 9415 3840
rect 9351 3780 9355 3836
rect 9355 3780 9411 3836
rect 9411 3780 9415 3836
rect 9351 3776 9415 3780
rect 4215 3292 4279 3296
rect 4215 3236 4219 3292
rect 4219 3236 4275 3292
rect 4275 3236 4279 3292
rect 4215 3232 4279 3236
rect 4295 3292 4359 3296
rect 4295 3236 4299 3292
rect 4299 3236 4355 3292
rect 4355 3236 4359 3292
rect 4295 3232 4359 3236
rect 4375 3292 4439 3296
rect 4375 3236 4379 3292
rect 4379 3236 4435 3292
rect 4435 3236 4439 3292
rect 4375 3232 4439 3236
rect 4455 3292 4519 3296
rect 4455 3236 4459 3292
rect 4459 3236 4515 3292
rect 4515 3236 4519 3292
rect 4455 3232 4519 3236
rect 7479 3292 7543 3296
rect 7479 3236 7483 3292
rect 7483 3236 7539 3292
rect 7539 3236 7543 3292
rect 7479 3232 7543 3236
rect 7559 3292 7623 3296
rect 7559 3236 7563 3292
rect 7563 3236 7619 3292
rect 7619 3236 7623 3292
rect 7559 3232 7623 3236
rect 7639 3292 7703 3296
rect 7639 3236 7643 3292
rect 7643 3236 7699 3292
rect 7699 3236 7703 3292
rect 7639 3232 7703 3236
rect 7719 3292 7783 3296
rect 7719 3236 7723 3292
rect 7723 3236 7779 3292
rect 7779 3236 7783 3292
rect 7719 3232 7783 3236
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5847 2748 5911 2752
rect 5847 2692 5851 2748
rect 5851 2692 5907 2748
rect 5907 2692 5911 2748
rect 5847 2688 5911 2692
rect 5927 2748 5991 2752
rect 5927 2692 5931 2748
rect 5931 2692 5987 2748
rect 5987 2692 5991 2748
rect 5927 2688 5991 2692
rect 6007 2748 6071 2752
rect 6007 2692 6011 2748
rect 6011 2692 6067 2748
rect 6067 2692 6071 2748
rect 6007 2688 6071 2692
rect 6087 2748 6151 2752
rect 6087 2692 6091 2748
rect 6091 2692 6147 2748
rect 6147 2692 6151 2748
rect 6087 2688 6151 2692
rect 9111 2748 9175 2752
rect 9111 2692 9115 2748
rect 9115 2692 9171 2748
rect 9171 2692 9175 2748
rect 9111 2688 9175 2692
rect 9191 2748 9255 2752
rect 9191 2692 9195 2748
rect 9195 2692 9251 2748
rect 9251 2692 9255 2748
rect 9191 2688 9255 2692
rect 9271 2748 9335 2752
rect 9271 2692 9275 2748
rect 9275 2692 9331 2748
rect 9331 2692 9335 2748
rect 9271 2688 9335 2692
rect 9351 2748 9415 2752
rect 9351 2692 9355 2748
rect 9355 2692 9411 2748
rect 9411 2692 9415 2748
rect 9351 2688 9415 2692
rect 4215 2204 4279 2208
rect 4215 2148 4219 2204
rect 4219 2148 4275 2204
rect 4275 2148 4279 2204
rect 4215 2144 4279 2148
rect 4295 2204 4359 2208
rect 4295 2148 4299 2204
rect 4299 2148 4355 2204
rect 4355 2148 4359 2204
rect 4295 2144 4359 2148
rect 4375 2204 4439 2208
rect 4375 2148 4379 2204
rect 4379 2148 4435 2204
rect 4435 2148 4439 2204
rect 4375 2144 4439 2148
rect 4455 2204 4519 2208
rect 4455 2148 4459 2204
rect 4459 2148 4515 2204
rect 4515 2148 4519 2204
rect 4455 2144 4519 2148
rect 7479 2204 7543 2208
rect 7479 2148 7483 2204
rect 7483 2148 7539 2204
rect 7539 2148 7543 2204
rect 7479 2144 7543 2148
rect 7559 2204 7623 2208
rect 7559 2148 7563 2204
rect 7563 2148 7619 2204
rect 7619 2148 7623 2204
rect 7559 2144 7623 2148
rect 7639 2204 7703 2208
rect 7639 2148 7643 2204
rect 7643 2148 7699 2204
rect 7699 2148 7703 2204
rect 7639 2144 7703 2148
rect 7719 2204 7783 2208
rect 7719 2148 7723 2204
rect 7723 2148 7779 2204
rect 7779 2148 7783 2204
rect 7719 2144 7783 2148
<< metal4 >>
rect 2575 77824 2896 77840
rect 2575 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2575 76736 2896 77760
rect 2575 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2575 75648 2896 76672
rect 2575 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2575 74560 2896 75584
rect 2575 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2575 73472 2896 74496
rect 2575 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2575 72384 2896 73408
rect 2575 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2575 71296 2896 72320
rect 2575 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2575 70208 2896 71232
rect 2575 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2575 69120 2896 70144
rect 2575 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2575 68032 2896 69056
rect 2575 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2575 66944 2896 67968
rect 2575 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2575 65856 2896 66880
rect 2575 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2575 64768 2896 65792
rect 2575 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2575 63680 2896 64704
rect 2575 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2575 62592 2896 63616
rect 4207 77280 4527 77840
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 76192 4527 77216
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 75104 4527 76128
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 74016 4527 75040
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 72928 4527 73952
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 71840 4527 72864
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 70752 4527 71776
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 69664 4527 70688
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 68576 4527 69600
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 67488 4527 68512
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 66400 4527 67424
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 65312 4527 66336
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 64224 4527 65248
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 63136 4527 64160
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 3555 62796 3621 62797
rect 3555 62732 3556 62796
rect 3620 62732 3621 62796
rect 3555 62731 3621 62732
rect 2575 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2575 61504 2896 62528
rect 2575 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2575 60416 2896 61440
rect 2575 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2575 59328 2896 60352
rect 3371 59532 3437 59533
rect 3371 59468 3372 59532
rect 3436 59468 3437 59532
rect 3371 59467 3437 59468
rect 2575 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2575 58240 2896 59264
rect 2575 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2575 57152 2896 58176
rect 2575 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2575 56064 2896 57088
rect 2575 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2575 54976 2896 56000
rect 2575 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2575 53888 2896 54912
rect 2575 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2575 52800 2896 53824
rect 2575 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2575 51712 2896 52736
rect 2575 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2575 50624 2896 51648
rect 3187 51236 3253 51237
rect 3187 51172 3188 51236
rect 3252 51172 3253 51236
rect 3187 51171 3253 51172
rect 3190 50965 3250 51171
rect 3187 50964 3253 50965
rect 3187 50900 3188 50964
rect 3252 50900 3253 50964
rect 3187 50899 3253 50900
rect 2575 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2575 49536 2896 50560
rect 2575 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2575 48448 2896 49472
rect 2575 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2575 47360 2896 48384
rect 2575 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2575 46272 2896 47296
rect 2575 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2575 45184 2896 46208
rect 2575 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2575 44096 2896 45120
rect 2575 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2575 43008 2896 44032
rect 2575 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2575 41920 2896 42944
rect 2575 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2575 40832 2896 41856
rect 2575 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2575 39744 2896 40768
rect 2575 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2575 38656 2896 39680
rect 2575 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2575 37568 2896 38592
rect 2575 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2575 36480 2896 37504
rect 3374 37229 3434 59467
rect 3558 44437 3618 62731
rect 4207 62048 4527 63072
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 60960 4527 61984
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 59872 4527 60896
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 58784 4527 59808
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 57696 4527 58720
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 4207 56608 4527 57632
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 55520 4527 56544
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 54432 4527 55456
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 53344 4527 54368
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 52256 4527 53280
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 51168 4527 52192
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 3739 50964 3805 50965
rect 3739 50900 3740 50964
rect 3804 50900 3805 50964
rect 3739 50899 3805 50900
rect 3742 45389 3802 50899
rect 4207 50080 4527 51104
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 48992 4527 50016
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 47904 4527 48928
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 46816 4527 47840
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 45728 4527 46752
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 3739 45388 3805 45389
rect 3739 45324 3740 45388
rect 3804 45324 3805 45388
rect 3739 45323 3805 45324
rect 4207 44640 4527 45664
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 3555 44436 3621 44437
rect 3555 44372 3556 44436
rect 3620 44372 3621 44436
rect 3555 44371 3621 44372
rect 4207 43552 4527 44576
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 42464 4527 43488
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 41376 4527 42400
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 40288 4527 41312
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 39200 4527 40224
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 38112 4527 39136
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 3371 37228 3437 37229
rect 3371 37164 3372 37228
rect 3436 37164 3437 37228
rect 3371 37163 3437 37164
rect 2575 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2575 35392 2896 36416
rect 2575 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2575 34304 2896 35328
rect 2575 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2575 33216 2896 34240
rect 2575 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2575 32128 2896 33152
rect 2575 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2575 31040 2896 32064
rect 2575 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2575 29952 2896 30976
rect 2575 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2575 28864 2896 29888
rect 2575 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2575 27776 2896 28800
rect 2575 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2575 26688 2896 27712
rect 2575 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2575 25600 2896 26624
rect 2575 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2575 24512 2896 25536
rect 2575 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2575 23424 2896 24448
rect 2575 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2575 22336 2896 23360
rect 2575 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2575 21248 2896 22272
rect 2575 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2575 20160 2896 21184
rect 2575 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2575 19072 2896 20096
rect 2575 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2575 17984 2896 19008
rect 2575 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2575 16896 2896 17920
rect 2575 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2575 15808 2896 16832
rect 2575 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2575 14720 2896 15744
rect 2575 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2575 13632 2896 14656
rect 2575 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2575 12544 2896 13568
rect 2575 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2575 11456 2896 12480
rect 2575 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2575 10368 2896 11392
rect 2575 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2575 9280 2896 10304
rect 2575 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2575 8192 2896 9216
rect 2575 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2575 7104 2896 8128
rect 2575 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2575 6016 2896 7040
rect 2575 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2575 4928 2896 5952
rect 2575 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2575 3840 2896 4864
rect 2575 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2575 2752 2896 3776
rect 2575 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2575 2128 2896 2688
rect 4207 37024 4527 38048
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 35936 4527 36960
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 34848 4527 35872
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 33760 4527 34784
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 32672 4527 33696
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 31584 4527 32608
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 30496 4527 31520
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 29408 4527 30432
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 28320 4527 29344
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 27232 4527 28256
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 26144 4527 27168
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 25056 4527 26080
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 23968 4527 24992
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 22880 4527 23904
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 21792 4527 22816
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 20704 4527 21728
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 19616 4527 20640
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 18528 4527 19552
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 17440 4527 18464
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 16352 4527 17376
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 15264 4527 16288
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 14176 4527 15200
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 13088 4527 14112
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 12000 4527 13024
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 10912 4527 11936
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 9824 4527 10848
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 8736 4527 9760
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 7648 4527 8672
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 6560 4527 7584
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 5472 4527 6496
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 4384 4527 5408
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 3296 4527 4320
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 2208 4527 3232
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2128 4527 2144
rect 5839 77824 6159 77840
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 76736 6159 77760
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 75648 6159 76672
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 74560 6159 75584
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 73472 6159 74496
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 72384 6159 73408
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 71296 6159 72320
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 70208 6159 71232
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 69120 6159 70144
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 68032 6159 69056
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 66944 6159 67968
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 65856 6159 66880
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 64768 6159 65792
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 63680 6159 64704
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 62592 6159 63616
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 61504 6159 62528
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 60416 6159 61440
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 59328 6159 60352
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 58240 6159 59264
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 57152 6159 58176
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 56064 6159 57088
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 54976 6159 56000
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 53888 6159 54912
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 52800 6159 53824
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 51712 6159 52736
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 50624 6159 51648
rect 7471 77280 7791 77840
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 76192 7791 77216
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 75104 7791 76128
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 74016 7791 75040
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 72928 7791 73952
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 71840 7791 72864
rect 9103 77824 9423 77840
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 76736 9423 77760
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 75648 9423 76672
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 9103 74560 9423 75584
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 73472 9423 74496
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 72384 9423 73408
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 8523 71908 8589 71909
rect 8523 71844 8524 71908
rect 8588 71844 8589 71908
rect 8523 71843 8589 71844
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 70752 7791 71776
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 69664 7791 70688
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 68576 7791 69600
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 67488 7791 68512
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 66400 7791 67424
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 65312 7791 66336
rect 8339 66332 8405 66333
rect 8339 66268 8340 66332
rect 8404 66268 8405 66332
rect 8339 66267 8405 66268
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 64224 7791 65248
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 63136 7791 64160
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 62048 7791 63072
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 60960 7791 61984
rect 8155 61300 8221 61301
rect 8155 61236 8156 61300
rect 8220 61236 8221 61300
rect 8155 61235 8221 61236
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 59872 7791 60896
rect 8158 60621 8218 61235
rect 8155 60620 8221 60621
rect 8155 60556 8156 60620
rect 8220 60556 8221 60620
rect 8155 60555 8221 60556
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 58784 7791 59808
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 57696 7791 58720
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 56608 7791 57632
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 55520 7791 56544
rect 7971 55860 8037 55861
rect 7971 55796 7972 55860
rect 8036 55796 8037 55860
rect 7971 55795 8037 55796
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 54432 7791 55456
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 53344 7791 54368
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 52256 7791 53280
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7051 51508 7117 51509
rect 7051 51444 7052 51508
rect 7116 51444 7117 51508
rect 7051 51443 7117 51444
rect 6683 51236 6749 51237
rect 6683 51172 6684 51236
rect 6748 51172 6749 51236
rect 6683 51171 6749 51172
rect 6686 50965 6746 51171
rect 6683 50964 6749 50965
rect 6683 50900 6684 50964
rect 6748 50900 6749 50964
rect 6683 50899 6749 50900
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 49536 6159 50560
rect 7054 49605 7114 51443
rect 7471 51168 7791 52192
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 50080 7791 51104
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7051 49604 7117 49605
rect 7051 49540 7052 49604
rect 7116 49540 7117 49604
rect 7051 49539 7117 49540
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5839 48448 6159 49472
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5839 47360 6159 48384
rect 7471 48992 7791 50016
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7235 48108 7301 48109
rect 7235 48044 7236 48108
rect 7300 48044 7301 48108
rect 7235 48043 7301 48044
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 46272 6159 47296
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 45184 6159 46208
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 44096 6159 45120
rect 7238 44301 7298 48043
rect 7471 47904 7791 48928
rect 7974 48517 8034 55795
rect 8155 53548 8221 53549
rect 8155 53484 8156 53548
rect 8220 53484 8221 53548
rect 8155 53483 8221 53484
rect 8158 51237 8218 53483
rect 8155 51236 8221 51237
rect 8155 51172 8156 51236
rect 8220 51172 8221 51236
rect 8155 51171 8221 51172
rect 8155 50420 8221 50421
rect 8155 50356 8156 50420
rect 8220 50356 8221 50420
rect 8155 50355 8221 50356
rect 8158 48789 8218 50355
rect 8155 48788 8221 48789
rect 8155 48724 8156 48788
rect 8220 48724 8221 48788
rect 8155 48723 8221 48724
rect 7971 48516 8037 48517
rect 7971 48452 7972 48516
rect 8036 48452 8037 48516
rect 7971 48451 8037 48452
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 7471 46816 7791 47840
rect 8155 47700 8221 47701
rect 8155 47636 8156 47700
rect 8220 47636 8221 47700
rect 8155 47635 8221 47636
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 45728 7791 46752
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 44640 7791 45664
rect 7971 44844 8037 44845
rect 7971 44780 7972 44844
rect 8036 44780 8037 44844
rect 7971 44779 8037 44780
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7235 44300 7301 44301
rect 7235 44236 7236 44300
rect 7300 44236 7301 44300
rect 7235 44235 7301 44236
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 43008 6159 44032
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 41920 6159 42944
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5839 40832 6159 41856
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 39744 6159 40768
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 38656 6159 39680
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 37568 6159 38592
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 36480 6159 37504
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 35392 6159 36416
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 34304 6159 35328
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 33216 6159 34240
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 32128 6159 33152
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 31040 6159 32064
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 29952 6159 30976
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 28864 6159 29888
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 27776 6159 28800
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 26688 6159 27712
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 25600 6159 26624
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 24512 6159 25536
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 23424 6159 24448
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 22336 6159 23360
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 21248 6159 22272
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 20160 6159 21184
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 19072 6159 20096
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 17984 6159 19008
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 16896 6159 17920
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 15808 6159 16832
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 14720 6159 15744
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 13632 6159 14656
rect 7471 43552 7791 44576
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 42464 7791 43488
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 41376 7791 42400
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 7471 40288 7791 41312
rect 7974 40493 8034 44779
rect 8158 43077 8218 47635
rect 8155 43076 8221 43077
rect 8155 43012 8156 43076
rect 8220 43012 8221 43076
rect 8155 43011 8221 43012
rect 8342 42805 8402 66267
rect 8339 42804 8405 42805
rect 8339 42740 8340 42804
rect 8404 42740 8405 42804
rect 8339 42739 8405 42740
rect 8155 41580 8221 41581
rect 8155 41516 8156 41580
rect 8220 41516 8221 41580
rect 8155 41515 8221 41516
rect 8158 41309 8218 41515
rect 8155 41308 8221 41309
rect 8155 41244 8156 41308
rect 8220 41244 8221 41308
rect 8155 41243 8221 41244
rect 8526 40765 8586 71843
rect 9103 71296 9423 72320
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 70208 9423 71232
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 8891 69324 8957 69325
rect 8891 69260 8892 69324
rect 8956 69260 8957 69324
rect 8891 69259 8957 69260
rect 8707 67692 8773 67693
rect 8707 67628 8708 67692
rect 8772 67628 8773 67692
rect 8707 67627 8773 67628
rect 8523 40764 8589 40765
rect 8523 40700 8524 40764
rect 8588 40700 8589 40764
rect 8523 40699 8589 40700
rect 7971 40492 8037 40493
rect 7971 40428 7972 40492
rect 8036 40428 8037 40492
rect 7971 40427 8037 40428
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 7471 39200 7791 40224
rect 8523 39540 8589 39541
rect 8523 39476 8524 39540
rect 8588 39476 8589 39540
rect 8523 39475 8589 39476
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 38112 7791 39136
rect 8526 38317 8586 39475
rect 8339 38316 8405 38317
rect 8339 38252 8340 38316
rect 8404 38252 8405 38316
rect 8339 38251 8405 38252
rect 8523 38316 8589 38317
rect 8523 38252 8524 38316
rect 8588 38252 8589 38316
rect 8523 38251 8589 38252
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 37024 7791 38048
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 35936 7791 36960
rect 8342 36277 8402 38251
rect 8523 37908 8589 37909
rect 8523 37844 8524 37908
rect 8588 37844 8589 37908
rect 8523 37843 8589 37844
rect 8339 36276 8405 36277
rect 8339 36212 8340 36276
rect 8404 36212 8405 36276
rect 8339 36211 8405 36212
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 34848 7791 35872
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 33760 7791 34784
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 32672 7791 33696
rect 8526 33557 8586 37843
rect 8710 34509 8770 67627
rect 8894 38861 8954 69259
rect 9103 69120 9423 70144
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 68032 9423 69056
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 66944 9423 67968
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 65856 9423 66880
rect 9627 66604 9693 66605
rect 9627 66540 9628 66604
rect 9692 66540 9693 66604
rect 9627 66539 9693 66540
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 64768 9423 65792
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 63680 9423 64704
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 62592 9423 63616
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 61504 9423 62528
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 60416 9423 61440
rect 9630 61301 9690 66539
rect 9627 61300 9693 61301
rect 9627 61236 9628 61300
rect 9692 61236 9693 61300
rect 9627 61235 9693 61236
rect 9627 60620 9693 60621
rect 9627 60556 9628 60620
rect 9692 60556 9693 60620
rect 9627 60555 9693 60556
rect 10179 60620 10245 60621
rect 10179 60556 10180 60620
rect 10244 60556 10245 60620
rect 10179 60555 10245 60556
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 59328 9423 60352
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 58240 9423 59264
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 57152 9423 58176
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 56064 9423 57088
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 54976 9423 56000
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 53888 9423 54912
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 52800 9423 53824
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 51712 9423 52736
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 50624 9423 51648
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 49536 9423 50560
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 48448 9423 49472
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 47360 9423 48384
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 46272 9423 47296
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 45184 9423 46208
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 44096 9423 45120
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 43008 9423 44032
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 41920 9423 42944
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 40832 9423 41856
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 39744 9423 40768
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 8891 38860 8957 38861
rect 8891 38796 8892 38860
rect 8956 38796 8957 38860
rect 8891 38795 8957 38796
rect 9103 38656 9423 39680
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 8891 38180 8957 38181
rect 8891 38116 8892 38180
rect 8956 38116 8957 38180
rect 8891 38115 8957 38116
rect 8894 36005 8954 38115
rect 9103 37568 9423 38592
rect 9630 37773 9690 60555
rect 9995 46340 10061 46341
rect 9995 46276 9996 46340
rect 10060 46276 10061 46340
rect 9995 46275 10061 46276
rect 9811 38588 9877 38589
rect 9811 38524 9812 38588
rect 9876 38524 9877 38588
rect 9811 38523 9877 38524
rect 9627 37772 9693 37773
rect 9627 37708 9628 37772
rect 9692 37708 9693 37772
rect 9627 37707 9693 37708
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 36480 9423 37504
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 8891 36004 8957 36005
rect 8891 35940 8892 36004
rect 8956 35940 8957 36004
rect 8891 35939 8957 35940
rect 9103 35392 9423 36416
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 8707 34508 8773 34509
rect 8707 34444 8708 34508
rect 8772 34444 8773 34508
rect 8707 34443 8773 34444
rect 9103 34304 9423 35328
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 8523 33556 8589 33557
rect 8523 33492 8524 33556
rect 8588 33492 8589 33556
rect 8523 33491 8589 33492
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 31584 7791 32608
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 30496 7791 31520
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 29408 7791 30432
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 7471 28320 7791 29344
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 27232 7791 28256
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 26144 7791 27168
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 25056 7791 26080
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 23968 7791 24992
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 22880 7791 23904
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 21792 7791 22816
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 20704 7791 21728
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 19616 7791 20640
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 18528 7791 19552
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 17440 7791 18464
rect 9103 33216 9423 34240
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 32128 9423 33152
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 31040 9423 32064
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 29952 9423 30976
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 28864 9423 29888
rect 9814 29749 9874 38523
rect 9998 30837 10058 46275
rect 10182 40493 10242 60555
rect 10731 56268 10797 56269
rect 10731 56204 10732 56268
rect 10796 56204 10797 56268
rect 10731 56203 10797 56204
rect 10363 53276 10429 53277
rect 10363 53212 10364 53276
rect 10428 53212 10429 53276
rect 10363 53211 10429 53212
rect 10366 42397 10426 53211
rect 10734 50149 10794 56203
rect 11467 54364 11533 54365
rect 11467 54300 11468 54364
rect 11532 54300 11533 54364
rect 11467 54299 11533 54300
rect 10915 52460 10981 52461
rect 10915 52396 10916 52460
rect 10980 52396 10981 52460
rect 10915 52395 10981 52396
rect 10731 50148 10797 50149
rect 10731 50084 10732 50148
rect 10796 50084 10797 50148
rect 10731 50083 10797 50084
rect 10731 42668 10797 42669
rect 10731 42604 10732 42668
rect 10796 42604 10797 42668
rect 10731 42603 10797 42604
rect 10547 42532 10613 42533
rect 10547 42468 10548 42532
rect 10612 42468 10613 42532
rect 10547 42467 10613 42468
rect 10363 42396 10429 42397
rect 10363 42332 10364 42396
rect 10428 42332 10429 42396
rect 10363 42331 10429 42332
rect 10179 40492 10245 40493
rect 10179 40428 10180 40492
rect 10244 40428 10245 40492
rect 10179 40427 10245 40428
rect 10550 40221 10610 42467
rect 10547 40220 10613 40221
rect 10547 40156 10548 40220
rect 10612 40156 10613 40220
rect 10547 40155 10613 40156
rect 10363 39676 10429 39677
rect 10363 39612 10364 39676
rect 10428 39612 10429 39676
rect 10363 39611 10429 39612
rect 10179 36684 10245 36685
rect 10179 36620 10180 36684
rect 10244 36620 10245 36684
rect 10179 36619 10245 36620
rect 9995 30836 10061 30837
rect 9995 30772 9996 30836
rect 10060 30772 10061 30836
rect 9995 30771 10061 30772
rect 9811 29748 9877 29749
rect 9811 29684 9812 29748
rect 9876 29684 9877 29748
rect 9811 29683 9877 29684
rect 10182 29613 10242 36619
rect 10179 29612 10245 29613
rect 10179 29548 10180 29612
rect 10244 29548 10245 29612
rect 10179 29547 10245 29548
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 27776 9423 28800
rect 10366 28253 10426 39611
rect 10547 36820 10613 36821
rect 10547 36756 10548 36820
rect 10612 36756 10613 36820
rect 10547 36755 10613 36756
rect 10550 33421 10610 36755
rect 10547 33420 10613 33421
rect 10547 33356 10548 33420
rect 10612 33356 10613 33420
rect 10547 33355 10613 33356
rect 10547 33148 10613 33149
rect 10547 33084 10548 33148
rect 10612 33084 10613 33148
rect 10547 33083 10613 33084
rect 10550 31789 10610 33083
rect 10734 32605 10794 42603
rect 10918 42125 10978 52395
rect 11470 50557 11530 54299
rect 11467 50556 11533 50557
rect 11467 50492 11468 50556
rect 11532 50492 11533 50556
rect 11467 50491 11533 50492
rect 11099 44436 11165 44437
rect 11099 44372 11100 44436
rect 11164 44372 11165 44436
rect 11099 44371 11165 44372
rect 10915 42124 10981 42125
rect 10915 42060 10916 42124
rect 10980 42060 10981 42124
rect 10915 42059 10981 42060
rect 10915 39676 10981 39677
rect 10915 39612 10916 39676
rect 10980 39612 10981 39676
rect 10915 39611 10981 39612
rect 10731 32604 10797 32605
rect 10731 32540 10732 32604
rect 10796 32540 10797 32604
rect 10731 32539 10797 32540
rect 10731 32060 10797 32061
rect 10731 31996 10732 32060
rect 10796 31996 10797 32060
rect 10731 31995 10797 31996
rect 10547 31788 10613 31789
rect 10547 31724 10548 31788
rect 10612 31724 10613 31788
rect 10547 31723 10613 31724
rect 10734 30565 10794 31995
rect 10731 30564 10797 30565
rect 10731 30500 10732 30564
rect 10796 30500 10797 30564
rect 10731 30499 10797 30500
rect 10918 29341 10978 39611
rect 10915 29340 10981 29341
rect 10915 29276 10916 29340
rect 10980 29276 10981 29340
rect 10915 29275 10981 29276
rect 11102 28930 11162 44371
rect 11467 43484 11533 43485
rect 11467 43420 11468 43484
rect 11532 43420 11533 43484
rect 11467 43419 11533 43420
rect 11470 38725 11530 43419
rect 11467 38724 11533 38725
rect 11467 38660 11468 38724
rect 11532 38660 11533 38724
rect 11467 38659 11533 38660
rect 11651 36820 11717 36821
rect 11651 36756 11652 36820
rect 11716 36756 11717 36820
rect 11651 36755 11717 36756
rect 11654 29749 11714 36755
rect 11651 29748 11717 29749
rect 11651 29684 11652 29748
rect 11716 29684 11717 29748
rect 11651 29683 11717 29684
rect 10918 28870 11162 28930
rect 10363 28252 10429 28253
rect 10363 28188 10364 28252
rect 10428 28188 10429 28252
rect 10363 28187 10429 28188
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 26688 9423 27712
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 25600 9423 26624
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 24512 9423 25536
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 23424 9423 24448
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 22336 9423 23360
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 21248 9423 22272
rect 10918 22269 10978 28870
rect 10915 22268 10981 22269
rect 10915 22204 10916 22268
rect 10980 22204 10981 22268
rect 10915 22203 10981 22204
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 20160 9423 21184
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 19072 9423 20096
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 8891 18460 8957 18461
rect 8891 18396 8892 18460
rect 8956 18396 8957 18460
rect 8891 18395 8957 18396
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 16352 7791 17376
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 15264 7791 16288
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7235 14652 7301 14653
rect 7235 14588 7236 14652
rect 7300 14588 7301 14652
rect 7235 14587 7301 14588
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 12544 6159 13568
rect 7238 13565 7298 14587
rect 7471 14176 7791 15200
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7235 13564 7301 13565
rect 7235 13500 7236 13564
rect 7300 13500 7301 13564
rect 7235 13499 7301 13500
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 11456 6159 12480
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 10368 6159 11392
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 9280 6159 10304
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 8192 6159 9216
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 7104 6159 8128
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 6016 6159 7040
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 4928 6159 5952
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 3840 6159 4864
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 2752 6159 3776
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2128 6159 2688
rect 7471 13088 7791 14112
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 12000 7791 13024
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 10912 7791 11936
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 9824 7791 10848
rect 8894 10165 8954 18395
rect 9103 17984 9423 19008
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 16896 9423 17920
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 15808 9423 16832
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 14720 9423 15744
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 13632 9423 14656
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 12544 9423 13568
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 11456 9423 12480
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 10368 9423 11392
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 8891 10164 8957 10165
rect 8891 10100 8892 10164
rect 8956 10100 8957 10164
rect 8891 10099 8957 10100
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 8736 7791 9760
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 7648 7791 8672
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 6560 7791 7584
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 5472 7791 6496
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 4384 7791 5408
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 3296 7791 4320
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 7471 2208 7791 3232
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2128 7791 2144
rect 9103 9280 9423 10304
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 8192 9423 9216
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 7104 9423 8128
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 6016 9423 7040
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 4928 9423 5952
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 3840 9423 4864
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 2752 9423 3776
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2128 9423 2688
use sky130_fd_sc_hd__buf_2  output214 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1635444444
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1635444444
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output178 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1635444444
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1635444444
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1635444444
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 1635444444
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1635444444
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1635444444
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 1635444444
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1635444444
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1635444444
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1635444444
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input112 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 7544 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8372 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1635444444
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1635444444
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1635444444
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1635444444
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1635444444
transform 1 0 9292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_7
timestamp 1635444444
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1635444444
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1635444444
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1635444444
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1635444444
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1635444444
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1635444444
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1635444444
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1635444444
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1635444444
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1635444444
transform 1 0 9292 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_3_19
timestamp 1635444444
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_7
timestamp 1635444444
transform 1 0 1748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1635444444
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_31
timestamp 1635444444
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1635444444
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1635444444
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1635444444
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_81
timestamp 1635444444
transform 1 0 8556 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1635444444
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1635444444
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1635444444
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input113
timestamp 1635444444
transform 1 0 9292 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1635444444
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_7
timestamp 1635444444
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1635444444
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1635444444
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1635444444
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1635444444
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1635444444
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1635444444
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1635444444
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9200 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1635444444
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9384 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1635444444
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_7
timestamp 1635444444
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1635444444
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_31
timestamp 1635444444
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1635444444
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635444444
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_69
timestamp 1635444444
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp 1635444444
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1635444444
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1635444444
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1635444444
transform 1 0 8096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1635444444
transform 1 0 9200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1635444444
transform 1 0 9016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1635444444
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _115_
timestamp 1635444444
transform 1 0 9384 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1635444444
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1635444444
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_19
timestamp 1635444444
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_7
timestamp 1635444444
transform 1 0 1748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1635444444
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1635444444
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1635444444
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1635444444
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1635444444
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_31
timestamp 1635444444
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1635444444
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1635444444
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1635444444
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1635444444
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1635444444
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_73
timestamp 1635444444
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1635444444
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1635444444
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1635444444
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_2  _037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _038_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _114_
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_90
timestamp 1635444444
transform 1 0 9384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1635444444
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1635444444
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1635444444
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1635444444
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_94
timestamp 1635444444
transform 1 0 9752 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_102
timestamp 1635444444
transform 1 0 10488 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1635444444
transform 1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1635444444
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1635444444
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635444444
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1635444444
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1635444444
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1635444444
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1635444444
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1635444444
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1635444444
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1635444444
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1635444444
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _116_
timestamp 1635444444
transform 1 0 9384 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1635444444
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_7
timestamp 1635444444
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1635444444
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1635444444
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1635444444
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1635444444
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1635444444
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1635444444
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1635444444
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_89
timestamp 1635444444
transform 1 0 9292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1635444444
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp 1635444444
transform 1 0 9384 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1635444444
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1635444444
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1635444444
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1635444444
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1635444444
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1635444444
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1635444444
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1635444444
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1635444444
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1635444444
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1635444444
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_99
timestamp 1635444444
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input67 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_19
timestamp 1635444444
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_7
timestamp 1635444444
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1635444444
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1635444444
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1635444444
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1635444444
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1635444444
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1635444444
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp 1635444444
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_90
timestamp 1635444444
transform 1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_b_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input68
timestamp 1635444444
transform 1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1635444444
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1635444444
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1635444444
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1635444444
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1635444444
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1635444444
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1635444444
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1635444444
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1635444444
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1635444444
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1635444444
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_91
timestamp 1635444444
transform 1 0 9476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1635444444
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1635444444
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1635444444
transform 1 0 9108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1635444444
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1635444444
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1635444444
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_7
timestamp 1635444444
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1635444444
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1635444444
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1635444444
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1635444444
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1635444444
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1635444444
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1635444444
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1635444444
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1635444444
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_77
timestamp 1635444444
transform 1 0 8188 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_68
timestamp 1635444444
transform 1 0 7360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_76
timestamp 1635444444
transform 1 0 8096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1635444444
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_a_clk_i
timestamp 1635444444
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1635444444
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1635444444
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net199_2
timestamp 1635444444
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input74
timestamp 1635444444
transform 1 0 9660 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _127_
timestamp 1635444444
transform 1 0 9384 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1635444444
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_85
timestamp 1635444444
transform 1 0 8924 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_99
timestamp 1635444444
transform 1 0 10212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1635444444
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_19
timestamp 1635444444
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_7
timestamp 1635444444
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1635444444
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_31
timestamp 1635444444
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1635444444
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1635444444
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1635444444
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_66
timestamp 1635444444
transform 1 0 7176 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_72
timestamp 1635444444
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_76
timestamp 1635444444
transform 1 0 8096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _045_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _113_
timestamp 1635444444
transform 1 0 8464 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1635444444
transform 1 0 7820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1635444444
transform 1 0 10488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_89
timestamp 1635444444
transform 1 0 9292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _128_
timestamp 1635444444
transform 1 0 9384 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1635444444
transform 1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1635444444
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1635444444
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1635444444
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1635444444
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1635444444
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1635444444
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1635444444
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_57
timestamp 1635444444
transform 1 0 6348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_61
timestamp 1635444444
transform 1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1635444444
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_68
timestamp 1635444444
transform 1 0 7360 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1635444444
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1635444444
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _025_
timestamp 1635444444
transform 1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1635444444
transform 1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1635444444
transform 1 0 9200 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1635444444
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_101
timestamp 1635444444
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_90
timestamp 1635444444
transform 1 0 9384 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_98
timestamp 1635444444
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_19
timestamp 1635444444
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_7
timestamp 1635444444
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1635444444
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_31
timestamp 1635444444
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_43
timestamp 1635444444
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1635444444
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6532 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_75
timestamp 1635444444
transform 1 0 8004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_a_clk_i
timestamp 1635444444
transform 1 0 8372 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1635444444
transform 1 0 10212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1635444444
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_7
timestamp 1635444444
transform 1 0 1748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1635444444
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635444444
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1635444444
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 1635444444
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 1635444444
transform 1 0 5612 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1635444444
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_60
timestamp 1635444444
transform 1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _026_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1635444444
transform 1 0 5704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1635444444
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _178_
timestamp 1635444444
transform 1 0 6992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1635444444
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1635444444
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1635444444
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 1635444444
transform 1 0 9384 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1635444444
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1635444444
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 1635444444
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1635444444
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1635444444
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1635444444
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp 1635444444
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1635444444
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1635444444
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _046_
timestamp 1635444444
transform 1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _041_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 5336 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_45
timestamp 1635444444
transform 1 0 5244 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp 1635444444
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _172_
timestamp 1635444444
transform 1 0 6440 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _031__1
timestamp 1635444444
transform 1 0 6532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_54
timestamp 1635444444
transform 1 0 6072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1635444444
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1635444444
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 1635444444
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_67
timestamp 1635444444
transform 1 0 7268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1635444444
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _159_
timestamp 1635444444
transform 1 0 7176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _168_
timestamp 1635444444
transform 1 0 7636 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_b_clk_i
timestamp 1635444444
transform 1 0 8372 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1635444444
transform 1 0 9200 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1635444444
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1635444444
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _130_
timestamp 1635444444
transform 1 0 9384 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1635444444
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_7
timestamp 1635444444
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1635444444
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1635444444
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_43
timestamp 1635444444
transform 1 0 5060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1635444444
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_60
timestamp 1635444444
transform 1 0 6624 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1635444444
transform 1 0 5612 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1635444444
transform 1 0 7820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _170_
timestamp 1635444444
transform 1 0 8188 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _173_
timestamp 1635444444
transform 1 0 6992 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1635444444
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1635444444
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _131_
timestamp 1635444444
transform 1 0 9384 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1635444444
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_7
timestamp 1635444444
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1635444444
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1635444444
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1635444444
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_41
timestamp 1635444444
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_48
timestamp 1635444444
transform 1 0 5520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_55
timestamp 1635444444
transform 1 0 6164 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_b_clk_i
timestamp 1635444444
transform 1 0 6532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1635444444
transform 1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1635444444
transform 1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_63
timestamp 1635444444
transform 1 0 6900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1635444444
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1635444444
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__and4b_1  _032_
timestamp 1635444444
transform 1 0 7268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1635444444
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1635444444
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1635444444
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_19
timestamp 1635444444
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_7
timestamp 1635444444
transform 1 0 1748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1635444444
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1635444444
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_43
timestamp 1635444444
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1635444444
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1635444444
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1635444444
transform 1 0 6808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_65
timestamp 1635444444
transform 1 0 7084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_73
timestamp 1635444444
transform 1 0 7820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 1635444444
transform 1 0 8188 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_a_clk_i
timestamp 1635444444
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1635444444
transform 1 0 9200 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_86
timestamp 1635444444
transform 1 0 9016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1635444444
transform 1 0 10212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _133_
timestamp 1635444444
transform 1 0 9384 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1635444444
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_7
timestamp 1635444444
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1635444444
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1635444444
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1635444444
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_53
timestamp 1635444444
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_62
timestamp 1635444444
transform 1 0 6808 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1635444444
transform 1 0 6532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1635444444
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1635444444
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _039_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 7820 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1635444444
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1635444444
transform 1 0 9200 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1635444444
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1635444444
transform 1 0 9384 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1635444444
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1635444444
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1635444444
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1635444444
transform 1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1635444444
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1635444444
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1635444444
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1635444444
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _177_
timestamp 1635444444
transform 1 0 7544 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform 1 0 6900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1635444444
transform 1 0 9016 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1635444444
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 1635444444
transform 1 0 9384 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1635444444
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_7
timestamp 1635444444
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_19
timestamp 1635444444
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_7
timestamp 1635444444
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1635444444
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1635444444
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1635444444
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1635444444
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_31
timestamp 1635444444
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _036_
timestamp 1635444444
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp 1635444444
transform 1 0 6440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_61
timestamp 1635444444
transform 1 0 6716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1635444444
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_61
timestamp 1635444444
transform 1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_57
timestamp 1635444444
transform 1 0 6348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1635444444
transform 1 0 5980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_43
timestamp 1635444444
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1635444444
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1635444444
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_68
timestamp 1635444444
transform 1 0 7360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _027__3
timestamp 1635444444
transform 1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _029_
timestamp 1635444444
transform 1 0 7728 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _035_
timestamp 1635444444
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _175_
timestamp 1635444444
transform 1 0 7728 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _171_
timestamp 1635444444
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _135_
timestamp 1635444444
transform 1 0 9384 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_88
timestamp 1635444444
transform 1 0 9200 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1635444444
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _028_
timestamp 1635444444
transform 1 0 10212 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_102
timestamp 1635444444
transform 1 0 10488 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_96
timestamp 1635444444
transform 1 0 9936 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_102
timestamp 1635444444
transform 1 0 10488 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1635444444
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_7
timestamp 1635444444
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1635444444
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1635444444
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1635444444
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_53
timestamp 1635444444
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_62
timestamp 1635444444
transform 1 0 6808 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _027__4
timestamp 1635444444
transform 1 0 6532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_70
timestamp 1635444444
transform 1 0 7544 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1635444444
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _043_
timestamp 1635444444
transform 1 0 7728 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1635444444
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_99
timestamp 1635444444
transform 1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _047_
timestamp 1635444444
transform 1 0 9384 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_19
timestamp 1635444444
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_7
timestamp 1635444444
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1635444444
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1635444444
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1635444444
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1635444444
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_68
timestamp 1635444444
transform 1 0 7360 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_76
timestamp 1635444444
transform 1 0 8096 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_80
timestamp 1635444444
transform 1 0 8464 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1635444444
transform 1 0 8188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1635444444
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1635444444
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1635444444
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1635444444
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_90
timestamp 1635444444
transform 1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_98
timestamp 1635444444
transform 1 0 10120 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1635444444
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1635444444
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1635444444
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1635444444
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1635444444
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_65
timestamp 1635444444
transform 1 0 7084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_69
timestamp 1635444444
transform 1 0 7452 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1635444444
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1635444444
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1635444444
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1635444444
transform 1 0 7544 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1635444444
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_102
timestamp 1635444444
transform 1 0 10488 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _139_
timestamp 1635444444
transform 1 0 9384 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1635444444
transform 1 0 10212 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_19
timestamp 1635444444
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_7
timestamp 1635444444
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1635444444
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1635444444
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1635444444
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1635444444
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1635444444
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_75
timestamp 1635444444
transform 1 0 8004 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1635444444
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1635444444
transform 1 0 8740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1635444444
transform 1 0 8096 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_86
timestamp 1635444444
transform 1 0 9016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1635444444
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1635444444
transform 1 0 9108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9384 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp 1635444444
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_7
timestamp 1635444444
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1635444444
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1635444444
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1635444444
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1635444444
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1635444444
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1635444444
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1635444444
transform 1 0 8188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1635444444
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1635444444
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _136_
timestamp 1635444444
transform 1 0 9384 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_19
timestamp 1635444444
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_7
timestamp 1635444444
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1635444444
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_7
timestamp 1635444444
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1635444444
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1635444444
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_31
timestamp 1635444444
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1635444444
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1635444444
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_43
timestamp 1635444444
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1635444444
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1635444444
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_69
timestamp 1635444444
transform 1 0 7452 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_75
timestamp 1635444444
transform 1 0 8004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1635444444
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1635444444
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1635444444
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1635444444
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1635444444
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1635444444
transform 1 0 8096 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1635444444
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_90
timestamp 1635444444
transform 1 0 9384 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_86
timestamp 1635444444
transform 1 0 9016 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1635444444
transform 1 0 9200 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1635444444
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_98
timestamp 1635444444
transform 1 0 10120 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1635444444
transform 1 0 10396 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1635444444
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1635444444
transform 1 0 9292 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_35_19
timestamp 1635444444
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_7
timestamp 1635444444
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1635444444
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_31
timestamp 1635444444
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_43
timestamp 1635444444
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1635444444
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1635444444
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_69
timestamp 1635444444
transform 1 0 7452 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_75
timestamp 1635444444
transform 1 0 8004 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _140_
timestamp 1635444444
transform 1 0 8096 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp 1635444444
transform 1 0 8924 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1635444444
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input91
timestamp 1635444444
transform 1 0 9292 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1635444444
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1635444444
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1635444444
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1635444444
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1635444444
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1635444444
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_65
timestamp 1635444444
transform 1 0 7084 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_73
timestamp 1635444444
transform 1 0 7820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1635444444
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1635444444
transform 1 0 8096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1635444444
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input92
timestamp 1635444444
transform 1 0 9292 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_37_19
timestamp 1635444444
transform 1 0 2852 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_7
timestamp 1635444444
transform 1 0 1748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1635444444
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_31
timestamp 1635444444
transform 1 0 3956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_43
timestamp 1635444444
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1635444444
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1635444444
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp 1635444444
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _141_
timestamp 1635444444
transform 1 0 8188 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1635444444
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1635444444
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _137_
timestamp 1635444444
transform 1 0 9384 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_38_19
timestamp 1635444444
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_7
timestamp 1635444444
transform 1 0 1748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1635444444
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1635444444
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1635444444
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1635444444
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1635444444
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1635444444
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1635444444
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1635444444
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1635444444
transform 1 0 9292 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1635444444
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _138_
timestamp 1635444444
transform 1 0 9384 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_39_19
timestamp 1635444444
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_7
timestamp 1635444444
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1635444444
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1635444444
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1635444444
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1635444444
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_31
timestamp 1635444444
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1635444444
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1635444444
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1635444444
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1635444444
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1635444444
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1635444444
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1635444444
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_81
timestamp 1635444444
transform 1 0 8556 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1635444444
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1635444444
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1635444444
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1635444444
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input97
timestamp 1635444444
transform 1 0 9108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _142_
timestamp 1635444444
transform 1 0 9384 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_91
timestamp 1635444444
transform 1 0 9476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1635444444
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_86
timestamp 1635444444
transform 1 0 9016 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1635444444
transform 1 0 9200 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1635444444
transform 1 0 9844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1635444444
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1635444444
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_19
timestamp 1635444444
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_7
timestamp 1635444444
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1635444444
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_31
timestamp 1635444444
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_43
timestamp 1635444444
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1635444444
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1635444444
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_81
timestamp 1635444444
transform 1 0 8556 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_91
timestamp 1635444444
transform 1 0 9476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1635444444
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1635444444
transform 1 0 9844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1635444444
transform 1 0 9108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1635444444
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1635444444
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1635444444
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1635444444
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1635444444
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1635444444
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1635444444
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1635444444
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_89
timestamp 1635444444
transform 1 0 9292 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1635444444
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 10856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _143_
timestamp 1635444444
transform 1 0 9384 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_43_19
timestamp 1635444444
transform 1 0 2852 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_7
timestamp 1635444444
transform 1 0 1748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1635444444
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_31
timestamp 1635444444
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_43
timestamp 1635444444
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1635444444
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1635444444
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1635444444
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_81
timestamp 1635444444
transform 1 0 8556 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_91
timestamp 1635444444
transform 1 0 9476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1635444444
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1635444444
transform 1 0 9844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1635444444
transform 1 0 9108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1635444444
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_7
timestamp 1635444444
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1635444444
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1635444444
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1635444444
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1635444444
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1635444444
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1635444444
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1635444444
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1635444444
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_93
timestamp 1635444444
transform 1 0 9660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_99
timestamp 1635444444
transform 1 0 10212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1635444444
transform 1 0 9844 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_19
timestamp 1635444444
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1635444444
transform 1 0 1748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1635444444
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_31
timestamp 1635444444
transform 1 0 3956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_43
timestamp 1635444444
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1635444444
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1635444444
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1635444444
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1635444444
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_93
timestamp 1635444444
transform 1 0 9660 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1635444444
transform 1 0 10212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1635444444
transform 1 0 9844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_19
timestamp 1635444444
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_7
timestamp 1635444444
transform 1 0 1748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1635444444
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1635444444
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1635444444
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1635444444
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1635444444
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1635444444
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1635444444
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1635444444
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1635444444
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1635444444
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1635444444
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1635444444
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1635444444
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1635444444
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1635444444
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1635444444
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1635444444
transform 1 0 9844 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1635444444
transform 1 0 9844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1635444444
transform 1 0 10212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1635444444
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_93
timestamp 1635444444
transform 1 0 9660 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1635444444
transform 1 0 9660 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1635444444
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_7
timestamp 1635444444
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1635444444
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1635444444
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1635444444
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1635444444
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1635444444
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1635444444
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1635444444
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1635444444
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1635444444
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_91
timestamp 1635444444
transform 1 0 9476 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_99
timestamp 1635444444
transform 1 0 10212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1635444444
transform 1 0 9844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1635444444
transform 1 0 9108 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_19
timestamp 1635444444
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_7
timestamp 1635444444
transform 1 0 1748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1635444444
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_31
timestamp 1635444444
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_43
timestamp 1635444444
transform 1 0 5060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1635444444
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1635444444
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_81
timestamp 1635444444
transform 1 0 8556 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1635444444
transform 1 0 8648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1635444444
transform 1 0 9200 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_86
timestamp 1635444444
transform 1 0 9016 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1635444444
transform 1 0 10212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _144_
timestamp 1635444444
transform 1 0 9384 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1635444444
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_7
timestamp 1635444444
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1635444444
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1635444444
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1635444444
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1635444444
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1635444444
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1635444444
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1635444444
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1635444444
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_91
timestamp 1635444444
transform 1 0 9476 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_99
timestamp 1635444444
transform 1 0 10212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1635444444
transform 1 0 9844 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1635444444
transform 1 0 9108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_19
timestamp 1635444444
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_7
timestamp 1635444444
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1635444444
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_31
timestamp 1635444444
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_43
timestamp 1635444444
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1635444444
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1635444444
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1635444444
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1635444444
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_93
timestamp 1635444444
transform 1 0 9660 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_99
timestamp 1635444444
transform 1 0 10212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1635444444
transform 1 0 9844 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 1635444444
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_7
timestamp 1635444444
transform 1 0 1748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1635444444
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1635444444
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1635444444
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1635444444
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1635444444
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1635444444
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1635444444
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1635444444
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1635444444
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1635444444
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1635444444
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1635444444
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1635444444
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1635444444
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1635444444
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_81
timestamp 1635444444
transform 1 0 8556 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _146_
timestamp 1635444444
transform 1 0 9384 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_89
timestamp 1635444444
transform 1 0 9292 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1635444444
transform 1 0 9660 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1635444444
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1635444444
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1635444444
transform 1 0 9844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1635444444
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_18
timestamp 1635444444
transform 1 0 2760 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1635444444
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635444444
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1635444444
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1635444444
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1635444444
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1635444444
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1635444444
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1635444444
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1635444444
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1635444444
transform 1 0 10212 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1635444444
transform 1 0 9200 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_101
timestamp 1635444444
transform 1 0 10396 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_90
timestamp 1635444444
transform 1 0 9384 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_98
timestamp 1635444444
transform 1 0 10120 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_18
timestamp 1635444444
transform 1 0 2760 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_6
timestamp 1635444444
transform 1 0 1656 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635444444
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_30
timestamp 1635444444
transform 1 0 3864 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_42
timestamp 1635444444
transform 1 0 4968 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1635444444
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1635444444
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_81
timestamp 1635444444
transform 1 0 8556 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1635444444
transform 1 0 8648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1635444444
transform 1 0 10212 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1635444444
transform 1 0 9200 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1635444444
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_86
timestamp 1635444444
transform 1 0 9016 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_90
timestamp 1635444444
transform 1 0 9384 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_98
timestamp 1635444444
transform 1 0 10120 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_10
timestamp 1635444444
transform 1 0 2024 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1635444444
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_6
timestamp 1635444444
transform 1 0 1656 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _048_
timestamp 1635444444
transform 1 0 2116 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1635444444
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1635444444
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1635444444
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1635444444
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1635444444
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1635444444
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1635444444
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _145_
timestamp 1635444444
transform 1 0 9384 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1635444444
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1635444444
transform 1 0 9016 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_13
timestamp 1635444444
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1635444444
transform 1 0 1380 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_57_25
timestamp 1635444444
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_37
timestamp 1635444444
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1635444444
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1635444444
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1635444444
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1635444444
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_81
timestamp 1635444444
transform 1 0 8556 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1635444444
transform 1 0 8648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1635444444
transform 1 0 9200 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_86
timestamp 1635444444
transform 1 0 9016 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_99
timestamp 1635444444
transform 1 0 10212 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 10856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _147_
timestamp 1635444444
transform 1 0 9384 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_58_13
timestamp 1635444444
transform 1 0 2300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1635444444
transform 1 0 1380 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_58_25
timestamp 1635444444
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1635444444
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1635444444
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1635444444
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1635444444
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1635444444
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1635444444
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_91
timestamp 1635444444
transform 1 0 9476 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_99
timestamp 1635444444
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1635444444
transform 1 0 9844 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1635444444
transform 1 0 9108 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_3
timestamp 1635444444
transform 1 0 1380 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1635444444
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_6
timestamp 1635444444
transform 1 0 1656 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _049_
timestamp 1635444444
transform 1 0 2024 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1635444444
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_23
timestamp 1635444444
transform 1 0 3220 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_35
timestamp 1635444444
transform 1 0 4324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1635444444
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1635444444
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1635444444
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_47
timestamp 1635444444
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1635444444
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1635444444
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1635444444
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1635444444
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_81
timestamp 1635444444
transform 1 0 8556 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1635444444
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1635444444
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1635444444
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1635444444
transform 1 0 9108 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _148_
timestamp 1635444444
transform 1 0 9384 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_91
timestamp 1635444444
transform 1 0 9476 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_87
timestamp 1635444444
transform 1 0 9108 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1635444444
transform 1 0 9200 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1635444444
transform 1 0 9844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1635444444
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_99
timestamp 1635444444
transform 1 0 10212 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1635444444
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1635444444
transform 1 0 1656 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635444444
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1635444444
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1635444444
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1635444444
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1635444444
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_81
timestamp 1635444444
transform 1 0 8556 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_91
timestamp 1635444444
transform 1 0 9476 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_99
timestamp 1635444444
transform 1 0 10212 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1635444444
transform 1 0 9844 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1635444444
transform 1 0 9108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_6
timestamp 1635444444
transform 1 0 1656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _082_
timestamp 1635444444
transform 1 0 2024 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635444444
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_22
timestamp 1635444444
transform 1 0 3128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1635444444
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1635444444
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1635444444
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1635444444
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1635444444
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1635444444
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_102
timestamp 1635444444
transform 1 0 10488 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_94
timestamp 1635444444
transform 1 0 9752 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 10856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _053_
timestamp 1635444444
transform 1 0 8924 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_63_13
timestamp 1635444444
transform 1 0 2300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1635444444
transform 1 0 1380 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_63_25
timestamp 1635444444
transform 1 0 3404 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_37
timestamp 1635444444
transform 1 0 4508 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 1635444444
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1635444444
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_73
timestamp 1635444444
transform 1 0 7820 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_78
timestamp 1635444444
transform 1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1635444444
transform 1 0 8648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1635444444
transform 1 0 7912 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1635444444
transform 1 0 9200 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1635444444
transform 1 0 10212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_101
timestamp 1635444444
transform 1 0 10396 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_86
timestamp 1635444444
transform 1 0 9016 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _149_
timestamp 1635444444
transform 1 0 9384 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_16
timestamp 1635444444
transform 1 0 2576 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _050_
timestamp 1635444444
transform 1 0 1748 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1635444444
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1635444444
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1635444444
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_65
timestamp 1635444444
transform 1 0 7084 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_73
timestamp 1635444444
transform 1 0 7820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1635444444
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1635444444
transform 1 0 8096 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_102
timestamp 1635444444
transform 1 0 10488 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1635444444
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_96
timestamp 1635444444
transform 1 0 9936 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _054_
timestamp 1635444444
transform 1 0 9108 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_19
timestamp 1635444444
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_7
timestamp 1635444444
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1635444444
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_31
timestamp 1635444444
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_43
timestamp 1635444444
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1635444444
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1635444444
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_69
timestamp 1635444444
transform 1 0 7452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_77
timestamp 1635444444
transform 1 0 8188 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_82
timestamp 1635444444
transform 1 0 8648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1635444444
transform 1 0 8280 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_95
timestamp 1635444444
transform 1 0 9844 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 10856 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _055_
timestamp 1635444444
transform 1 0 9016 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1635444444
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_7
timestamp 1635444444
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_19
timestamp 1635444444
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_7
timestamp 1635444444
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1635444444
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1635444444
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1635444444
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1635444444
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1635444444
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1635444444
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1635444444
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1635444444
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1635444444
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_65
timestamp 1635444444
transform 1 0 7084 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_73
timestamp 1635444444
transform 1 0 7820 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1635444444
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_69
timestamp 1635444444
transform 1 0 7452 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_77
timestamp 1635444444
transform 1 0 8188 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_82
timestamp 1635444444
transform 1 0 8648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1635444444
transform 1 0 8096 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1635444444
transform 1 0 8280 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_102
timestamp 1635444444
transform 1 0 10488 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_94
timestamp 1635444444
transform 1 0 9752 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_95
timestamp 1635444444
transform 1 0 9844 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _086_
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _088_
timestamp 1635444444
transform 1 0 9016 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_68_16
timestamp 1635444444
transform 1 0 2576 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1635444444
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _083_
timestamp 1635444444
transform 1 0 1748 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_68_29
timestamp 1635444444
transform 1 0 3772 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_37
timestamp 1635444444
transform 1 0 4508 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _051_
timestamp 1635444444
transform 1 0 4692 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_68_48
timestamp 1635444444
transform 1 0 5520 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_60
timestamp 1635444444
transform 1 0 6624 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_72
timestamp 1635444444
transform 1 0 7728 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_102
timestamp 1635444444
transform 1 0 10488 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_96
timestamp 1635444444
transform 1 0 9936 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 10856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _087_
timestamp 1635444444
transform 1 0 9108 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_69_13
timestamp 1635444444
transform 1 0 2300 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1635444444
transform 1 0 1380 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_69_25
timestamp 1635444444
transform 1 0 3404 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_37
timestamp 1635444444
transform 1 0 4508 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_49
timestamp 1635444444
transform 1 0 5612 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1635444444
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_57
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _052_
timestamp 1635444444
transform 1 0 6440 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_69_67
timestamp 1635444444
transform 1 0 7268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_79
timestamp 1635444444
transform 1 0 8372 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1635444444
transform 1 0 8464 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1635444444
transform 1 0 9200 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1635444444
transform 1 0 10212 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1635444444
transform 1 0 9016 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_101
timestamp 1635444444
transform 1 0 10396 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_84
timestamp 1635444444
transform 1 0 8832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _150_
timestamp 1635444444
transform 1 0 9384 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_11
timestamp 1635444444
transform 1 0 2116 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1635444444
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1635444444
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1635444444
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1635444444
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1635444444
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1635444444
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1635444444
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1635444444
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1635444444
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1635444444
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_85
timestamp 1635444444
transform 1 0 8924 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_91
timestamp 1635444444
transform 1 0 9476 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_99
timestamp 1635444444
transform 1 0 10212 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 10856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1635444444
transform 1 0 9844 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1635444444
transform 1 0 9108 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_11
timestamp 1635444444
transform 1 0 2116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1635444444
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1635444444
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_23
timestamp 1635444444
transform 1 0 3220 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_35
timestamp 1635444444
transform 1 0 4324 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_47
timestamp 1635444444
transform 1 0 5428 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1635444444
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1635444444
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1635444444
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_93
timestamp 1635444444
transform 1 0 9660 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_99
timestamp 1635444444
transform 1 0 10212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1635444444
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_19
timestamp 1635444444
transform 1 0 2852 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_7
timestamp 1635444444
transform 1 0 1748 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_19
timestamp 1635444444
transform 1 0 2852 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_7
timestamp 1635444444
transform 1 0 1748 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1635444444
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1635444444
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1635444444
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1635444444
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1635444444
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_31
timestamp 1635444444
transform 1 0 3956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _084_
timestamp 1635444444
transform 1 0 4692 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1635444444
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_48
timestamp 1635444444
transform 1 0 5520 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1635444444
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1635444444
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1635444444
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1635444444
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_81
timestamp 1635444444
transform 1 0 8556 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input160
timestamp 1635444444
transform 1 0 9108 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_91
timestamp 1635444444
transform 1 0 9476 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_85
timestamp 1635444444
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1635444444
transform 1 0 9844 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input122
timestamp 1635444444
transform 1 0 9844 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_99
timestamp 1635444444
transform 1 0 10212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_99
timestamp 1635444444
transform 1 0 10212 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_93
timestamp 1635444444
transform 1 0 9660 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 10856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 10856 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_19
timestamp 1635444444
transform 1 0 2852 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_7
timestamp 1635444444
transform 1 0 1748 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1635444444
transform 1 0 1380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1635444444
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1635444444
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1635444444
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_53
timestamp 1635444444
transform 1 0 5980 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_57
timestamp 1635444444
transform 1 0 6348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _085_
timestamp 1635444444
transform 1 0 6440 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_74_67
timestamp 1635444444
transform 1 0 7268 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_79
timestamp 1635444444
transform 1 0 8372 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1635444444
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1635444444
transform 1 0 9200 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1635444444
transform 1 0 10212 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1635444444
transform 1 0 9016 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_101
timestamp 1635444444
transform 1 0 10396 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_85
timestamp 1635444444
transform 1 0 8924 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _151_
timestamp 1635444444
transform 1 0 9384 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_11
timestamp 1635444444
transform 1 0 2116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1635444444
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1635444444
transform 1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_23
timestamp 1635444444
transform 1 0 3220 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_35
timestamp 1635444444
transform 1 0 4324 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_47
timestamp 1635444444
transform 1 0 5428 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1635444444
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1635444444
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_69
timestamp 1635444444
transform 1 0 7452 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_77
timestamp 1635444444
transform 1 0 8188 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_83
timestamp 1635444444
transform 1 0 8740 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1635444444
transform 1 0 8372 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1635444444
transform 1 0 9660 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_91
timestamp 1635444444
transform 1 0 9476 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_99
timestamp 1635444444
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input155
timestamp 1635444444
transform 1 0 9844 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1635444444
transform 1 0 9108 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1635444444
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1635444444
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1635444444
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1635444444
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _119_
timestamp 1635444444
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1635444444
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_65
timestamp 1635444444
transform 1 0 7084 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_80
timestamp 1635444444
transform 1 0 8464 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _056_
timestamp 1635444444
transform 1 0 7636 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_99
timestamp 1635444444
transform 1 0 10212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _122_
timestamp 1635444444
transform 1 0 9108 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_11
timestamp 1635444444
transform 1 0 2116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_3
timestamp 1635444444
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1635444444
transform 1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_23
timestamp 1635444444
transform 1 0 3220 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_35
timestamp 1635444444
transform 1 0 4324 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_47
timestamp 1635444444
transform 1 0 5428 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1635444444
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_69
timestamp 1635444444
transform 1 0 7452 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_77
timestamp 1635444444
transform 1 0 8188 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_83
timestamp 1635444444
transform 1 0 8740 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input157
timestamp 1635444444
transform 1 0 8372 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_99
timestamp 1635444444
transform 1 0 10212 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _123_
timestamp 1635444444
transform 1 0 9108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_11
timestamp 1635444444
transform 1 0 2116 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1635444444
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1635444444
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1635444444
transform 1 0 3220 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1635444444
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1635444444
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1635444444
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1635444444
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1635444444
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1635444444
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1635444444
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1635444444
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1635444444
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 10856 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _121_
timestamp 1635444444
transform 1 0 9108 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_19
timestamp 1635444444
transform 1 0 2852 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_7
timestamp 1635444444
transform 1 0 1748 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1635444444
transform 1 0 2116 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1635444444
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1635444444
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _160_
timestamp 1635444444
transform 1 0 2944 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1635444444
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1635444444
transform 1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_29
timestamp 1635444444
transform 1 0 3772 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_41
timestamp 1635444444
transform 1 0 4876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1635444444
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1635444444
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1635444444
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1635444444
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1635444444
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1635444444
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1635444444
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_81
timestamp 1635444444
transform 1 0 8556 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1635444444
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1635444444
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1635444444
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input158
timestamp 1635444444
transform 1 0 8648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _152_
timestamp 1635444444
transform 1 0 9384 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_89
timestamp 1635444444
transform 1 0 9292 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_85
timestamp 1635444444
transform 1 0 8924 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_90
timestamp 1635444444
transform 1 0 9384 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_86
timestamp 1635444444
transform 1 0 9016 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1635444444
transform 1 0 9200 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1635444444
transform -1 0 10856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 10856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_99
timestamp 1635444444
transform 1 0 10212 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_98
timestamp 1635444444
transform 1 0 10120 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_101
timestamp 1635444444
transform 1 0 10396 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1635444444
transform 1 0 10212 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1635444444
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1635444444
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1635444444
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1635444444
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _120_
timestamp 1635444444
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1635444444
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1635444444
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1635444444
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_69
timestamp 1635444444
transform 1 0 7452 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_75
timestamp 1635444444
transform 1 0 8004 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _089_
timestamp 1635444444
transform 1 0 8096 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_81_85
timestamp 1635444444
transform 1 0 8924 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_89
timestamp 1635444444
transform 1 0 9292 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1635444444
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1635444444
transform -1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 1635444444
transform 1 0 9384 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_82_11
timestamp 1635444444
transform 1 0 2116 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1635444444
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1635444444
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1635444444
transform 1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_23
timestamp 1635444444
transform 1 0 3220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1635444444
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1635444444
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1635444444
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1635444444
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1635444444
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_80
timestamp 1635444444
transform 1 0 8464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1635444444
transform 1 0 8188 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_85
timestamp 1635444444
transform 1 0 8924 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_89
timestamp 1635444444
transform 1 0 9292 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_99
timestamp 1635444444
transform 1 0 10212 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1635444444
transform -1 0 10856 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _163_
timestamp 1635444444
transform 1 0 9384 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_83_11
timestamp 1635444444
transform 1 0 2116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_3
timestamp 1635444444
transform 1 0 1380 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1635444444
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1635444444
transform 1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_23
timestamp 1635444444
transform 1 0 3220 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_35
timestamp 1635444444
transform 1 0 4324 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _161_
timestamp 1635444444
transform 1 0 4692 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_83_48
timestamp 1635444444
transform 1 0 5520 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1635444444
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1635444444
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_81
timestamp 1635444444
transform 1 0 8556 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1635444444
transform 1 0 8648 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_101
timestamp 1635444444
transform 1 0 10396 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_85
timestamp 1635444444
transform 1 0 8924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1635444444
transform -1 0 10856 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _164_
timestamp 1635444444
transform 1 0 9292 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1635444444
transform 1 0 10120 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1635444444
transform 1 0 9016 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_11
timestamp 1635444444
transform 1 0 2116 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_3
timestamp 1635444444
transform 1 0 1380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1635444444
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1635444444
transform 1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_23
timestamp 1635444444
transform 1 0 3220 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1635444444
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1635444444
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1635444444
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1635444444
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1635444444
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_80
timestamp 1635444444
transform 1 0 8464 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1635444444
transform 1 0 8188 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_84_102
timestamp 1635444444
transform 1 0 10488 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_85
timestamp 1635444444
transform 1 0 8924 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_98
timestamp 1635444444
transform 1 0 10120 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1635444444
transform -1 0 10856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _124_
timestamp 1635444444
transform 1 0 9016 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_11
timestamp 1635444444
transform 1 0 2116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_3
timestamp 1635444444
transform 1 0 1380 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_11
timestamp 1635444444
transform 1 0 2116 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_3
timestamp 1635444444
transform 1 0 1380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1635444444
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1635444444
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1635444444
transform 1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1635444444
transform 1 0 1748 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_23
timestamp 1635444444
transform 1 0 3220 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_35
timestamp 1635444444
transform 1 0 4324 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_23
timestamp 1635444444
transform 1 0 3220 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1635444444
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1635444444
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1635444444
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_47
timestamp 1635444444
transform 1 0 5428 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1635444444
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1635444444
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1635444444
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_69
timestamp 1635444444
transform 1 0 7452 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_75
timestamp 1635444444
transform 1 0 8004 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_79
timestamp 1635444444
transform 1 0 8372 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1635444444
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_80
timestamp 1635444444
transform 1 0 8464 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _125_
timestamp 1635444444
transform 1 0 8740 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1635444444
transform 1 0 8096 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1635444444
transform 1 0 8188 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_85_95
timestamp 1635444444
transform 1 0 9844 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_86_97
timestamp 1635444444
transform 1 0 10028 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1635444444
transform -1 0 10856 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1635444444
transform -1 0 10856 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _126_
timestamp 1635444444
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1635444444
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1635444444
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1635444444
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1635444444
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1635444444
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1635444444
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1635444444
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1635444444
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1635444444
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_81
timestamp 1635444444
transform 1 0 8556 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input123
timestamp 1635444444
transform 1 0 8648 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_86
timestamp 1635444444
transform 1 0 9016 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_99
timestamp 1635444444
transform 1 0 10212 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1635444444
transform -1 0 10856 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _153_
timestamp 1635444444
transform 1 0 9384 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_88_11
timestamp 1635444444
transform 1 0 2116 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_3
timestamp 1635444444
transform 1 0 1380 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1635444444
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1635444444
transform 1 0 1748 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_23
timestamp 1635444444
transform 1 0 3220 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1635444444
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1635444444
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1635444444
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1635444444
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_65
timestamp 1635444444
transform 1 0 7084 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_73
timestamp 1635444444
transform 1 0 7820 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_80
timestamp 1635444444
transform 1 0 8464 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input134
timestamp 1635444444
transform 1 0 8096 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_102
timestamp 1635444444
transform 1 0 10488 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_85
timestamp 1635444444
transform 1 0 8924 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_96
timestamp 1635444444
transform 1 0 9936 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1635444444
transform -1 0 10856 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _165_
timestamp 1635444444
transform 1 0 9108 0 1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_89_11
timestamp 1635444444
transform 1 0 2116 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_18
timestamp 1635444444
transform 1 0 2760 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_3
timestamp 1635444444
transform 1 0 1380 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1635444444
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1635444444
transform 1 0 2484 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1635444444
transform 1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_30
timestamp 1635444444
transform 1 0 3864 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_42
timestamp 1635444444
transform 1 0 4968 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_54
timestamp 1635444444
transform 1 0 6072 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1635444444
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1635444444
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_81
timestamp 1635444444
transform 1 0 8556 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1635444444
transform 1 0 8740 0 -1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_89_92
timestamp 1635444444
transform 1 0 9568 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_99
timestamp 1635444444
transform 1 0 10212 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1635444444
transform -1 0 10856 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1635444444
transform 1 0 9936 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_90_19
timestamp 1635444444
transform 1 0 2852 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_7
timestamp 1635444444
transform 1 0 1748 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1635444444
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1635444444
transform 1 0 1380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1635444444
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1635444444
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1635444444
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1635444444
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1635444444
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1635444444
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1635444444
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_102
timestamp 1635444444
transform 1 0 10488 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_94
timestamp 1635444444
transform 1 0 9752 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1635444444
transform -1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _167_
timestamp 1635444444
transform 1 0 8924 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_91_11
timestamp 1635444444
transform 1 0 2116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_3
timestamp 1635444444
transform 1 0 1380 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1635444444
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1635444444
transform 1 0 1748 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_23
timestamp 1635444444
transform 1 0 3220 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_35
timestamp 1635444444
transform 1 0 4324 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_47
timestamp 1635444444
transform 1 0 5428 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1635444444
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1635444444
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1635444444
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_81
timestamp 1635444444
transform 1 0 8556 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_91_91
timestamp 1635444444
transform 1 0 9476 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_99
timestamp 1635444444
transform 1 0 10212 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1635444444
transform -1 0 10856 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input145
timestamp 1635444444
transform 1 0 9844 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input149
timestamp 1635444444
transform 1 0 9108 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_14
timestamp 1635444444
transform 1 0 2392 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1635444444
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_19
timestamp 1635444444
transform 1 0 2852 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_7
timestamp 1635444444
transform 1 0 1748 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1635444444
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1635444444
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _061_
timestamp 1635444444
transform 1 0 1564 0 1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  output179
timestamp 1635444444
transform 1 0 2760 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1635444444
transform 1 0 1380 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_21
timestamp 1635444444
transform 1 0 3036 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1635444444
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1635444444
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1635444444
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_31
timestamp 1635444444
transform 1 0 3956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1635444444
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_43
timestamp 1635444444
transform 1 0 5060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1635444444
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1635444444
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1635444444
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1635444444
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1635444444
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1635444444
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_81
timestamp 1635444444
transform 1 0 8556 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input150
timestamp 1635444444
transform 1 0 9108 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _154_
timestamp 1635444444
transform 1 0 9384 0 -1 53312
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_89
timestamp 1635444444
transform 1 0 9292 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_91
timestamp 1635444444
transform 1 0 9476 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_85
timestamp 1635444444
transform 1 0 8924 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1635444444
transform 1 0 9660 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input148
timestamp 1635444444
transform 1 0 9844 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1635444444
transform -1 0 10856 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1635444444
transform -1 0 10856 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_99
timestamp 1635444444
transform 1 0 10212 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_99
timestamp 1635444444
transform 1 0 10212 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_19
timestamp 1635444444
transform 1 0 2852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_7
timestamp 1635444444
transform 1 0 1748 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1635444444
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1635444444
transform 1 0 1380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1635444444
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1635444444
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1635444444
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1635444444
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1635444444
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1635444444
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1635444444
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1635444444
transform 1 0 9660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_85
timestamp 1635444444
transform 1 0 8924 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_91
timestamp 1635444444
transform 1 0 9476 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_99
timestamp 1635444444
transform 1 0 10212 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1635444444
transform -1 0 10856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input151
timestamp 1635444444
transform 1 0 9844 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input154
timestamp 1635444444
transform 1 0 9108 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_17
timestamp 1635444444
transform 1 0 2668 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_3
timestamp 1635444444
transform 1 0 1380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_7
timestamp 1635444444
transform 1 0 1748 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1635444444
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _072_
timestamp 1635444444
transform 1 0 1840 0 -1 54400
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_95_29
timestamp 1635444444
transform 1 0 3772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_41
timestamp 1635444444
transform 1 0 4876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_53
timestamp 1635444444
transform 1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1635444444
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1635444444
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_81
timestamp 1635444444
transform 1 0 8556 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1635444444
transform 1 0 9660 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_91
timestamp 1635444444
transform 1 0 9476 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_99
timestamp 1635444444
transform 1 0 10212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1635444444
transform -1 0 10856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input152
timestamp 1635444444
transform 1 0 9844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1635444444
transform 1 0 9108 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_14
timestamp 1635444444
transform 1 0 2392 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_3
timestamp 1635444444
transform 1 0 1380 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1635444444
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _094_
timestamp 1635444444
transform 1 0 1564 0 1 54400
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_96_26
timestamp 1635444444
transform 1 0 3496 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1635444444
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1635444444
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1635444444
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1635444444
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1635444444
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1635444444
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_85
timestamp 1635444444
transform 1 0 8924 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_93
timestamp 1635444444
transform 1 0 9660 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_99
timestamp 1635444444
transform 1 0 10212 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1635444444
transform -1 0 10856 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1635444444
transform 1 0 9844 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_19
timestamp 1635444444
transform 1 0 2852 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_7
timestamp 1635444444
transform 1 0 1748 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1635444444
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1635444444
transform 1 0 1380 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_31
timestamp 1635444444
transform 1 0 3956 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_43
timestamp 1635444444
transform 1 0 5060 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1635444444
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1635444444
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1635444444
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1635444444
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_93
timestamp 1635444444
transform 1 0 9660 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_99
timestamp 1635444444
transform 1 0 10212 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1635444444
transform -1 0 10856 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input125
timestamp 1635444444
transform 1 0 9844 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_19
timestamp 1635444444
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_7
timestamp 1635444444
transform 1 0 1748 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1635444444
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1635444444
transform 1 0 1380 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1635444444
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1635444444
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1635444444
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1635444444
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1635444444
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1635444444
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1635444444
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1635444444
transform 1 0 9660 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_98_85
timestamp 1635444444
transform 1 0 8924 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_99
timestamp 1635444444
transform 1 0 10212 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1635444444
transform -1 0 10856 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input126
timestamp 1635444444
transform 1 0 9844 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_19
timestamp 1635444444
transform 1 0 2852 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_7
timestamp 1635444444
transform 1 0 1748 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_19
timestamp 1635444444
transform 1 0 2852 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_7
timestamp 1635444444
transform 1 0 1748 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1635444444
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1635444444
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1635444444
transform 1 0 1380 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1635444444
transform 1 0 1380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1635444444
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1635444444
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1635444444
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_31
timestamp 1635444444
transform 1 0 3956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1635444444
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_43
timestamp 1635444444
transform 1 0 5060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1635444444
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1635444444
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1635444444
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1635444444
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1635444444
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1635444444
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1635444444
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _155_
timestamp 1635444444
transform 1 0 9384 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_93
timestamp 1635444444
transform 1 0 9660 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_89
timestamp 1635444444
transform 1 0 9292 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_85
timestamp 1635444444
transform 1 0 8924 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input127
timestamp 1635444444
transform 1 0 9844 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1635444444
transform -1 0 10856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1635444444
transform -1 0 10856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_99
timestamp 1635444444
transform 1 0 10212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_99
timestamp 1635444444
transform 1 0 10212 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_19
timestamp 1635444444
transform 1 0 2852 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_7
timestamp 1635444444
transform 1 0 1748 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1635444444
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1635444444
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_31
timestamp 1635444444
transform 1 0 3956 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_43
timestamp 1635444444
transform 1 0 5060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1635444444
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1635444444
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1635444444
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_81
timestamp 1635444444
transform 1 0 8556 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_91
timestamp 1635444444
transform 1 0 9476 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_99
timestamp 1635444444
transform 1 0 10212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1635444444
transform -1 0 10856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input128
timestamp 1635444444
transform 1 0 9844 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1635444444
transform 1 0 9108 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_102_19
timestamp 1635444444
transform 1 0 2852 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_7
timestamp 1635444444
transform 1 0 1748 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1635444444
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1635444444
transform 1 0 1380 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1635444444
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1635444444
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1635444444
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1635444444
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1635444444
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1635444444
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1635444444
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1635444444
transform 1 0 9660 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_102_85
timestamp 1635444444
transform 1 0 8924 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_102_99
timestamp 1635444444
transform 1 0 10212 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1635444444
transform -1 0 10856 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1635444444
transform 1 0 9844 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_19
timestamp 1635444444
transform 1 0 2852 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_7
timestamp 1635444444
transform 1 0 1748 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1635444444
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1635444444
transform 1 0 1380 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_31
timestamp 1635444444
transform 1 0 3956 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_43
timestamp 1635444444
transform 1 0 5060 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1635444444
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1635444444
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1635444444
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1635444444
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_93
timestamp 1635444444
transform 1 0 9660 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_99
timestamp 1635444444
transform 1 0 10212 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1635444444
transform -1 0 10856 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1635444444
transform 1 0 9844 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1635444444
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1635444444
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1635444444
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1635444444
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1635444444
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1635444444
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1635444444
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1635444444
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1635444444
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1635444444
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_85
timestamp 1635444444
transform 1 0 8924 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_104_93
timestamp 1635444444
transform 1 0 9660 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_104_99
timestamp 1635444444
transform 1 0 10212 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1635444444
transform -1 0 10856 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input132
timestamp 1635444444
transform 1 0 9844 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_11
timestamp 1635444444
transform 1 0 2116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_3
timestamp 1635444444
transform 1 0 1380 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_11
timestamp 1635444444
transform 1 0 2116 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_3
timestamp 1635444444
transform 1 0 1380 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1635444444
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1635444444
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1635444444
transform 1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1635444444
transform 1 0 1748 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_23
timestamp 1635444444
transform 1 0 3220 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_35
timestamp 1635444444
transform 1 0 4324 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_23
timestamp 1635444444
transform 1 0 3220 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1635444444
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1635444444
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1635444444
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_47
timestamp 1635444444
transform 1 0 5428 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1635444444
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1635444444
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1635444444
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1635444444
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_81
timestamp 1635444444
transform 1 0 8556 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_106_65
timestamp 1635444444
transform 1 0 7084 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_106_80
timestamp 1635444444
transform 1 0 8464 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _066_
timestamp 1635444444
transform 1 0 7636 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input136
timestamp 1635444444
transform 1 0 9108 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_85
timestamp 1635444444
transform 1 0 8924 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_105_91
timestamp 1635444444
transform 1 0 9476 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input135
timestamp 1635444444
transform 1 0 9844 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1635444444
transform 1 0 9844 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_99
timestamp 1635444444
transform 1 0 10212 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_93
timestamp 1635444444
transform 1 0 9660 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_99
timestamp 1635444444
transform 1 0 10212 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1635444444
transform -1 0 10856 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1635444444
transform -1 0 10856 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_13
timestamp 1635444444
transform 1 0 2300 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_3
timestamp 1635444444
transform 1 0 1380 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1635444444
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _073_
timestamp 1635444444
transform 1 0 1472 0 -1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1635444444
transform 1 0 2668 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_21
timestamp 1635444444
transform 1 0 3036 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_33
timestamp 1635444444
transform 1 0 4140 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_45
timestamp 1635444444
transform 1 0 5244 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_53
timestamp 1635444444
transform 1 0 5980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1635444444
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1635444444
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input137
timestamp 1635444444
transform 1 0 8556 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_85
timestamp 1635444444
transform 1 0 8924 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_99
timestamp 1635444444
transform 1 0 10212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1635444444
transform -1 0 10856 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input138
timestamp 1635444444
transform 1 0 9292 0 -1 60928
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_108_3
timestamp 1635444444
transform 1 0 1380 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1635444444
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _062_
timestamp 1635444444
transform 1 0 1932 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_21
timestamp 1635444444
transform 1 0 3036 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1635444444
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1635444444
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1635444444
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1635444444
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1635444444
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1635444444
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1635444444
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_85
timestamp 1635444444
transform 1 0 8924 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_99
timestamp 1635444444
transform 1 0 10212 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1635444444
transform -1 0 10856 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _156_
timestamp 1635444444
transform 1 0 9108 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_11
timestamp 1635444444
transform 1 0 2116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_3
timestamp 1635444444
transform 1 0 1380 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1635444444
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1635444444
transform 1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_23
timestamp 1635444444
transform 1 0 3220 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_35
timestamp 1635444444
transform 1 0 4324 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_47
timestamp 1635444444
transform 1 0 5428 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1635444444
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1635444444
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1635444444
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_81
timestamp 1635444444
transform 1 0 8556 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_109_99
timestamp 1635444444
transform 1 0 10212 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1635444444
transform -1 0 10856 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input139
timestamp 1635444444
transform 1 0 9292 0 -1 62016
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_110_11
timestamp 1635444444
transform 1 0 2116 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_3
timestamp 1635444444
transform 1 0 1380 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1635444444
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1635444444
transform 1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_23
timestamp 1635444444
transform 1 0 3220 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1635444444
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1635444444
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1635444444
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1635444444
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_65
timestamp 1635444444
transform 1 0 7084 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_110_80
timestamp 1635444444
transform 1 0 8464 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp 1635444444
transform 1 0 7636 0 1 62016
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_110_85
timestamp 1635444444
transform 1 0 8924 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_99
timestamp 1635444444
transform 1 0 10212 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1635444444
transform -1 0 10856 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input140
timestamp 1635444444
transform 1 0 9292 0 1 62016
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_111_18
timestamp 1635444444
transform 1 0 2760 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_3
timestamp 1635444444
transform 1 0 1380 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1635444444
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _095_
timestamp 1635444444
transform 1 0 1932 0 -1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_111_30
timestamp 1635444444
transform 1 0 3864 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_42
timestamp 1635444444
transform 1 0 4968 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_54
timestamp 1635444444
transform 1 0 6072 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_111_57
timestamp 1635444444
transform 1 0 6348 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_111_65
timestamp 1635444444
transform 1 0 7084 0 -1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_111_76
timestamp 1635444444
transform 1 0 8096 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_82
timestamp 1635444444
transform 1 0 8648 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _058_
timestamp 1635444444
transform 1 0 8740 0 -1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _059_
timestamp 1635444444
transform 1 0 7268 0 -1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_111_92
timestamp 1635444444
transform 1 0 9568 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_99
timestamp 1635444444
transform 1 0 10212 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1635444444
transform -1 0 10856 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1635444444
transform 1 0 9936 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_112_7
timestamp 1635444444
transform 1 0 1748 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_19
timestamp 1635444444
transform 1 0 2852 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_7
timestamp 1635444444
transform 1 0 1748 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1635444444
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1635444444
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _067_
timestamp 1635444444
transform 1 0 2484 0 1 63104
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1635444444
transform 1 0 1380 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input61
timestamp 1635444444
transform 1 0 1380 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_24
timestamp 1635444444
transform 1 0 3312 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_29
timestamp 1635444444
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_41
timestamp 1635444444
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_31
timestamp 1635444444
transform 1 0 3956 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_53
timestamp 1635444444
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_43
timestamp 1635444444
transform 1 0 5060 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1635444444
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1635444444
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_65
timestamp 1635444444
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1635444444
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1635444444
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1635444444
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_81
timestamp 1635444444
transform 1 0 8556 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp 1635444444
transform 1 0 8740 0 -1 64192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_112_85
timestamp 1635444444
transform 1 0 8924 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1635444444
transform 1 0 9292 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_113_92
timestamp 1635444444
transform 1 0 9568 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_92
timestamp 1635444444
transform 1 0 9568 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1635444444
transform 1 0 9936 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1635444444
transform 1 0 9936 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_113_99
timestamp 1635444444
transform 1 0 10212 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_99
timestamp 1635444444
transform 1 0 10212 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1635444444
transform -1 0 10856 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1635444444
transform -1 0 10856 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_114_19
timestamp 1635444444
transform 1 0 2852 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_7
timestamp 1635444444
transform 1 0 1748 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1635444444
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1635444444
transform 1 0 1380 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1635444444
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1635444444
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1635444444
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1635444444
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1635444444
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1635444444
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1635444444
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_114_85
timestamp 1635444444
transform 1 0 8924 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_114_99
timestamp 1635444444
transform 1 0 10212 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1635444444
transform -1 0 10856 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _157_
timestamp 1635444444
transform 1 0 9108 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_11
timestamp 1635444444
transform 1 0 2116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_3
timestamp 1635444444
transform 1 0 1380 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1635444444
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1635444444
transform 1 0 1748 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_23
timestamp 1635444444
transform 1 0 3220 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_35
timestamp 1635444444
transform 1 0 4324 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_47
timestamp 1635444444
transform 1 0 5428 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1635444444
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_57
timestamp 1635444444
transform 1 0 6348 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_115_65
timestamp 1635444444
transform 1 0 7084 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_115_76
timestamp 1635444444
transform 1 0 8096 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_80
timestamp 1635444444
transform 1 0 8464 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _092_
timestamp 1635444444
transform 1 0 7268 0 -1 65280
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1635444444
transform 1 0 8556 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_84
timestamp 1635444444
transform 1 0 8832 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_91
timestamp 1635444444
transform 1 0 9476 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_99
timestamp 1635444444
transform 1 0 10212 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1635444444
transform -1 0 10856 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1635444444
transform 1 0 9200 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1635444444
transform 1 0 9844 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_13
timestamp 1635444444
transform 1 0 2300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_6
timestamp 1635444444
transform 1 0 1656 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1635444444
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1635444444
transform 1 0 1380 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635444444
transform 1 0 2024 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_116_25
timestamp 1635444444
transform 1 0 3404 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_29
timestamp 1635444444
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_41
timestamp 1635444444
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_53
timestamp 1635444444
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_65
timestamp 1635444444
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1635444444
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1635444444
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_116_85
timestamp 1635444444
transform 1 0 8924 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_116_99
timestamp 1635444444
transform 1 0 10212 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1635444444
transform -1 0 10856 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _158_
timestamp 1635444444
transform 1 0 9108 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_15
timestamp 1635444444
transform 1 0 2484 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1635444444
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _060_
timestamp 1635444444
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _100_
timestamp 1635444444
transform 1 0 2852 0 -1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_117_28
timestamp 1635444444
transform 1 0 3680 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_40
timestamp 1635444444
transform 1 0 4784 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_52
timestamp 1635444444
transform 1 0 5888 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1635444444
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1635444444
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_81
timestamp 1635444444
transform 1 0 8556 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_117_91
timestamp 1635444444
transform 1 0 9476 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_99
timestamp 1635444444
transform 1 0 10212 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1635444444
transform -1 0 10856 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1635444444
transform 1 0 9844 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1635444444
transform 1 0 9108 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_118_19
timestamp 1635444444
transform 1 0 2852 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_118_3
timestamp 1635444444
transform 1 0 1380 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_12
timestamp 1635444444
transform 1 0 2208 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_19
timestamp 1635444444
transform 1 0 2852 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1635444444
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1635444444
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _068_
timestamp 1635444444
transform 1 0 1748 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _093_
timestamp 1635444444
transform 1 0 1380 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1635444444
transform 1 0 2576 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1635444444
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1635444444
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1635444444
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_31
timestamp 1635444444
transform 1 0 3956 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_53
timestamp 1635444444
transform 1 0 5980 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_61
timestamp 1635444444
transform 1 0 6716 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_43
timestamp 1635444444
transform 1 0 5060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1635444444
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1635444444
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _063_
timestamp 1635444444
transform 1 0 6808 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_74
timestamp 1635444444
transform 1 0 7912 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_118_82
timestamp 1635444444
transform 1 0 8648 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_119_69
timestamp 1635444444
transform 1 0 7452 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_77
timestamp 1635444444
transform 1 0 8188 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 1635444444
transform 1 0 8648 0 -1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1635444444
transform 1 0 8280 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_119_91
timestamp 1635444444
transform 1 0 9476 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_118_85
timestamp 1635444444
transform 1 0 8924 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1635444444
transform 1 0 9660 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1635444444
transform 1 0 9844 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1635444444
transform -1 0 10856 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1635444444
transform -1 0 10856 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_99
timestamp 1635444444
transform 1 0 10212 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_99
timestamp 1635444444
transform 1 0 10212 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _057_
timestamp 1635444444
transform 1 0 9108 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_13
timestamp 1635444444
transform 1 0 2300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1635444444
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1635444444
transform 1 0 1380 0 1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_120_25
timestamp 1635444444
transform 1 0 3404 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1635444444
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1635444444
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1635444444
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_65
timestamp 1635444444
transform 1 0 7084 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_73
timestamp 1635444444
transform 1 0 7820 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_80
timestamp 1635444444
transform 1 0 8464 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output280
timestamp 1635444444
transform 1 0 8096 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_102
timestamp 1635444444
transform 1 0 10488 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_85
timestamp 1635444444
transform 1 0 8924 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_98
timestamp 1635444444
transform 1 0 10120 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1635444444
transform -1 0 10856 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _065_
timestamp 1635444444
transform 1 0 9292 0 1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_121_18
timestamp 1635444444
transform 1 0 2760 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_6
timestamp 1635444444
transform 1 0 1656 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1635444444
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform 1 0 1380 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_121_22
timestamp 1635444444
transform 1 0 3128 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_35
timestamp 1635444444
transform 1 0 4324 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _070_
timestamp 1635444444
transform 1 0 3220 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_47
timestamp 1635444444
transform 1 0 5428 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1635444444
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1635444444
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1635444444
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1635444444
transform 1 0 8556 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1635444444
transform 1 0 9108 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_121_85
timestamp 1635444444
transform 1 0 8924 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_121_89
timestamp 1635444444
transform 1 0 9292 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_121_99
timestamp 1635444444
transform 1 0 10212 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1635444444
transform -1 0 10856 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _064_
timestamp 1635444444
transform 1 0 9384 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_122_6
timestamp 1635444444
transform 1 0 1656 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1635444444
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _077_
timestamp 1635444444
transform 1 0 2208 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1635444444
transform 1 0 1380 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_24
timestamp 1635444444
transform 1 0 3312 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1635444444
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1635444444
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_53
timestamp 1635444444
transform 1 0 5980 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_61
timestamp 1635444444
transform 1 0 6716 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _096_
timestamp 1635444444
transform 1 0 6808 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_122_71
timestamp 1635444444
transform 1 0 7636 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_75
timestamp 1635444444
transform 1 0 8004 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_80
timestamp 1635444444
transform 1 0 8464 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output283
timestamp 1635444444
transform 1 0 8096 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1635444444
transform -1 0 10396 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1635444444
transform -1 0 9384 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_122_101
timestamp 1635444444
transform 1 0 10396 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_122_85
timestamp 1635444444
transform 1 0 8924 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_90
timestamp 1635444444
transform 1 0 9384 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_98
timestamp 1635444444
transform 1 0 10120 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1635444444
transform -1 0 10856 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_13
timestamp 1635444444
transform 1 0 2300 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_3
timestamp 1635444444
transform 1 0 1380 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1635444444
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _076_
timestamp 1635444444
transform 1 0 2668 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp 1635444444
transform 1 0 1472 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_123_29
timestamp 1635444444
transform 1 0 3772 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_41
timestamp 1635444444
transform 1 0 4876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_53
timestamp 1635444444
transform 1 0 5980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1635444444
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_69
timestamp 1635444444
transform 1 0 7452 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_123_77
timestamp 1635444444
transform 1 0 8188 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_123_83
timestamp 1635444444
transform 1 0 8740 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output284
timestamp 1635444444
transform 1 0 8372 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1635444444
transform -1 0 10856 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _098_
timestamp 1635444444
transform 1 0 9384 0 -1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1635444444
transform 1 0 10212 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1635444444
transform 1 0 9016 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_15
timestamp 1635444444
transform 1 0 2484 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1635444444
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _071_
timestamp 1635444444
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635444444
transform 1 0 2852 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_124_22
timestamp 1635444444
transform 1 0 3128 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_124_32
timestamp 1635444444
transform 1 0 4048 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform 1 0 3772 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_44
timestamp 1635444444
transform 1 0 5152 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_56
timestamp 1635444444
transform 1 0 6256 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_68
timestamp 1635444444
transform 1 0 7360 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_80
timestamp 1635444444
transform 1 0 8464 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1635444444
transform -1 0 9384 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_124_85
timestamp 1635444444
transform 1 0 8924 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_99
timestamp 1635444444
transform 1 0 10212 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1635444444
transform -1 0 10856 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _097_
timestamp 1635444444
transform 1 0 9384 0 1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_125_3
timestamp 1635444444
transform 1 0 1380 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_126_13
timestamp 1635444444
transform 1 0 2300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1635444444
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1635444444
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _074_
timestamp 1635444444
transform 1 0 1932 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1635444444
transform 1 0 1380 0 1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_125_21
timestamp 1635444444
transform 1 0 3036 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_33
timestamp 1635444444
transform 1 0 4140 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_126_25
timestamp 1635444444
transform 1 0 3404 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_126_38
timestamp 1635444444
transform 1 0 4600 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _103_
timestamp 1635444444
transform 1 0 3772 0 1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_125_45
timestamp 1635444444
transform 1 0 5244 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_53
timestamp 1635444444
transform 1 0 5980 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_125_57
timestamp 1635444444
transform 1 0 6348 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_50
timestamp 1635444444
transform 1 0 5704 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_62
timestamp 1635444444
transform 1 0 6808 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_77
timestamp 1635444444
transform 1 0 8188 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_126_74
timestamp 1635444444
transform 1 0 7912 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_126_82
timestamp 1635444444
transform 1 0 8648 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_4  _069_
timestamp 1635444444
transform 1 0 7084 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_126_85
timestamp 1635444444
transform 1 0 8924 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_125_90
timestamp 1635444444
transform 1 0 9384 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_85
timestamp 1635444444
transform 1 0 8924 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1635444444
transform 1 0 9200 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1635444444
transform 1 0 9844 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_126_99
timestamp 1635444444
transform 1 0 10212 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_126_93
timestamp 1635444444
transform 1 0 9660 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_125_98
timestamp 1635444444
transform 1 0 10120 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_125_101
timestamp 1635444444
transform 1 0 10396 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1635444444
transform 1 0 10212 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1635444444
transform -1 0 10856 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1635444444
transform -1 0 10856 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_18
timestamp 1635444444
transform 1 0 2760 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_6
timestamp 1635444444
transform 1 0 1656 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1635444444
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform 1 0 1380 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_30
timestamp 1635444444
transform 1 0 3864 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_42
timestamp 1635444444
transform 1 0 4968 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_54
timestamp 1635444444
transform 1 0 6072 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1635444444
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1635444444
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1635444444
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_93
timestamp 1635444444
transform 1 0 9660 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_127_99
timestamp 1635444444
transform 1 0 10212 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1635444444
transform -1 0 10856 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1635444444
transform 1 0 9844 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_128_13
timestamp 1635444444
transform 1 0 2300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_128_6
timestamp 1635444444
transform 1 0 1656 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1635444444
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform 1 0 1380 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1635444444
transform 1 0 2024 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_128_25
timestamp 1635444444
transform 1 0 3404 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1635444444
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  _075_
timestamp 1635444444
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_53
timestamp 1635444444
transform 1 0 5980 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _079_
timestamp 1635444444
transform 1 0 6072 0 1 71808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_128_63
timestamp 1635444444
transform 1 0 6900 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_75
timestamp 1635444444
transform 1 0 8004 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1635444444
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1635444444
transform 1 0 9660 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_128_85
timestamp 1635444444
transform 1 0 8924 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_128_91
timestamp 1635444444
transform 1 0 9476 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_128_99
timestamp 1635444444
transform 1 0 10212 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1635444444
transform -1 0 10856 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1635444444
transform 1 0 9844 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1635444444
transform 1 0 9108 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_12
timestamp 1635444444
transform 1 0 2208 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1635444444
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _104_
timestamp 1635444444
transform 1 0 1380 0 -1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 1635444444
transform 1 0 2576 0 -1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_129_25
timestamp 1635444444
transform 1 0 3404 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_37
timestamp 1635444444
transform 1 0 4508 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_49
timestamp 1635444444
transform 1 0 5612 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1635444444
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1635444444
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1635444444
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_81
timestamp 1635444444
transform 1 0 8556 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_129_91
timestamp 1635444444
transform 1 0 9476 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_99
timestamp 1635444444
transform 1 0 10212 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1635444444
transform -1 0 10856 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1635444444
transform 1 0 9844 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1635444444
transform 1 0 9108 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_130_13
timestamp 1635444444
transform 1 0 2300 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_130_20
timestamp 1635444444
transform 1 0 2944 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_3
timestamp 1635444444
transform 1 0 1380 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1635444444
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _106_
timestamp 1635444444
transform 1 0 1472 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1635444444
transform 1 0 2668 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1635444444
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1635444444
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1635444444
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_74
timestamp 1635444444
transform 1 0 7912 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_130_82
timestamp 1635444444
transform 1 0 8648 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp 1635444444
transform 1 0 7084 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_130_85
timestamp 1635444444
transform 1 0 8924 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_89
timestamp 1635444444
transform 1 0 9292 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_130_99
timestamp 1635444444
transform 1 0 10212 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1635444444
transform -1 0 10856 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _078_
timestamp 1635444444
transform 1 0 9384 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_131_14
timestamp 1635444444
transform 1 0 2392 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_131_3
timestamp 1635444444
transform 1 0 1380 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1635444444
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _105_
timestamp 1635444444
transform 1 0 1564 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_131_22
timestamp 1635444444
transform 1 0 3128 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_131_33
timestamp 1635444444
transform 1 0 4140 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _108_
timestamp 1635444444
transform 1 0 3312 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_131_45
timestamp 1635444444
transform 1 0 5244 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_131_53
timestamp 1635444444
transform 1 0 5980 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1635444444
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1635444444
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_81
timestamp 1635444444
transform 1 0 8556 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_131_91
timestamp 1635444444
transform 1 0 9476 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_131_99
timestamp 1635444444
transform 1 0 10212 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1635444444
transform -1 0 10856 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1635444444
transform 1 0 9844 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1635444444
transform 1 0 9108 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform 1 0 1380 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _107_
timestamp 1635444444
transform 1 0 1932 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1635444444
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1635444444
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_133_6
timestamp 1635444444
transform 1 0 1656 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_132_3
timestamp 1635444444
transform 1 0 1380 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform 1 0 2024 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _109_
timestamp 1635444444
transform 1 0 2668 0 -1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_133_13
timestamp 1635444444
transform 1 0 2300 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_132_18
timestamp 1635444444
transform 1 0 2760 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_132_26
timestamp 1635444444
transform 1 0 3496 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_132_29
timestamp 1635444444
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_41
timestamp 1635444444
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_26
timestamp 1635444444
transform 1 0 3496 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_38
timestamp 1635444444
transform 1 0 4600 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_132_53
timestamp 1635444444
transform 1 0 5980 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_133_50
timestamp 1635444444
transform 1 0 5704 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1635444444
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 1635444444
transform 1 0 6072 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_132_63
timestamp 1635444444
transform 1 0 6900 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_75
timestamp 1635444444
transform 1 0 8004 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1635444444
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1635444444
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1635444444
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _111_
timestamp 1635444444
transform 1 0 9384 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_133_93
timestamp 1635444444
transform 1 0 9660 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_132_89
timestamp 1635444444
transform 1 0 9292 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_132_85
timestamp 1635444444
transform 1 0 8924 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1635444444
transform 1 0 9844 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1635444444
transform -1 0 10856 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1635444444
transform -1 0 10856 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_133_99
timestamp 1635444444
transform 1 0 10212 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_132_99
timestamp 1635444444
transform 1 0 10212 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_134_11
timestamp 1635444444
transform 1 0 2116 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_3
timestamp 1635444444
transform 1 0 1380 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1635444444
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1635444444
transform 1 0 1748 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_134_23
timestamp 1635444444
transform 1 0 3220 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1635444444
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1635444444
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1635444444
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1635444444
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1635444444
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1635444444
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1635444444
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_85
timestamp 1635444444
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_134_93
timestamp 1635444444
transform 1 0 9660 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_134_99
timestamp 1635444444
transform 1 0 10212 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1635444444
transform -1 0 10856 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1635444444
transform 1 0 9844 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_13
timestamp 1635444444
transform 1 0 2300 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1635444444
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1635444444
transform 1 0 1380 0 -1 76160
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_135_25
timestamp 1635444444
transform 1 0 3404 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_37
timestamp 1635444444
transform 1 0 4508 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_49
timestamp 1635444444
transform 1 0 5612 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1635444444
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1635444444
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1635444444
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_81
timestamp 1635444444
transform 1 0 8556 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_135_91
timestamp 1635444444
transform 1 0 9476 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_135_99
timestamp 1635444444
transform 1 0 10212 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1635444444
transform -1 0 10856 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1635444444
transform 1 0 9844 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1635444444
transform 1 0 9108 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_136_18
timestamp 1635444444
transform 1 0 2760 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_6
timestamp 1635444444
transform 1 0 1656 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1635444444
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform 1 0 1380 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_136_26
timestamp 1635444444
transform 1 0 3496 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_136_29
timestamp 1635444444
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_41
timestamp 1635444444
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_53
timestamp 1635444444
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_65
timestamp 1635444444
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1635444444
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1635444444
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_136_85
timestamp 1635444444
transform 1 0 8924 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_136_91
timestamp 1635444444
transform 1 0 9476 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_136_99
timestamp 1635444444
transform 1 0 10212 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1635444444
transform -1 0 10856 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1635444444
transform 1 0 9844 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1635444444
transform 1 0 9108 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_13
timestamp 1635444444
transform 1 0 2300 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_20
timestamp 1635444444
transform 1 0 2944 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_6
timestamp 1635444444
transform 1 0 1656 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1635444444
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform 1 0 1380 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform 1 0 2024 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1635444444
transform 1 0 2668 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_32
timestamp 1635444444
transform 1 0 4048 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_44
timestamp 1635444444
transform 1 0 5152 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1635444444
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_69
timestamp 1635444444
transform 1 0 7452 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_137_77
timestamp 1635444444
transform 1 0 8188 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_137_83
timestamp 1635444444
transform 1 0 8740 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1635444444
transform 1 0 8372 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_91
timestamp 1635444444
transform 1 0 9476 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_99
timestamp 1635444444
transform 1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1635444444
transform -1 0 10856 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1635444444
transform 1 0 9844 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1635444444
transform 1 0 9108 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_13
timestamp 1635444444
transform 1 0 2300 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_138_20
timestamp 1635444444
transform 1 0 2944 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1635444444
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform 1 0 2668 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1635444444
transform 1 0 1380 0 1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_138_29
timestamp 1635444444
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_41
timestamp 1635444444
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_138_53
timestamp 1635444444
transform 1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_138_57
timestamp 1635444444
transform 1 0 6348 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_138_65
timestamp 1635444444
transform 1 0 7084 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_72
timestamp 1635444444
transform 1 0 7728 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_80
timestamp 1635444444
transform 1 0 8464 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1635444444
transform 1 0 8096 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1635444444
transform 1 0 7360 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_138_85
timestamp 1635444444
transform 1 0 8924 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_138_91
timestamp 1635444444
transform 1 0 9476 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_99
timestamp 1635444444
transform 1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1635444444
transform -1 0 10856 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1635444444
transform 1 0 9844 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1635444444
transform 1 0 9108 0 1 77248
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 4904 800 5024 6 ram_addr0[0]
port 0 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 ram_addr0[1]
port 1 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 ram_addr0[2]
port 2 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 ram_addr0[3]
port 3 nsew signal tristate
rlabel metal3 s 0 7488 800 7608 6 ram_addr0[4]
port 4 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 ram_addr0[5]
port 5 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 ram_addr0[6]
port 6 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 ram_addr0[7]
port 7 nsew signal tristate
rlabel metal3 s 0 53728 800 53848 6 ram_addr1[0]
port 8 nsew signal tristate
rlabel metal3 s 0 54408 800 54528 6 ram_addr1[1]
port 9 nsew signal tristate
rlabel metal3 s 0 55088 800 55208 6 ram_addr1[2]
port 10 nsew signal tristate
rlabel metal3 s 0 55768 800 55888 6 ram_addr1[3]
port 11 nsew signal tristate
rlabel metal3 s 0 56448 800 56568 6 ram_addr1[4]
port 12 nsew signal tristate
rlabel metal3 s 0 56992 800 57112 6 ram_addr1[5]
port 13 nsew signal tristate
rlabel metal3 s 0 57672 800 57792 6 ram_addr1[6]
port 14 nsew signal tristate
rlabel metal3 s 0 58352 800 58472 6 ram_addr1[7]
port 15 nsew signal tristate
rlabel metal3 s 0 280 800 400 6 ram_clk0
port 16 nsew signal tristate
rlabel metal3 s 0 52368 800 52488 6 ram_clk1
port 17 nsew signal tristate
rlabel metal3 s 0 824 800 944 6 ram_csb0
port 18 nsew signal tristate
rlabel metal3 s 0 53048 800 53168 6 ram_csb1
port 19 nsew signal tristate
rlabel metal3 s 0 10072 800 10192 6 ram_din0[0]
port 20 nsew signal tristate
rlabel metal3 s 0 16736 800 16856 6 ram_din0[10]
port 21 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 ram_din0[11]
port 22 nsew signal tristate
rlabel metal3 s 0 18096 800 18216 6 ram_din0[12]
port 23 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 ram_din0[13]
port 24 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 ram_din0[14]
port 25 nsew signal tristate
rlabel metal3 s 0 20000 800 20120 6 ram_din0[15]
port 26 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 ram_din0[16]
port 27 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 ram_din0[17]
port 28 nsew signal tristate
rlabel metal3 s 0 22040 800 22160 6 ram_din0[18]
port 29 nsew signal tristate
rlabel metal3 s 0 22720 800 22840 6 ram_din0[19]
port 30 nsew signal tristate
rlabel metal3 s 0 10752 800 10872 6 ram_din0[1]
port 31 nsew signal tristate
rlabel metal3 s 0 23400 800 23520 6 ram_din0[20]
port 32 nsew signal tristate
rlabel metal3 s 0 23944 800 24064 6 ram_din0[21]
port 33 nsew signal tristate
rlabel metal3 s 0 24624 800 24744 6 ram_din0[22]
port 34 nsew signal tristate
rlabel metal3 s 0 25304 800 25424 6 ram_din0[23]
port 35 nsew signal tristate
rlabel metal3 s 0 25984 800 26104 6 ram_din0[24]
port 36 nsew signal tristate
rlabel metal3 s 0 26664 800 26784 6 ram_din0[25]
port 37 nsew signal tristate
rlabel metal3 s 0 27344 800 27464 6 ram_din0[26]
port 38 nsew signal tristate
rlabel metal3 s 0 28024 800 28144 6 ram_din0[27]
port 39 nsew signal tristate
rlabel metal3 s 0 28568 800 28688 6 ram_din0[28]
port 40 nsew signal tristate
rlabel metal3 s 0 29248 800 29368 6 ram_din0[29]
port 41 nsew signal tristate
rlabel metal3 s 0 11432 800 11552 6 ram_din0[2]
port 42 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 ram_din0[30]
port 43 nsew signal tristate
rlabel metal3 s 0 30608 800 30728 6 ram_din0[31]
port 44 nsew signal tristate
rlabel metal3 s 0 12112 800 12232 6 ram_din0[3]
port 45 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 ram_din0[4]
port 46 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 ram_din0[5]
port 47 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 ram_din0[6]
port 48 nsew signal tristate
rlabel metal3 s 0 14696 800 14816 6 ram_din0[7]
port 49 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 ram_din0[8]
port 50 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 ram_din0[9]
port 51 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 ram_dout0[0]
port 52 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 ram_dout0[10]
port 53 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 ram_dout0[11]
port 54 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 ram_dout0[12]
port 55 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 ram_dout0[13]
port 56 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 ram_dout0[14]
port 57 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 ram_dout0[15]
port 58 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 ram_dout0[16]
port 59 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 ram_dout0[17]
port 60 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 ram_dout0[18]
port 61 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 ram_dout0[19]
port 62 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 ram_dout0[1]
port 63 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 ram_dout0[20]
port 64 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 ram_dout0[21]
port 65 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 ram_dout0[22]
port 66 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 ram_dout0[23]
port 67 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 ram_dout0[24]
port 68 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 ram_dout0[25]
port 69 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 ram_dout0[26]
port 70 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 ram_dout0[27]
port 71 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 ram_dout0[28]
port 72 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 ram_dout0[29]
port 73 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 ram_dout0[2]
port 74 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 ram_dout0[30]
port 75 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 ram_dout0[31]
port 76 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 ram_dout0[3]
port 77 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 ram_dout0[4]
port 78 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 ram_dout0[5]
port 79 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 ram_dout0[6]
port 80 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 ram_dout0[7]
port 81 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 ram_dout0[8]
port 82 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 ram_dout0[9]
port 83 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 ram_dout1[0]
port 84 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 ram_dout1[10]
port 85 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 ram_dout1[11]
port 86 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 ram_dout1[12]
port 87 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 ram_dout1[13]
port 88 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 ram_dout1[14]
port 89 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 ram_dout1[15]
port 90 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 ram_dout1[16]
port 91 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 ram_dout1[17]
port 92 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 ram_dout1[18]
port 93 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 ram_dout1[19]
port 94 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 ram_dout1[1]
port 95 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 ram_dout1[20]
port 96 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 ram_dout1[21]
port 97 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 ram_dout1[22]
port 98 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 ram_dout1[23]
port 99 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 ram_dout1[24]
port 100 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 ram_dout1[25]
port 101 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 ram_dout1[26]
port 102 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 ram_dout1[27]
port 103 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 ram_dout1[28]
port 104 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 ram_dout1[29]
port 105 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 ram_dout1[2]
port 106 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 ram_dout1[30]
port 107 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 ram_dout1[31]
port 108 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 ram_dout1[3]
port 109 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 ram_dout1[4]
port 110 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 ram_dout1[5]
port 111 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 ram_dout1[6]
port 112 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 ram_dout1[7]
port 113 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 ram_dout1[8]
port 114 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 ram_dout1[9]
port 115 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 ram_web0
port 116 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 ram_wmask0[0]
port 117 nsew signal tristate
rlabel metal3 s 0 2864 800 2984 6 ram_wmask0[1]
port 118 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 ram_wmask0[2]
port 119 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 ram_wmask0[3]
port 120 nsew signal tristate
rlabel metal4 s 2575 2128 2895 77840 6 vccd1
port 121 nsew power input
rlabel metal4 s 5839 2128 6159 77840 6 vccd1
port 121 nsew power input
rlabel metal4 s 9103 2128 9423 77840 6 vccd1
port 121 nsew power input
rlabel metal4 s 4207 2128 4527 77840 6 vssd1
port 122 nsew ground input
rlabel metal4 s 7471 2128 7791 77840 6 vssd1
port 122 nsew ground input
rlabel metal3 s 11200 552 12000 672 6 wb_a_clk_i
port 123 nsew signal input
rlabel metal3 s 11200 960 12000 1080 6 wb_a_rst_i
port 124 nsew signal input
rlabel metal3 s 11200 40264 12000 40384 6 wb_b_clk_i
port 125 nsew signal input
rlabel metal3 s 11200 40808 12000 40928 6 wb_b_rst_i
port 126 nsew signal input
rlabel metal3 s 11200 2864 12000 2984 6 wbs_a_ack_o
port 127 nsew signal tristate
rlabel metal3 s 11200 5312 12000 5432 6 wbs_a_adr_i[0]
port 128 nsew signal input
rlabel metal3 s 11200 5720 12000 5840 6 wbs_a_adr_i[1]
port 129 nsew signal input
rlabel metal3 s 11200 6264 12000 6384 6 wbs_a_adr_i[2]
port 130 nsew signal input
rlabel metal3 s 11200 6672 12000 6792 6 wbs_a_adr_i[3]
port 131 nsew signal input
rlabel metal3 s 11200 7216 12000 7336 6 wbs_a_adr_i[4]
port 132 nsew signal input
rlabel metal3 s 11200 7624 12000 7744 6 wbs_a_adr_i[5]
port 133 nsew signal input
rlabel metal3 s 11200 8168 12000 8288 6 wbs_a_adr_i[6]
port 134 nsew signal input
rlabel metal3 s 11200 8576 12000 8696 6 wbs_a_adr_i[7]
port 135 nsew signal input
rlabel metal3 s 11200 9120 12000 9240 6 wbs_a_adr_i[8]
port 136 nsew signal input
rlabel metal3 s 11200 9528 12000 9648 6 wbs_a_adr_i[9]
port 137 nsew signal input
rlabel metal3 s 11200 1912 12000 2032 6 wbs_a_cyc_i
port 138 nsew signal input
rlabel metal3 s 11200 10072 12000 10192 6 wbs_a_dat_i[0]
port 139 nsew signal input
rlabel metal3 s 11200 14696 12000 14816 6 wbs_a_dat_i[10]
port 140 nsew signal input
rlabel metal3 s 11200 15240 12000 15360 6 wbs_a_dat_i[11]
port 141 nsew signal input
rlabel metal3 s 11200 15648 12000 15768 6 wbs_a_dat_i[12]
port 142 nsew signal input
rlabel metal3 s 11200 16192 12000 16312 6 wbs_a_dat_i[13]
port 143 nsew signal input
rlabel metal3 s 11200 16600 12000 16720 6 wbs_a_dat_i[14]
port 144 nsew signal input
rlabel metal3 s 11200 17144 12000 17264 6 wbs_a_dat_i[15]
port 145 nsew signal input
rlabel metal3 s 11200 17552 12000 17672 6 wbs_a_dat_i[16]
port 146 nsew signal input
rlabel metal3 s 11200 18096 12000 18216 6 wbs_a_dat_i[17]
port 147 nsew signal input
rlabel metal3 s 11200 18504 12000 18624 6 wbs_a_dat_i[18]
port 148 nsew signal input
rlabel metal3 s 11200 19048 12000 19168 6 wbs_a_dat_i[19]
port 149 nsew signal input
rlabel metal3 s 11200 10480 12000 10600 6 wbs_a_dat_i[1]
port 150 nsew signal input
rlabel metal3 s 11200 19456 12000 19576 6 wbs_a_dat_i[20]
port 151 nsew signal input
rlabel metal3 s 11200 20000 12000 20120 6 wbs_a_dat_i[21]
port 152 nsew signal input
rlabel metal3 s 11200 20408 12000 20528 6 wbs_a_dat_i[22]
port 153 nsew signal input
rlabel metal3 s 11200 20952 12000 21072 6 wbs_a_dat_i[23]
port 154 nsew signal input
rlabel metal3 s 11200 21360 12000 21480 6 wbs_a_dat_i[24]
port 155 nsew signal input
rlabel metal3 s 11200 21904 12000 22024 6 wbs_a_dat_i[25]
port 156 nsew signal input
rlabel metal3 s 11200 22312 12000 22432 6 wbs_a_dat_i[26]
port 157 nsew signal input
rlabel metal3 s 11200 22856 12000 22976 6 wbs_a_dat_i[27]
port 158 nsew signal input
rlabel metal3 s 11200 23264 12000 23384 6 wbs_a_dat_i[28]
port 159 nsew signal input
rlabel metal3 s 11200 23672 12000 23792 6 wbs_a_dat_i[29]
port 160 nsew signal input
rlabel metal3 s 11200 11024 12000 11144 6 wbs_a_dat_i[2]
port 161 nsew signal input
rlabel metal3 s 11200 24216 12000 24336 6 wbs_a_dat_i[30]
port 162 nsew signal input
rlabel metal3 s 11200 24624 12000 24744 6 wbs_a_dat_i[31]
port 163 nsew signal input
rlabel metal3 s 11200 11432 12000 11552 6 wbs_a_dat_i[3]
port 164 nsew signal input
rlabel metal3 s 11200 11840 12000 11960 6 wbs_a_dat_i[4]
port 165 nsew signal input
rlabel metal3 s 11200 12384 12000 12504 6 wbs_a_dat_i[5]
port 166 nsew signal input
rlabel metal3 s 11200 12792 12000 12912 6 wbs_a_dat_i[6]
port 167 nsew signal input
rlabel metal3 s 11200 13336 12000 13456 6 wbs_a_dat_i[7]
port 168 nsew signal input
rlabel metal3 s 11200 13744 12000 13864 6 wbs_a_dat_i[8]
port 169 nsew signal input
rlabel metal3 s 11200 14288 12000 14408 6 wbs_a_dat_i[9]
port 170 nsew signal input
rlabel metal3 s 11200 25168 12000 25288 6 wbs_a_dat_o[0]
port 171 nsew signal tristate
rlabel metal3 s 11200 29928 12000 30048 6 wbs_a_dat_o[10]
port 172 nsew signal tristate
rlabel metal3 s 11200 30336 12000 30456 6 wbs_a_dat_o[11]
port 173 nsew signal tristate
rlabel metal3 s 11200 30880 12000 31000 6 wbs_a_dat_o[12]
port 174 nsew signal tristate
rlabel metal3 s 11200 31288 12000 31408 6 wbs_a_dat_o[13]
port 175 nsew signal tristate
rlabel metal3 s 11200 31832 12000 31952 6 wbs_a_dat_o[14]
port 176 nsew signal tristate
rlabel metal3 s 11200 32240 12000 32360 6 wbs_a_dat_o[15]
port 177 nsew signal tristate
rlabel metal3 s 11200 32784 12000 32904 6 wbs_a_dat_o[16]
port 178 nsew signal tristate
rlabel metal3 s 11200 33192 12000 33312 6 wbs_a_dat_o[17]
port 179 nsew signal tristate
rlabel metal3 s 11200 33736 12000 33856 6 wbs_a_dat_o[18]
port 180 nsew signal tristate
rlabel metal3 s 11200 34144 12000 34264 6 wbs_a_dat_o[19]
port 181 nsew signal tristate
rlabel metal3 s 11200 25576 12000 25696 6 wbs_a_dat_o[1]
port 182 nsew signal tristate
rlabel metal3 s 11200 34552 12000 34672 6 wbs_a_dat_o[20]
port 183 nsew signal tristate
rlabel metal3 s 11200 35096 12000 35216 6 wbs_a_dat_o[21]
port 184 nsew signal tristate
rlabel metal3 s 11200 35504 12000 35624 6 wbs_a_dat_o[22]
port 185 nsew signal tristate
rlabel metal3 s 11200 36048 12000 36168 6 wbs_a_dat_o[23]
port 186 nsew signal tristate
rlabel metal3 s 11200 36456 12000 36576 6 wbs_a_dat_o[24]
port 187 nsew signal tristate
rlabel metal3 s 11200 37000 12000 37120 6 wbs_a_dat_o[25]
port 188 nsew signal tristate
rlabel metal3 s 11200 37408 12000 37528 6 wbs_a_dat_o[26]
port 189 nsew signal tristate
rlabel metal3 s 11200 37952 12000 38072 6 wbs_a_dat_o[27]
port 190 nsew signal tristate
rlabel metal3 s 11200 38360 12000 38480 6 wbs_a_dat_o[28]
port 191 nsew signal tristate
rlabel metal3 s 11200 38904 12000 39024 6 wbs_a_dat_o[29]
port 192 nsew signal tristate
rlabel metal3 s 11200 26120 12000 26240 6 wbs_a_dat_o[2]
port 193 nsew signal tristate
rlabel metal3 s 11200 39312 12000 39432 6 wbs_a_dat_o[30]
port 194 nsew signal tristate
rlabel metal3 s 11200 39856 12000 39976 6 wbs_a_dat_o[31]
port 195 nsew signal tristate
rlabel metal3 s 11200 26528 12000 26648 6 wbs_a_dat_o[3]
port 196 nsew signal tristate
rlabel metal3 s 11200 27072 12000 27192 6 wbs_a_dat_o[4]
port 197 nsew signal tristate
rlabel metal3 s 11200 27480 12000 27600 6 wbs_a_dat_o[5]
port 198 nsew signal tristate
rlabel metal3 s 11200 28024 12000 28144 6 wbs_a_dat_o[6]
port 199 nsew signal tristate
rlabel metal3 s 11200 28432 12000 28552 6 wbs_a_dat_o[7]
port 200 nsew signal tristate
rlabel metal3 s 11200 28976 12000 29096 6 wbs_a_dat_o[8]
port 201 nsew signal tristate
rlabel metal3 s 11200 29384 12000 29504 6 wbs_a_dat_o[9]
port 202 nsew signal tristate
rlabel metal3 s 11200 3408 12000 3528 6 wbs_a_sel_i[0]
port 203 nsew signal input
rlabel metal3 s 11200 3816 12000 3936 6 wbs_a_sel_i[1]
port 204 nsew signal input
rlabel metal3 s 11200 4360 12000 4480 6 wbs_a_sel_i[2]
port 205 nsew signal input
rlabel metal3 s 11200 4768 12000 4888 6 wbs_a_sel_i[3]
port 206 nsew signal input
rlabel metal3 s 11200 1504 12000 1624 6 wbs_a_stb_i
port 207 nsew signal input
rlabel metal3 s 11200 2456 12000 2576 6 wbs_a_we_i
port 208 nsew signal input
rlabel metal3 s 11200 42712 12000 42832 6 wbs_b_ack_o
port 209 nsew signal tristate
rlabel metal3 s 11200 45024 12000 45144 6 wbs_b_adr_i[0]
port 210 nsew signal input
rlabel metal3 s 11200 45568 12000 45688 6 wbs_b_adr_i[1]
port 211 nsew signal input
rlabel metal3 s 11200 45976 12000 46096 6 wbs_b_adr_i[2]
port 212 nsew signal input
rlabel metal3 s 11200 46384 12000 46504 6 wbs_b_adr_i[3]
port 213 nsew signal input
rlabel metal3 s 11200 46928 12000 47048 6 wbs_b_adr_i[4]
port 214 nsew signal input
rlabel metal3 s 11200 47336 12000 47456 6 wbs_b_adr_i[5]
port 215 nsew signal input
rlabel metal3 s 11200 47880 12000 48000 6 wbs_b_adr_i[6]
port 216 nsew signal input
rlabel metal3 s 11200 48288 12000 48408 6 wbs_b_adr_i[7]
port 217 nsew signal input
rlabel metal3 s 11200 48832 12000 48952 6 wbs_b_adr_i[8]
port 218 nsew signal input
rlabel metal3 s 11200 49240 12000 49360 6 wbs_b_adr_i[9]
port 219 nsew signal input
rlabel metal3 s 11200 41760 12000 41880 6 wbs_b_cyc_i
port 220 nsew signal input
rlabel metal3 s 11200 49784 12000 49904 6 wbs_b_dat_i[0]
port 221 nsew signal input
rlabel metal3 s 11200 54544 12000 54664 6 wbs_b_dat_i[10]
port 222 nsew signal input
rlabel metal3 s 11200 54952 12000 55072 6 wbs_b_dat_i[11]
port 223 nsew signal input
rlabel metal3 s 11200 55496 12000 55616 6 wbs_b_dat_i[12]
port 224 nsew signal input
rlabel metal3 s 11200 55904 12000 56024 6 wbs_b_dat_i[13]
port 225 nsew signal input
rlabel metal3 s 11200 56448 12000 56568 6 wbs_b_dat_i[14]
port 226 nsew signal input
rlabel metal3 s 11200 56856 12000 56976 6 wbs_b_dat_i[15]
port 227 nsew signal input
rlabel metal3 s 11200 57264 12000 57384 6 wbs_b_dat_i[16]
port 228 nsew signal input
rlabel metal3 s 11200 57808 12000 57928 6 wbs_b_dat_i[17]
port 229 nsew signal input
rlabel metal3 s 11200 58216 12000 58336 6 wbs_b_dat_i[18]
port 230 nsew signal input
rlabel metal3 s 11200 58760 12000 58880 6 wbs_b_dat_i[19]
port 231 nsew signal input
rlabel metal3 s 11200 50192 12000 50312 6 wbs_b_dat_i[1]
port 232 nsew signal input
rlabel metal3 s 11200 59168 12000 59288 6 wbs_b_dat_i[20]
port 233 nsew signal input
rlabel metal3 s 11200 59712 12000 59832 6 wbs_b_dat_i[21]
port 234 nsew signal input
rlabel metal3 s 11200 60120 12000 60240 6 wbs_b_dat_i[22]
port 235 nsew signal input
rlabel metal3 s 11200 60664 12000 60784 6 wbs_b_dat_i[23]
port 236 nsew signal input
rlabel metal3 s 11200 61072 12000 61192 6 wbs_b_dat_i[24]
port 237 nsew signal input
rlabel metal3 s 11200 61616 12000 61736 6 wbs_b_dat_i[25]
port 238 nsew signal input
rlabel metal3 s 11200 62024 12000 62144 6 wbs_b_dat_i[26]
port 239 nsew signal input
rlabel metal3 s 11200 62568 12000 62688 6 wbs_b_dat_i[27]
port 240 nsew signal input
rlabel metal3 s 11200 62976 12000 63096 6 wbs_b_dat_i[28]
port 241 nsew signal input
rlabel metal3 s 11200 63520 12000 63640 6 wbs_b_dat_i[29]
port 242 nsew signal input
rlabel metal3 s 11200 50736 12000 50856 6 wbs_b_dat_i[2]
port 243 nsew signal input
rlabel metal3 s 11200 63928 12000 64048 6 wbs_b_dat_i[30]
port 244 nsew signal input
rlabel metal3 s 11200 64472 12000 64592 6 wbs_b_dat_i[31]
port 245 nsew signal input
rlabel metal3 s 11200 51144 12000 51264 6 wbs_b_dat_i[3]
port 246 nsew signal input
rlabel metal3 s 11200 51688 12000 51808 6 wbs_b_dat_i[4]
port 247 nsew signal input
rlabel metal3 s 11200 52096 12000 52216 6 wbs_b_dat_i[5]
port 248 nsew signal input
rlabel metal3 s 11200 52640 12000 52760 6 wbs_b_dat_i[6]
port 249 nsew signal input
rlabel metal3 s 11200 53048 12000 53168 6 wbs_b_dat_i[7]
port 250 nsew signal input
rlabel metal3 s 11200 53592 12000 53712 6 wbs_b_dat_i[8]
port 251 nsew signal input
rlabel metal3 s 11200 54000 12000 54120 6 wbs_b_dat_i[9]
port 252 nsew signal input
rlabel metal3 s 11200 64880 12000 65000 6 wbs_b_dat_o[0]
port 253 nsew signal tristate
rlabel metal3 s 11200 69640 12000 69760 6 wbs_b_dat_o[10]
port 254 nsew signal tristate
rlabel metal3 s 11200 70048 12000 70168 6 wbs_b_dat_o[11]
port 255 nsew signal tristate
rlabel metal3 s 11200 70592 12000 70712 6 wbs_b_dat_o[12]
port 256 nsew signal tristate
rlabel metal3 s 11200 71000 12000 71120 6 wbs_b_dat_o[13]
port 257 nsew signal tristate
rlabel metal3 s 11200 71544 12000 71664 6 wbs_b_dat_o[14]
port 258 nsew signal tristate
rlabel metal3 s 11200 71952 12000 72072 6 wbs_b_dat_o[15]
port 259 nsew signal tristate
rlabel metal3 s 11200 72496 12000 72616 6 wbs_b_dat_o[16]
port 260 nsew signal tristate
rlabel metal3 s 11200 72904 12000 73024 6 wbs_b_dat_o[17]
port 261 nsew signal tristate
rlabel metal3 s 11200 73448 12000 73568 6 wbs_b_dat_o[18]
port 262 nsew signal tristate
rlabel metal3 s 11200 73856 12000 73976 6 wbs_b_dat_o[19]
port 263 nsew signal tristate
rlabel metal3 s 11200 65424 12000 65544 6 wbs_b_dat_o[1]
port 264 nsew signal tristate
rlabel metal3 s 11200 74400 12000 74520 6 wbs_b_dat_o[20]
port 265 nsew signal tristate
rlabel metal3 s 11200 74808 12000 74928 6 wbs_b_dat_o[21]
port 266 nsew signal tristate
rlabel metal3 s 11200 75352 12000 75472 6 wbs_b_dat_o[22]
port 267 nsew signal tristate
rlabel metal3 s 11200 75760 12000 75880 6 wbs_b_dat_o[23]
port 268 nsew signal tristate
rlabel metal3 s 11200 76304 12000 76424 6 wbs_b_dat_o[24]
port 269 nsew signal tristate
rlabel metal3 s 11200 76712 12000 76832 6 wbs_b_dat_o[25]
port 270 nsew signal tristate
rlabel metal3 s 11200 77256 12000 77376 6 wbs_b_dat_o[26]
port 271 nsew signal tristate
rlabel metal3 s 11200 77664 12000 77784 6 wbs_b_dat_o[27]
port 272 nsew signal tristate
rlabel metal3 s 11200 78208 12000 78328 6 wbs_b_dat_o[28]
port 273 nsew signal tristate
rlabel metal3 s 11200 78616 12000 78736 6 wbs_b_dat_o[29]
port 274 nsew signal tristate
rlabel metal3 s 11200 65832 12000 65952 6 wbs_b_dat_o[2]
port 275 nsew signal tristate
rlabel metal3 s 11200 79160 12000 79280 6 wbs_b_dat_o[30]
port 276 nsew signal tristate
rlabel metal3 s 11200 79568 12000 79688 6 wbs_b_dat_o[31]
port 277 nsew signal tristate
rlabel metal3 s 11200 66376 12000 66496 6 wbs_b_dat_o[3]
port 278 nsew signal tristate
rlabel metal3 s 11200 66784 12000 66904 6 wbs_b_dat_o[4]
port 279 nsew signal tristate
rlabel metal3 s 11200 67328 12000 67448 6 wbs_b_dat_o[5]
port 280 nsew signal tristate
rlabel metal3 s 11200 67736 12000 67856 6 wbs_b_dat_o[6]
port 281 nsew signal tristate
rlabel metal3 s 11200 68280 12000 68400 6 wbs_b_dat_o[7]
port 282 nsew signal tristate
rlabel metal3 s 11200 68688 12000 68808 6 wbs_b_dat_o[8]
port 283 nsew signal tristate
rlabel metal3 s 11200 69096 12000 69216 6 wbs_b_dat_o[9]
port 284 nsew signal tristate
rlabel metal3 s 11200 43120 12000 43240 6 wbs_b_sel_i[0]
port 285 nsew signal input
rlabel metal3 s 11200 43664 12000 43784 6 wbs_b_sel_i[1]
port 286 nsew signal input
rlabel metal3 s 11200 44072 12000 44192 6 wbs_b_sel_i[2]
port 287 nsew signal input
rlabel metal3 s 11200 44616 12000 44736 6 wbs_b_sel_i[3]
port 288 nsew signal input
rlabel metal3 s 11200 41216 12000 41336 6 wbs_b_stb_i
port 289 nsew signal input
rlabel metal3 s 11200 42168 12000 42288 6 wbs_b_we_i
port 290 nsew signal input
rlabel metal3 s 11200 144 12000 264 6 writable_port_req
port 291 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
<< end >>
