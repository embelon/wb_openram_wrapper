magic
tech sky130A
magscale 1 2
timestamp 1635332841
<< locali >>
rect 6929 52139 6963 55709
rect 7389 55217 7423 56321
rect 7389 55183 7515 55217
rect 6929 36567 6963 51357
rect 7021 36635 7055 53533
rect 6929 36533 7055 36567
rect 6929 34051 6963 36465
rect 6929 30923 6963 33881
rect 7021 28475 7055 36533
rect 7113 28679 7147 50881
rect 6929 24395 6963 27625
rect 7021 23035 7055 27285
rect 7113 24939 7147 28373
rect 7205 27047 7239 51969
rect 7297 38743 7331 54621
rect 7389 47175 7423 50201
rect 7481 47243 7515 55183
rect 7573 51077 7607 55641
rect 7757 51077 7791 53125
rect 7573 51043 7699 51077
rect 7757 51043 7883 51077
rect 7389 47141 7515 47175
rect 7297 32011 7331 37145
rect 7297 28747 7331 31841
rect 7389 28815 7423 47005
rect 7481 42279 7515 47141
rect 7481 41531 7515 42109
rect 7481 38811 7515 41383
rect 7573 41259 7607 46461
rect 7665 40579 7699 51043
rect 7757 46767 7791 49861
rect 7757 41531 7791 46597
rect 7849 41327 7883 51043
rect 7941 41667 7975 54213
rect 7941 41395 7975 41497
rect 7757 41293 7883 41327
rect 7481 38777 7607 38811
rect 7481 30311 7515 38709
rect 7573 35071 7607 38777
rect 7665 36227 7699 40409
rect 7757 37315 7791 41293
rect 7573 31875 7607 33813
rect 7389 25959 7423 28645
rect 7481 25415 7515 28441
rect 7573 25483 7607 30141
rect 7665 26503 7699 34493
rect 7757 32963 7791 37145
rect 7849 29699 7883 41157
rect 7941 37179 7975 41225
rect 6963 23001 7055 23035
rect 6929 18955 6963 22049
rect 6929 16779 6963 17493
rect 7021 16711 7055 22933
rect 7113 21131 7147 23613
rect 7205 20043 7239 23681
rect 7757 23239 7791 28781
rect 7941 27591 7975 36601
rect 7297 17867 7331 21981
rect 6929 16677 7055 16711
rect 6929 16577 6963 16677
rect 6929 16543 7055 16577
rect 6929 11883 6963 14977
rect 6929 8823 6963 10013
rect 7021 8007 7055 16543
rect 7389 15147 7423 23137
rect 6929 6987 6963 7905
rect 6929 4131 6963 6613
rect 7021 5967 7055 7837
rect 7113 7055 7147 8925
rect 7113 4811 7147 6885
rect 7205 4743 7239 11237
rect 7297 6919 7331 14773
<< viali >>
rect 2329 57545 2363 57579
rect 3065 57545 3099 57579
rect 4261 57545 4295 57579
rect 4997 57545 5031 57579
rect 1409 57409 1443 57443
rect 2145 57409 2179 57443
rect 2881 57409 2915 57443
rect 4077 57409 4111 57443
rect 4813 57409 4847 57443
rect 5549 57409 5583 57443
rect 1593 57205 1627 57239
rect 5733 57205 5767 57239
rect 4537 57001 4571 57035
rect 5273 57001 5307 57035
rect 6009 57001 6043 57035
rect 1409 56797 1443 56831
rect 4353 56797 4387 56831
rect 5089 56797 5123 56831
rect 5825 56797 5859 56831
rect 1593 56661 1627 56695
rect 1593 56457 1627 56491
rect 1409 56321 1443 56355
rect 5549 56321 5583 56355
rect 7389 56321 7423 56355
rect 5733 56185 5767 56219
rect 4261 55913 4295 55947
rect 1409 55709 1443 55743
rect 4445 55709 4479 55743
rect 5825 55709 5859 55743
rect 6929 55709 6963 55743
rect 1593 55573 1627 55607
rect 6009 55573 6043 55607
rect 2145 55369 2179 55403
rect 2973 55369 3007 55403
rect 4077 55369 4111 55403
rect 4721 55369 4755 55403
rect 1409 55233 1443 55267
rect 2329 55233 2363 55267
rect 3157 55233 3191 55267
rect 4261 55233 4295 55267
rect 4905 55233 4939 55267
rect 5365 55233 5399 55267
rect 5549 55233 5583 55267
rect 5733 55097 5767 55131
rect 1593 55029 1627 55063
rect 2145 54825 2179 54859
rect 3801 54825 3835 54859
rect 1409 54621 1443 54655
rect 2329 54621 2363 54655
rect 3985 54621 4019 54655
rect 5825 54621 5859 54655
rect 1593 54485 1627 54519
rect 6009 54485 6043 54519
rect 3249 54281 3283 54315
rect 4905 54281 4939 54315
rect 3433 54145 3467 54179
rect 5089 54145 5123 54179
rect 5549 54145 5583 54179
rect 5733 54009 5767 54043
rect 1409 53533 1443 53567
rect 5733 53533 5767 53567
rect 5825 53533 5859 53567
rect 1593 53397 1627 53431
rect 6009 53397 6043 53431
rect 3433 53193 3467 53227
rect 1409 53057 1443 53091
rect 3617 53057 3651 53091
rect 5549 53057 5583 53091
rect 1593 52853 1627 52887
rect 5365 52853 5399 52887
rect 5733 52853 5767 52887
rect 3065 52649 3099 52683
rect 3249 52445 3283 52479
rect 5825 52445 5859 52479
rect 6009 52309 6043 52343
rect 7573 55641 7607 55675
rect 7297 54621 7331 54655
rect 3525 52105 3559 52139
rect 6929 52105 6963 52139
rect 7021 53533 7055 53567
rect 1409 51969 1443 52003
rect 3709 51969 3743 52003
rect 5549 51969 5583 52003
rect 1593 51833 1627 51867
rect 5733 51765 5767 51799
rect 1409 51357 1443 51391
rect 5733 51357 5767 51391
rect 5825 51357 5859 51391
rect 6929 51357 6963 51391
rect 1593 51221 1627 51255
rect 6009 51221 6043 51255
rect 2145 51017 2179 51051
rect 2789 51017 2823 51051
rect 1409 50881 1443 50915
rect 2329 50881 2363 50915
rect 2973 50881 3007 50915
rect 5549 50881 5583 50915
rect 1593 50677 1627 50711
rect 5733 50677 5767 50711
rect 1593 50473 1627 50507
rect 1777 50269 1811 50303
rect 5825 50269 5859 50303
rect 6009 50133 6043 50167
rect 2145 49929 2179 49963
rect 1409 49793 1443 49827
rect 2329 49793 2363 49827
rect 5549 49793 5583 49827
rect 5365 49725 5399 49759
rect 1593 49589 1627 49623
rect 5733 49589 5767 49623
rect 1409 49181 1443 49215
rect 5825 49181 5859 49215
rect 1593 49045 1627 49079
rect 6009 49045 6043 49079
rect 5549 48705 5583 48739
rect 5365 48501 5399 48535
rect 5733 48501 5767 48535
rect 3801 48229 3835 48263
rect 1409 48093 1443 48127
rect 3249 48093 3283 48127
rect 3985 48093 4019 48127
rect 5825 48093 5859 48127
rect 1593 47957 1627 47991
rect 3065 47957 3099 47991
rect 6009 47957 6043 47991
rect 1409 47617 1443 47651
rect 5549 47617 5583 47651
rect 5457 47481 5491 47515
rect 1593 47413 1627 47447
rect 5733 47413 5767 47447
rect 3801 47209 3835 47243
rect 1409 47005 1443 47039
rect 3985 47005 4019 47039
rect 5733 47005 5767 47039
rect 5825 47005 5859 47039
rect 1593 46869 1627 46903
rect 6009 46869 6043 46903
rect 2789 46665 2823 46699
rect 4169 46665 4203 46699
rect 2973 46529 3007 46563
rect 4353 46529 4387 46563
rect 5549 46529 5583 46563
rect 5733 46325 5767 46359
rect 1409 45917 1443 45951
rect 5825 45917 5859 45951
rect 1593 45781 1627 45815
rect 6009 45781 6043 45815
rect 1409 45441 1443 45475
rect 5549 45441 5583 45475
rect 1593 45237 1627 45271
rect 5365 45237 5399 45271
rect 5733 45237 5767 45271
rect 2329 45033 2363 45067
rect 2513 44829 2547 44863
rect 5825 44829 5859 44863
rect 6009 44693 6043 44727
rect 1409 44353 1443 44387
rect 5549 44353 5583 44387
rect 1593 44217 1627 44251
rect 5733 44149 5767 44183
rect 1409 43741 1443 43775
rect 5825 43741 5859 43775
rect 1593 43605 1627 43639
rect 6009 43605 6043 43639
rect 1409 43265 1443 43299
rect 5549 43265 5583 43299
rect 1593 43061 1627 43095
rect 5733 43061 5767 43095
rect 2145 42313 2179 42347
rect 1409 42177 1443 42211
rect 2329 42177 2363 42211
rect 5549 42177 5583 42211
rect 1593 42041 1627 42075
rect 5733 42041 5767 42075
rect 5457 41973 5491 42007
rect 3065 41769 3099 41803
rect 4353 41769 4387 41803
rect 5549 41633 5583 41667
rect 1409 41565 1443 41599
rect 3249 41565 3283 41599
rect 5273 41565 5307 41599
rect 4261 41497 4295 41531
rect 1593 41429 1627 41463
rect 1409 41089 1443 41123
rect 5273 41089 5307 41123
rect 4997 41021 5031 41055
rect 1593 40885 1627 40919
rect 5549 40545 5583 40579
rect 1409 40477 1443 40511
rect 5273 40477 5307 40511
rect 1593 40341 1627 40375
rect 5641 40137 5675 40171
rect 1869 40069 1903 40103
rect 2053 40001 2087 40035
rect 5825 40001 5859 40035
rect 5917 39593 5951 39627
rect 1409 39389 1443 39423
rect 6101 39389 6135 39423
rect 1593 39253 1627 39287
rect 5641 39049 5675 39083
rect 3985 38981 4019 39015
rect 4169 38913 4203 38947
rect 5825 38913 5859 38947
rect 1409 38301 1443 38335
rect 6101 38301 6135 38335
rect 4261 38233 4295 38267
rect 1593 38165 1627 38199
rect 4353 38165 4387 38199
rect 5917 38165 5951 38199
rect 1409 37825 1443 37859
rect 5273 37825 5307 37859
rect 4997 37757 5031 37791
rect 1593 37621 1627 37655
rect 5273 37281 5307 37315
rect 5549 37281 5583 37315
rect 2053 37213 2087 37247
rect 1869 37077 1903 37111
rect 1409 36737 1443 36771
rect 5273 36737 5307 36771
rect 4997 36669 5031 36703
rect 1593 36601 1627 36635
rect 7205 51969 7239 52003
rect 7021 36601 7055 36635
rect 7113 50881 7147 50915
rect 6929 36465 6963 36499
rect 5549 36193 5583 36227
rect 1409 36125 1443 36159
rect 5273 36125 5307 36159
rect 1593 35989 1627 36023
rect 4353 35785 4387 35819
rect 2053 35717 2087 35751
rect 1869 35649 1903 35683
rect 4537 35649 4571 35683
rect 5273 35649 5307 35683
rect 4997 35581 5031 35615
rect 5273 35037 5307 35071
rect 5549 35037 5583 35071
rect 2513 34697 2547 34731
rect 2053 34629 2087 34663
rect 1869 34561 1903 34595
rect 2697 34561 2731 34595
rect 5273 34561 5307 34595
rect 4997 34493 5031 34527
rect 3065 34153 3099 34187
rect 3801 34085 3835 34119
rect 2053 34017 2087 34051
rect 5549 34017 5583 34051
rect 6929 34017 6963 34051
rect 3249 33949 3283 33983
rect 3985 33949 4019 33983
rect 5273 33949 5307 33983
rect 1869 33881 1903 33915
rect 6929 33881 6963 33915
rect 2053 33541 2087 33575
rect 1869 33473 1903 33507
rect 5273 33473 5307 33507
rect 4997 33405 5031 33439
rect 5549 32929 5583 32963
rect 5273 32861 5307 32895
rect 2053 32453 2087 32487
rect 1869 32385 1903 32419
rect 5273 32385 5307 32419
rect 4997 32317 5031 32351
rect 2513 31977 2547 32011
rect 5917 31977 5951 32011
rect 2053 31841 2087 31875
rect 1869 31773 1903 31807
rect 2697 31773 2731 31807
rect 6101 31773 6135 31807
rect 5641 31433 5675 31467
rect 4629 31365 4663 31399
rect 4813 31297 4847 31331
rect 5825 31297 5859 31331
rect 5273 30889 5307 30923
rect 5917 30889 5951 30923
rect 6929 30889 6963 30923
rect 1685 30753 1719 30787
rect 1409 30685 1443 30719
rect 5457 30685 5491 30719
rect 6101 30685 6135 30719
rect 2053 30277 2087 30311
rect 5549 30277 5583 30311
rect 1869 30209 1903 30243
rect 2697 30209 2731 30243
rect 5365 30209 5399 30243
rect 2513 30073 2547 30107
rect 2881 29733 2915 29767
rect 5549 29665 5583 29699
rect 1593 29597 1627 29631
rect 5273 29597 5307 29631
rect 2697 29529 2731 29563
rect 1409 29461 1443 29495
rect 1409 29257 1443 29291
rect 2881 29189 2915 29223
rect 3065 29189 3099 29223
rect 1593 29121 1627 29155
rect 2145 29121 2179 29155
rect 5273 29121 5307 29155
rect 2329 29053 2363 29087
rect 4997 29053 5031 29087
rect 1777 28713 1811 28747
rect 5181 28713 5215 28747
rect 5917 28713 5951 28747
rect 1961 28509 1995 28543
rect 6101 28509 6135 28543
rect 7113 28645 7147 28679
rect 5089 28441 5123 28475
rect 7021 28441 7055 28475
rect 7113 28373 7147 28407
rect 1593 28169 1627 28203
rect 2237 28169 2271 28203
rect 1777 28033 1811 28067
rect 2421 28033 2455 28067
rect 5825 28033 5859 28067
rect 5641 27829 5675 27863
rect 5917 27625 5951 27659
rect 6929 27625 6963 27659
rect 4445 27557 4479 27591
rect 2053 27489 2087 27523
rect 5549 27421 5583 27455
rect 5825 27421 5859 27455
rect 1869 27353 1903 27387
rect 4261 27353 4295 27387
rect 6101 27285 6135 27319
rect 1409 27081 1443 27115
rect 3249 27081 3283 27115
rect 4905 27081 4939 27115
rect 3157 27013 3191 27047
rect 5825 27013 5859 27047
rect 1593 26945 1627 26979
rect 5089 26945 5123 26979
rect 5641 26945 5675 26979
rect 1409 26537 1443 26571
rect 5273 26537 5307 26571
rect 5917 26469 5951 26503
rect 1593 26333 1627 26367
rect 5457 26333 5491 26367
rect 6101 26333 6135 26367
rect 1409 25993 1443 26027
rect 4721 25993 4755 26027
rect 5365 25925 5399 25959
rect 5549 25925 5583 25959
rect 1593 25857 1627 25891
rect 4629 25857 4663 25891
rect 5917 25449 5951 25483
rect 5365 25381 5399 25415
rect 6101 25245 6135 25279
rect 5181 25177 5215 25211
rect 5641 24905 5675 24939
rect 1593 24769 1627 24803
rect 5825 24769 5859 24803
rect 1409 24633 1443 24667
rect 1501 24361 1535 24395
rect 4353 24361 4387 24395
rect 5917 24361 5951 24395
rect 6929 24361 6963 24395
rect 7021 27285 7055 27319
rect 5273 24293 5307 24327
rect 1685 24157 1719 24191
rect 5457 24157 5491 24191
rect 6101 24157 6135 24191
rect 4261 24089 4295 24123
rect 1409 23817 1443 23851
rect 1593 23681 1627 23715
rect 5181 23681 5215 23715
rect 5641 23681 5675 23715
rect 5549 23613 5583 23647
rect 5457 23477 5491 23511
rect 5825 23477 5859 23511
rect 1409 23273 1443 23307
rect 4905 23273 4939 23307
rect 5825 23273 5859 23307
rect 3249 23205 3283 23239
rect 4445 23137 4479 23171
rect 1593 23069 1627 23103
rect 5089 23069 5123 23103
rect 5549 23069 5583 23103
rect 5733 23069 5767 23103
rect 5825 23069 5859 23103
rect 7389 50201 7423 50235
rect 7941 54213 7975 54247
rect 7757 53125 7791 53159
rect 7481 47209 7515 47243
rect 7297 38709 7331 38743
rect 7389 47005 7423 47039
rect 7297 37145 7331 37179
rect 7297 31977 7331 32011
rect 7297 31841 7331 31875
rect 7481 42245 7515 42279
rect 7573 46461 7607 46495
rect 7481 42109 7515 42143
rect 7481 41497 7515 41531
rect 7481 41383 7515 41417
rect 7573 41225 7607 41259
rect 7757 49861 7791 49895
rect 7757 46733 7791 46767
rect 7757 46597 7791 46631
rect 7757 41497 7791 41531
rect 7941 41633 7975 41667
rect 7941 41497 7975 41531
rect 7941 41361 7975 41395
rect 7665 40545 7699 40579
rect 7665 40409 7699 40443
rect 7481 38709 7515 38743
rect 7941 41225 7975 41259
rect 7757 37281 7791 37315
rect 7849 41157 7883 41191
rect 7665 36193 7699 36227
rect 7757 37145 7791 37179
rect 7573 35037 7607 35071
rect 7665 34493 7699 34527
rect 7573 33813 7607 33847
rect 7573 31841 7607 31875
rect 7481 30277 7515 30311
rect 7389 28781 7423 28815
rect 7573 30141 7607 30175
rect 7297 28713 7331 28747
rect 7205 27013 7239 27047
rect 7389 28645 7423 28679
rect 7389 25925 7423 25959
rect 7481 28441 7515 28475
rect 7757 32929 7791 32963
rect 7941 37145 7975 37179
rect 7849 29665 7883 29699
rect 7941 36601 7975 36635
rect 7665 26469 7699 26503
rect 7757 28781 7791 28815
rect 7573 25449 7607 25483
rect 7481 25381 7515 25415
rect 7113 24905 7147 24939
rect 7205 23681 7239 23715
rect 3065 23001 3099 23035
rect 4261 23001 4295 23035
rect 6929 23001 6963 23035
rect 7113 23613 7147 23647
rect 6009 22933 6043 22967
rect 7021 22933 7055 22967
rect 1409 22729 1443 22763
rect 4997 22729 5031 22763
rect 5641 22729 5675 22763
rect 1593 22593 1627 22627
rect 5181 22593 5215 22627
rect 5825 22593 5859 22627
rect 5641 22185 5675 22219
rect 6101 22185 6135 22219
rect 4721 22049 4755 22083
rect 5825 22049 5859 22083
rect 6929 22049 6963 22083
rect 1593 21981 1627 22015
rect 5917 21981 5951 22015
rect 4537 21913 4571 21947
rect 5641 21913 5675 21947
rect 1409 21845 1443 21879
rect 5641 21641 5675 21675
rect 5825 21505 5859 21539
rect 1409 21097 1443 21131
rect 5917 21097 5951 21131
rect 1593 20893 1627 20927
rect 6101 20893 6135 20927
rect 1409 20553 1443 20587
rect 5641 20553 5675 20587
rect 1593 20417 1627 20451
rect 5825 20417 5859 20451
rect 5917 20009 5951 20043
rect 2053 19941 2087 19975
rect 6101 19805 6135 19839
rect 1869 19737 1903 19771
rect 1409 19465 1443 19499
rect 5641 19465 5675 19499
rect 3341 19397 3375 19431
rect 1593 19329 1627 19363
rect 5825 19329 5859 19363
rect 3525 19193 3559 19227
rect 1409 18921 1443 18955
rect 5917 18921 5951 18955
rect 6929 18921 6963 18955
rect 1593 18717 1627 18751
rect 6101 18717 6135 18751
rect 1409 18377 1443 18411
rect 1593 18241 1627 18275
rect 5825 18241 5859 18275
rect 5641 18037 5675 18071
rect 4629 17833 4663 17867
rect 5273 17833 5307 17867
rect 5457 17629 5491 17663
rect 6101 17629 6135 17663
rect 4537 17561 4571 17595
rect 5917 17493 5951 17527
rect 6929 17493 6963 17527
rect 1409 17289 1443 17323
rect 4445 17289 4479 17323
rect 1593 17153 1627 17187
rect 4353 17153 4387 17187
rect 5825 17153 5859 17187
rect 5641 16949 5675 16983
rect 4353 16745 4387 16779
rect 5917 16745 5951 16779
rect 6929 16745 6963 16779
rect 7113 21097 7147 21131
rect 7941 27557 7975 27591
rect 7757 23205 7791 23239
rect 7389 23137 7423 23171
rect 7205 20009 7239 20043
rect 7297 21981 7331 22015
rect 7297 17833 7331 17867
rect 5733 16609 5767 16643
rect 1593 16541 1627 16575
rect 5917 16541 5951 16575
rect 4261 16473 4295 16507
rect 5641 16473 5675 16507
rect 1409 16405 1443 16439
rect 6101 16405 6135 16439
rect 4905 16201 4939 16235
rect 4813 16065 4847 16099
rect 5825 16065 5859 16099
rect 5641 15861 5675 15895
rect 1409 15657 1443 15691
rect 5273 15657 5307 15691
rect 1593 15453 1627 15487
rect 5457 15453 5491 15487
rect 6101 15453 6135 15487
rect 5917 15317 5951 15351
rect 1409 15113 1443 15147
rect 5825 15113 5859 15147
rect 1593 14977 1627 15011
rect 5365 14977 5399 15011
rect 5641 14977 5675 15011
rect 6929 14977 6963 15011
rect 5549 14909 5583 14943
rect 5641 14773 5675 14807
rect 1409 14569 1443 14603
rect 5641 14569 5675 14603
rect 6101 14501 6135 14535
rect 1593 14365 1627 14399
rect 5641 14365 5675 14399
rect 5825 14365 5859 14399
rect 5917 14365 5951 14399
rect 5641 14025 5675 14059
rect 3341 13957 3375 13991
rect 3157 13889 3191 13923
rect 5825 13889 5859 13923
rect 1409 13481 1443 13515
rect 4445 13413 4479 13447
rect 1593 13277 1627 13311
rect 6101 13277 6135 13311
rect 4261 13209 4295 13243
rect 5917 13141 5951 13175
rect 1409 12937 1443 12971
rect 5641 12937 5675 12971
rect 5181 12869 5215 12903
rect 1593 12801 1627 12835
rect 4997 12801 5031 12835
rect 5825 12801 5859 12835
rect 6101 12189 6135 12223
rect 5917 12053 5951 12087
rect 1409 11849 1443 11883
rect 5825 11849 5859 11883
rect 6929 11849 6963 11883
rect 5365 11781 5399 11815
rect 1593 11713 1627 11747
rect 5641 11713 5675 11747
rect 5549 11645 5583 11679
rect 5641 11509 5675 11543
rect 5273 11305 5307 11339
rect 5917 11305 5951 11339
rect 4629 11237 4663 11271
rect 1409 11101 1443 11135
rect 4813 11101 4847 11135
rect 5457 11101 5491 11135
rect 6101 11101 6135 11135
rect 1593 10965 1627 10999
rect 4261 10761 4295 10795
rect 5273 10761 5307 10795
rect 1409 10625 1443 10659
rect 4445 10625 4479 10659
rect 5457 10625 5491 10659
rect 1593 10421 1627 10455
rect 3801 10217 3835 10251
rect 3985 10013 4019 10047
rect 5181 10013 5215 10047
rect 5825 10013 5859 10047
rect 6929 10013 6963 10047
rect 4997 9877 5031 9911
rect 5641 9877 5675 9911
rect 1409 9537 1443 9571
rect 5457 9537 5491 9571
rect 1593 9333 1627 9367
rect 5273 9333 5307 9367
rect 2145 9129 2179 9163
rect 1409 8925 1443 8959
rect 2329 8925 2363 8959
rect 5457 8925 5491 8959
rect 6101 8925 6135 8959
rect 1593 8789 1627 8823
rect 5273 8789 5307 8823
rect 5917 8789 5951 8823
rect 6929 8789 6963 8823
rect 3617 8585 3651 8619
rect 3801 8449 3835 8483
rect 4712 8449 4746 8483
rect 4445 8381 4479 8415
rect 5825 8245 5859 8279
rect 5273 8041 5307 8075
rect 7389 15113 7423 15147
rect 7297 14773 7331 14807
rect 7205 11237 7239 11271
rect 7021 7973 7055 8007
rect 7113 8925 7147 8959
rect 6929 7905 6963 7939
rect 1409 7837 1443 7871
rect 4813 7837 4847 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 6101 7837 6135 7871
rect 1593 7701 1627 7735
rect 4629 7701 4663 7735
rect 5917 7701 5951 7735
rect 3157 7497 3191 7531
rect 4629 7497 4663 7531
rect 1409 7361 1443 7395
rect 3341 7361 3375 7395
rect 3801 7361 3835 7395
rect 4445 7361 4479 7395
rect 5089 7361 5123 7395
rect 1593 7157 1627 7191
rect 3893 7157 3927 7191
rect 5181 7157 5215 7191
rect 3801 6953 3835 6987
rect 4997 6953 5031 6987
rect 6929 6953 6963 6987
rect 7021 7837 7055 7871
rect 5825 6885 5859 6919
rect 1409 6749 1443 6783
rect 3985 6749 4019 6783
rect 4905 6681 4939 6715
rect 5549 6681 5583 6715
rect 1593 6613 1627 6647
rect 6009 6613 6043 6647
rect 6929 6613 6963 6647
rect 2881 6409 2915 6443
rect 4169 6409 4203 6443
rect 3065 6273 3099 6307
rect 3985 6273 4019 6307
rect 4629 6273 4663 6307
rect 5457 6273 5491 6307
rect 5273 6137 5307 6171
rect 4721 6069 4755 6103
rect 1409 5661 1443 5695
rect 3249 5661 3283 5695
rect 4169 5593 4203 5627
rect 1593 5525 1627 5559
rect 3065 5525 3099 5559
rect 5457 5525 5491 5559
rect 2145 5321 2179 5355
rect 3433 5321 3467 5355
rect 5825 5321 5859 5355
rect 4712 5253 4746 5287
rect 1409 5185 1443 5219
rect 2329 5185 2363 5219
rect 3617 5185 3651 5219
rect 4445 5185 4479 5219
rect 1593 4981 1627 5015
rect 4721 4777 4755 4811
rect 5917 4777 5951 4811
rect 6101 4777 6135 4811
rect 1777 4573 1811 4607
rect 2513 4573 2547 4607
rect 4261 4573 4295 4607
rect 4721 4573 4755 4607
rect 4905 4573 4939 4607
rect 5457 4573 5491 4607
rect 5549 4573 5583 4607
rect 5917 4573 5951 4607
rect 1961 4437 1995 4471
rect 2605 4437 2639 4471
rect 4077 4437 4111 4471
rect 7113 7021 7147 7055
rect 7021 5933 7055 5967
rect 7113 6885 7147 6919
rect 7113 4777 7147 4811
rect 7297 6885 7331 6919
rect 7205 4709 7239 4743
rect 1409 4097 1443 4131
rect 2145 4097 2179 4131
rect 4261 4097 4295 4131
rect 4905 4097 4939 4131
rect 5825 4097 5859 4131
rect 6929 4097 6963 4131
rect 2329 3961 2363 3995
rect 4077 3961 4111 3995
rect 1593 3893 1627 3927
rect 4721 3893 4755 3927
rect 5641 3893 5675 3927
rect 4353 3689 4387 3723
rect 4997 3689 5031 3723
rect 1409 3485 1443 3519
rect 4537 3485 4571 3519
rect 5181 3485 5215 3519
rect 5825 3485 5859 3519
rect 1593 3349 1627 3383
rect 6009 3349 6043 3383
rect 4997 3145 5031 3179
rect 5641 3145 5675 3179
rect 3617 3077 3651 3111
rect 1409 3009 1443 3043
rect 3433 3009 3467 3043
rect 5181 3009 5215 3043
rect 5825 3009 5859 3043
rect 1593 2805 1627 2839
rect 4997 2601 5031 2635
rect 5641 2533 5675 2567
rect 1409 2397 1443 2431
rect 2329 2397 2363 2431
rect 5181 2397 5215 2431
rect 5825 2397 5859 2431
rect 1593 2261 1627 2295
rect 2145 2261 2179 2295
<< metal1 >>
rect 1104 57690 6808 57712
rect 1104 57638 2880 57690
rect 2932 57638 2944 57690
rect 2996 57638 3008 57690
rect 3060 57638 3072 57690
rect 3124 57638 3136 57690
rect 3188 57638 4811 57690
rect 4863 57638 4875 57690
rect 4927 57638 4939 57690
rect 4991 57638 5003 57690
rect 5055 57638 5067 57690
rect 5119 57638 6808 57690
rect 1104 57616 6808 57638
rect 2317 57579 2375 57585
rect 2317 57545 2329 57579
rect 2363 57576 2375 57579
rect 2774 57576 2780 57588
rect 2363 57548 2780 57576
rect 2363 57545 2375 57548
rect 2317 57539 2375 57545
rect 2774 57536 2780 57548
rect 2832 57536 2838 57588
rect 3053 57579 3111 57585
rect 3053 57545 3065 57579
rect 3099 57576 3111 57579
rect 3234 57576 3240 57588
rect 3099 57548 3240 57576
rect 3099 57545 3111 57548
rect 3053 57539 3111 57545
rect 3234 57536 3240 57548
rect 3292 57536 3298 57588
rect 4246 57576 4252 57588
rect 4207 57548 4252 57576
rect 4246 57536 4252 57548
rect 4304 57536 4310 57588
rect 4985 57579 5043 57585
rect 4985 57545 4997 57579
rect 5031 57576 5043 57579
rect 5442 57576 5448 57588
rect 5031 57548 5448 57576
rect 5031 57545 5043 57548
rect 4985 57539 5043 57545
rect 5442 57536 5448 57548
rect 5500 57536 5506 57588
rect 1397 57443 1455 57449
rect 1397 57409 1409 57443
rect 1443 57409 1455 57443
rect 1397 57403 1455 57409
rect 2133 57443 2191 57449
rect 2133 57409 2145 57443
rect 2179 57409 2191 57443
rect 2133 57403 2191 57409
rect 1412 57304 1440 57403
rect 2148 57372 2176 57403
rect 2774 57400 2780 57452
rect 2832 57440 2838 57452
rect 2869 57443 2927 57449
rect 2869 57440 2881 57443
rect 2832 57412 2881 57440
rect 2832 57400 2838 57412
rect 2869 57409 2881 57412
rect 2915 57409 2927 57443
rect 2869 57403 2927 57409
rect 4065 57443 4123 57449
rect 4065 57409 4077 57443
rect 4111 57440 4123 57443
rect 4246 57440 4252 57452
rect 4111 57412 4252 57440
rect 4111 57409 4123 57412
rect 4065 57403 4123 57409
rect 4246 57400 4252 57412
rect 4304 57400 4310 57452
rect 4801 57443 4859 57449
rect 4801 57409 4813 57443
rect 4847 57409 4859 57443
rect 5534 57440 5540 57452
rect 5495 57412 5540 57440
rect 4801 57403 4859 57409
rect 3234 57372 3240 57384
rect 2148 57344 3240 57372
rect 3234 57332 3240 57344
rect 3292 57332 3298 57384
rect 3418 57332 3424 57384
rect 3476 57372 3482 57384
rect 4816 57372 4844 57403
rect 5534 57400 5540 57412
rect 5592 57400 5598 57452
rect 3476 57344 4844 57372
rect 3476 57332 3482 57344
rect 4706 57304 4712 57316
rect 1412 57276 4712 57304
rect 4706 57264 4712 57276
rect 4764 57264 4770 57316
rect 1578 57236 1584 57248
rect 1539 57208 1584 57236
rect 1578 57196 1584 57208
rect 1636 57196 1642 57248
rect 5721 57239 5779 57245
rect 5721 57205 5733 57239
rect 5767 57236 5779 57239
rect 6178 57236 6184 57248
rect 5767 57208 6184 57236
rect 5767 57205 5779 57208
rect 5721 57199 5779 57205
rect 6178 57196 6184 57208
rect 6236 57196 6242 57248
rect 1104 57146 6808 57168
rect 1104 57094 1915 57146
rect 1967 57094 1979 57146
rect 2031 57094 2043 57146
rect 2095 57094 2107 57146
rect 2159 57094 2171 57146
rect 2223 57094 3846 57146
rect 3898 57094 3910 57146
rect 3962 57094 3974 57146
rect 4026 57094 4038 57146
rect 4090 57094 4102 57146
rect 4154 57094 5776 57146
rect 5828 57094 5840 57146
rect 5892 57094 5904 57146
rect 5956 57094 5968 57146
rect 6020 57094 6032 57146
rect 6084 57094 6808 57146
rect 1104 57072 6808 57094
rect 4522 57032 4528 57044
rect 4483 57004 4528 57032
rect 4522 56992 4528 57004
rect 4580 56992 4586 57044
rect 5258 57032 5264 57044
rect 5219 57004 5264 57032
rect 5258 56992 5264 57004
rect 5316 56992 5322 57044
rect 5997 57035 6055 57041
rect 5997 57001 6009 57035
rect 6043 57032 6055 57035
rect 6270 57032 6276 57044
rect 6043 57004 6276 57032
rect 6043 57001 6055 57004
rect 5997 56995 6055 57001
rect 6270 56992 6276 57004
rect 6328 56992 6334 57044
rect 1394 56828 1400 56840
rect 1355 56800 1400 56828
rect 1394 56788 1400 56800
rect 1452 56788 1458 56840
rect 4338 56828 4344 56840
rect 4299 56800 4344 56828
rect 4338 56788 4344 56800
rect 4396 56788 4402 56840
rect 4522 56788 4528 56840
rect 4580 56828 4586 56840
rect 5077 56831 5135 56837
rect 5077 56828 5089 56831
rect 4580 56800 5089 56828
rect 4580 56788 4586 56800
rect 5077 56797 5089 56800
rect 5123 56797 5135 56831
rect 5077 56791 5135 56797
rect 5626 56788 5632 56840
rect 5684 56828 5690 56840
rect 5813 56831 5871 56837
rect 5813 56828 5825 56831
rect 5684 56800 5825 56828
rect 5684 56788 5690 56800
rect 5813 56797 5825 56800
rect 5859 56797 5871 56831
rect 5813 56791 5871 56797
rect 1578 56692 1584 56704
rect 1539 56664 1584 56692
rect 1578 56652 1584 56664
rect 1636 56652 1642 56704
rect 1104 56602 6808 56624
rect 1104 56550 2880 56602
rect 2932 56550 2944 56602
rect 2996 56550 3008 56602
rect 3060 56550 3072 56602
rect 3124 56550 3136 56602
rect 3188 56550 4811 56602
rect 4863 56550 4875 56602
rect 4927 56550 4939 56602
rect 4991 56550 5003 56602
rect 5055 56550 5067 56602
rect 5119 56550 6808 56602
rect 1104 56528 6808 56550
rect 1581 56491 1639 56497
rect 1581 56457 1593 56491
rect 1627 56488 1639 56491
rect 3326 56488 3332 56500
rect 1627 56460 3332 56488
rect 1627 56457 1639 56460
rect 1581 56451 1639 56457
rect 3326 56448 3332 56460
rect 3384 56448 3390 56500
rect 1397 56355 1455 56361
rect 1397 56321 1409 56355
rect 1443 56352 1455 56355
rect 3326 56352 3332 56364
rect 1443 56324 3332 56352
rect 1443 56321 1455 56324
rect 1397 56315 1455 56321
rect 3326 56312 3332 56324
rect 3384 56312 3390 56364
rect 5537 56355 5595 56361
rect 5537 56321 5549 56355
rect 5583 56352 5595 56355
rect 7377 56355 7435 56361
rect 7377 56352 7389 56355
rect 5583 56324 7389 56352
rect 5583 56321 5595 56324
rect 5537 56315 5595 56321
rect 7377 56321 7389 56324
rect 7423 56321 7435 56355
rect 7377 56315 7435 56321
rect 5718 56216 5724 56228
rect 5679 56188 5724 56216
rect 5718 56176 5724 56188
rect 5776 56176 5782 56228
rect 1104 56058 6808 56080
rect 1104 56006 1915 56058
rect 1967 56006 1979 56058
rect 2031 56006 2043 56058
rect 2095 56006 2107 56058
rect 2159 56006 2171 56058
rect 2223 56006 3846 56058
rect 3898 56006 3910 56058
rect 3962 56006 3974 56058
rect 4026 56006 4038 56058
rect 4090 56006 4102 56058
rect 4154 56006 5776 56058
rect 5828 56006 5840 56058
rect 5892 56006 5904 56058
rect 5956 56006 5968 56058
rect 6020 56006 6032 56058
rect 6084 56006 6808 56058
rect 1104 55984 6808 56006
rect 4246 55944 4252 55956
rect 4207 55916 4252 55944
rect 4246 55904 4252 55916
rect 4304 55904 4310 55956
rect 1397 55743 1455 55749
rect 1397 55709 1409 55743
rect 1443 55740 1455 55743
rect 1670 55740 1676 55752
rect 1443 55712 1676 55740
rect 1443 55709 1455 55712
rect 1397 55703 1455 55709
rect 1670 55700 1676 55712
rect 1728 55700 1734 55752
rect 4430 55740 4436 55752
rect 4391 55712 4436 55740
rect 4430 55700 4436 55712
rect 4488 55700 4494 55752
rect 5813 55743 5871 55749
rect 5813 55709 5825 55743
rect 5859 55740 5871 55743
rect 6917 55743 6975 55749
rect 6917 55740 6929 55743
rect 5859 55712 6929 55740
rect 5859 55709 5871 55712
rect 5813 55703 5871 55709
rect 6917 55709 6929 55712
rect 6963 55709 6975 55743
rect 6917 55703 6975 55709
rect 4062 55632 4068 55684
rect 4120 55672 4126 55684
rect 7561 55675 7619 55681
rect 7561 55672 7573 55675
rect 4120 55644 7573 55672
rect 4120 55632 4126 55644
rect 7561 55641 7573 55644
rect 7607 55641 7619 55675
rect 7561 55635 7619 55641
rect 1578 55604 1584 55616
rect 1539 55576 1584 55604
rect 1578 55564 1584 55576
rect 1636 55564 1642 55616
rect 5994 55604 6000 55616
rect 5955 55576 6000 55604
rect 5994 55564 6000 55576
rect 6052 55564 6058 55616
rect 1104 55514 6808 55536
rect 1104 55462 2880 55514
rect 2932 55462 2944 55514
rect 2996 55462 3008 55514
rect 3060 55462 3072 55514
rect 3124 55462 3136 55514
rect 3188 55462 4811 55514
rect 4863 55462 4875 55514
rect 4927 55462 4939 55514
rect 4991 55462 5003 55514
rect 5055 55462 5067 55514
rect 5119 55462 6808 55514
rect 1104 55440 6808 55462
rect 2133 55403 2191 55409
rect 2133 55369 2145 55403
rect 2179 55400 2191 55403
rect 2774 55400 2780 55412
rect 2179 55372 2780 55400
rect 2179 55369 2191 55372
rect 2133 55363 2191 55369
rect 2774 55360 2780 55372
rect 2832 55360 2838 55412
rect 2961 55403 3019 55409
rect 2961 55369 2973 55403
rect 3007 55400 3019 55403
rect 3234 55400 3240 55412
rect 3007 55372 3240 55400
rect 3007 55369 3019 55372
rect 2961 55363 3019 55369
rect 3234 55360 3240 55372
rect 3292 55360 3298 55412
rect 4065 55403 4123 55409
rect 4065 55369 4077 55403
rect 4111 55369 4123 55403
rect 4065 55363 4123 55369
rect 4709 55403 4767 55409
rect 4709 55369 4721 55403
rect 4755 55400 4767 55403
rect 5534 55400 5540 55412
rect 4755 55372 5540 55400
rect 4755 55369 4767 55372
rect 4709 55363 4767 55369
rect 4080 55332 4108 55363
rect 5534 55360 5540 55372
rect 5592 55360 5598 55412
rect 5626 55332 5632 55344
rect 4080 55304 5632 55332
rect 5626 55292 5632 55304
rect 5684 55292 5690 55344
rect 1397 55267 1455 55273
rect 1397 55233 1409 55267
rect 1443 55264 1455 55267
rect 1486 55264 1492 55276
rect 1443 55236 1492 55264
rect 1443 55233 1455 55236
rect 1397 55227 1455 55233
rect 1486 55224 1492 55236
rect 1544 55224 1550 55276
rect 2317 55267 2375 55273
rect 2317 55233 2329 55267
rect 2363 55264 2375 55267
rect 2406 55264 2412 55276
rect 2363 55236 2412 55264
rect 2363 55233 2375 55236
rect 2317 55227 2375 55233
rect 2406 55224 2412 55236
rect 2464 55224 2470 55276
rect 3145 55267 3203 55273
rect 3145 55233 3157 55267
rect 3191 55264 3203 55267
rect 4062 55264 4068 55276
rect 3191 55236 4068 55264
rect 3191 55233 3203 55236
rect 3145 55227 3203 55233
rect 4062 55224 4068 55236
rect 4120 55224 4126 55276
rect 4246 55264 4252 55276
rect 4207 55236 4252 55264
rect 4246 55224 4252 55236
rect 4304 55224 4310 55276
rect 4893 55267 4951 55273
rect 4893 55264 4905 55267
rect 4356 55236 4905 55264
rect 4246 55088 4252 55140
rect 4304 55128 4310 55140
rect 4356 55128 4384 55236
rect 4893 55233 4905 55236
rect 4939 55233 4951 55267
rect 5350 55264 5356 55276
rect 5311 55236 5356 55264
rect 4893 55227 4951 55233
rect 5350 55224 5356 55236
rect 5408 55264 5414 55276
rect 5537 55267 5595 55273
rect 5537 55264 5549 55267
rect 5408 55236 5549 55264
rect 5408 55224 5414 55236
rect 5537 55233 5549 55236
rect 5583 55233 5595 55267
rect 5537 55227 5595 55233
rect 5718 55128 5724 55140
rect 4304 55100 4384 55128
rect 5679 55100 5724 55128
rect 4304 55088 4310 55100
rect 5718 55088 5724 55100
rect 5776 55088 5782 55140
rect 1578 55060 1584 55072
rect 1539 55032 1584 55060
rect 1578 55020 1584 55032
rect 1636 55020 1642 55072
rect 1104 54970 6808 54992
rect 1104 54918 1915 54970
rect 1967 54918 1979 54970
rect 2031 54918 2043 54970
rect 2095 54918 2107 54970
rect 2159 54918 2171 54970
rect 2223 54918 3846 54970
rect 3898 54918 3910 54970
rect 3962 54918 3974 54970
rect 4026 54918 4038 54970
rect 4090 54918 4102 54970
rect 4154 54918 5776 54970
rect 5828 54918 5840 54970
rect 5892 54918 5904 54970
rect 5956 54918 5968 54970
rect 6020 54918 6032 54970
rect 6084 54918 6808 54970
rect 1104 54896 6808 54918
rect 2133 54859 2191 54865
rect 2133 54825 2145 54859
rect 2179 54856 2191 54859
rect 3418 54856 3424 54868
rect 2179 54828 3424 54856
rect 2179 54825 2191 54828
rect 2133 54819 2191 54825
rect 3418 54816 3424 54828
rect 3476 54816 3482 54868
rect 3789 54859 3847 54865
rect 3789 54825 3801 54859
rect 3835 54856 3847 54859
rect 4522 54856 4528 54868
rect 3835 54828 4528 54856
rect 3835 54825 3847 54828
rect 3789 54819 3847 54825
rect 4522 54816 4528 54828
rect 4580 54816 4586 54868
rect 1397 54655 1455 54661
rect 1397 54621 1409 54655
rect 1443 54621 1455 54655
rect 1397 54615 1455 54621
rect 1412 54584 1440 54615
rect 1762 54612 1768 54664
rect 1820 54652 1826 54664
rect 2317 54655 2375 54661
rect 2317 54652 2329 54655
rect 1820 54624 2329 54652
rect 1820 54612 1826 54624
rect 2317 54621 2329 54624
rect 2363 54621 2375 54655
rect 2317 54615 2375 54621
rect 3510 54612 3516 54664
rect 3568 54652 3574 54664
rect 3973 54655 4031 54661
rect 3973 54652 3985 54655
rect 3568 54624 3985 54652
rect 3568 54612 3574 54624
rect 3973 54621 3985 54624
rect 4019 54621 4031 54655
rect 3973 54615 4031 54621
rect 5813 54655 5871 54661
rect 5813 54621 5825 54655
rect 5859 54652 5871 54655
rect 7285 54655 7343 54661
rect 7285 54652 7297 54655
rect 5859 54624 7297 54652
rect 5859 54621 5871 54624
rect 5813 54615 5871 54621
rect 7285 54621 7297 54624
rect 7331 54621 7343 54655
rect 7285 54615 7343 54621
rect 2774 54584 2780 54596
rect 1412 54556 2780 54584
rect 2774 54544 2780 54556
rect 2832 54544 2838 54596
rect 1578 54516 1584 54528
rect 1539 54488 1584 54516
rect 1578 54476 1584 54488
rect 1636 54476 1642 54528
rect 4614 54476 4620 54528
rect 4672 54516 4678 54528
rect 5350 54516 5356 54528
rect 4672 54488 5356 54516
rect 4672 54476 4678 54488
rect 5350 54476 5356 54488
rect 5408 54476 5414 54528
rect 5994 54516 6000 54528
rect 5955 54488 6000 54516
rect 5994 54476 6000 54488
rect 6052 54476 6058 54528
rect 1104 54426 6808 54448
rect 1104 54374 2880 54426
rect 2932 54374 2944 54426
rect 2996 54374 3008 54426
rect 3060 54374 3072 54426
rect 3124 54374 3136 54426
rect 3188 54374 4811 54426
rect 4863 54374 4875 54426
rect 4927 54374 4939 54426
rect 4991 54374 5003 54426
rect 5055 54374 5067 54426
rect 5119 54374 6808 54426
rect 1104 54352 6808 54374
rect 3237 54315 3295 54321
rect 3237 54281 3249 54315
rect 3283 54312 3295 54315
rect 3326 54312 3332 54324
rect 3283 54284 3332 54312
rect 3283 54281 3295 54284
rect 3237 54275 3295 54281
rect 3326 54272 3332 54284
rect 3384 54272 3390 54324
rect 4338 54272 4344 54324
rect 4396 54312 4402 54324
rect 4893 54315 4951 54321
rect 4893 54312 4905 54315
rect 4396 54284 4905 54312
rect 4396 54272 4402 54284
rect 4893 54281 4905 54284
rect 4939 54281 4951 54315
rect 4893 54275 4951 54281
rect 7929 54247 7987 54253
rect 7929 54244 7941 54247
rect 3436 54216 7941 54244
rect 3436 54185 3464 54216
rect 7929 54213 7941 54216
rect 7975 54213 7987 54247
rect 7929 54207 7987 54213
rect 3421 54179 3479 54185
rect 3421 54145 3433 54179
rect 3467 54145 3479 54179
rect 3421 54139 3479 54145
rect 5077 54179 5135 54185
rect 5077 54145 5089 54179
rect 5123 54176 5135 54179
rect 5350 54176 5356 54188
rect 5123 54148 5356 54176
rect 5123 54145 5135 54148
rect 5077 54139 5135 54145
rect 5350 54136 5356 54148
rect 5408 54136 5414 54188
rect 5537 54179 5595 54185
rect 5537 54145 5549 54179
rect 5583 54145 5595 54179
rect 5537 54139 5595 54145
rect 4522 54068 4528 54120
rect 4580 54108 4586 54120
rect 5552 54108 5580 54139
rect 4580 54080 5580 54108
rect 4580 54068 4586 54080
rect 5718 54040 5724 54052
rect 5679 54012 5724 54040
rect 5718 54000 5724 54012
rect 5776 54000 5782 54052
rect 1104 53882 6808 53904
rect 1104 53830 1915 53882
rect 1967 53830 1979 53882
rect 2031 53830 2043 53882
rect 2095 53830 2107 53882
rect 2159 53830 2171 53882
rect 2223 53830 3846 53882
rect 3898 53830 3910 53882
rect 3962 53830 3974 53882
rect 4026 53830 4038 53882
rect 4090 53830 4102 53882
rect 4154 53830 5776 53882
rect 5828 53830 5840 53882
rect 5892 53830 5904 53882
rect 5956 53830 5968 53882
rect 6020 53830 6032 53882
rect 6084 53830 6808 53882
rect 1104 53808 6808 53830
rect 1397 53567 1455 53573
rect 1397 53533 1409 53567
rect 1443 53564 1455 53567
rect 3418 53564 3424 53576
rect 1443 53536 3424 53564
rect 1443 53533 1455 53536
rect 1397 53527 1455 53533
rect 3418 53524 3424 53536
rect 3476 53524 3482 53576
rect 5721 53567 5779 53573
rect 5721 53533 5733 53567
rect 5767 53564 5779 53567
rect 5813 53567 5871 53573
rect 5813 53564 5825 53567
rect 5767 53536 5825 53564
rect 5767 53533 5779 53536
rect 5721 53527 5779 53533
rect 5813 53533 5825 53536
rect 5859 53564 5871 53567
rect 7009 53567 7067 53573
rect 7009 53564 7021 53567
rect 5859 53536 7021 53564
rect 5859 53533 5871 53536
rect 5813 53527 5871 53533
rect 7009 53533 7021 53536
rect 7055 53533 7067 53567
rect 7009 53527 7067 53533
rect 1578 53428 1584 53440
rect 1539 53400 1584 53428
rect 1578 53388 1584 53400
rect 1636 53388 1642 53440
rect 5994 53428 6000 53440
rect 5955 53400 6000 53428
rect 5994 53388 6000 53400
rect 6052 53388 6058 53440
rect 1104 53338 6808 53360
rect 1104 53286 2880 53338
rect 2932 53286 2944 53338
rect 2996 53286 3008 53338
rect 3060 53286 3072 53338
rect 3124 53286 3136 53338
rect 3188 53286 4811 53338
rect 4863 53286 4875 53338
rect 4927 53286 4939 53338
rect 4991 53286 5003 53338
rect 5055 53286 5067 53338
rect 5119 53286 6808 53338
rect 1104 53264 6808 53286
rect 3418 53224 3424 53236
rect 3379 53196 3424 53224
rect 3418 53184 3424 53196
rect 3476 53184 3482 53236
rect 7745 53159 7803 53165
rect 7745 53156 7757 53159
rect 3620 53128 7757 53156
rect 1397 53091 1455 53097
rect 1397 53057 1409 53091
rect 1443 53088 1455 53091
rect 2866 53088 2872 53100
rect 1443 53060 2872 53088
rect 1443 53057 1455 53060
rect 1397 53051 1455 53057
rect 2866 53048 2872 53060
rect 2924 53048 2930 53100
rect 3620 53097 3648 53128
rect 7745 53125 7757 53128
rect 7791 53125 7803 53159
rect 7745 53119 7803 53125
rect 3605 53091 3663 53097
rect 3605 53057 3617 53091
rect 3651 53057 3663 53091
rect 5537 53091 5595 53097
rect 5537 53088 5549 53091
rect 3605 53051 3663 53057
rect 5368 53060 5549 53088
rect 1578 52884 1584 52896
rect 1539 52856 1584 52884
rect 1578 52844 1584 52856
rect 1636 52844 1642 52896
rect 5258 52844 5264 52896
rect 5316 52884 5322 52896
rect 5368 52893 5396 53060
rect 5537 53057 5549 53060
rect 5583 53057 5595 53091
rect 5537 53051 5595 53057
rect 5353 52887 5411 52893
rect 5353 52884 5365 52887
rect 5316 52856 5365 52884
rect 5316 52844 5322 52856
rect 5353 52853 5365 52856
rect 5399 52853 5411 52887
rect 5353 52847 5411 52853
rect 5721 52887 5779 52893
rect 5721 52853 5733 52887
rect 5767 52884 5779 52887
rect 6178 52884 6184 52896
rect 5767 52856 6184 52884
rect 5767 52853 5779 52856
rect 5721 52847 5779 52853
rect 6178 52844 6184 52856
rect 6236 52844 6242 52896
rect 1104 52794 6808 52816
rect 1104 52742 1915 52794
rect 1967 52742 1979 52794
rect 2031 52742 2043 52794
rect 2095 52742 2107 52794
rect 2159 52742 2171 52794
rect 2223 52742 3846 52794
rect 3898 52742 3910 52794
rect 3962 52742 3974 52794
rect 4026 52742 4038 52794
rect 4090 52742 4102 52794
rect 4154 52742 5776 52794
rect 5828 52742 5840 52794
rect 5892 52742 5904 52794
rect 5956 52742 5968 52794
rect 6020 52742 6032 52794
rect 6084 52742 6808 52794
rect 1104 52720 6808 52742
rect 2774 52640 2780 52692
rect 2832 52680 2838 52692
rect 3053 52683 3111 52689
rect 3053 52680 3065 52683
rect 2832 52652 3065 52680
rect 2832 52640 2838 52652
rect 3053 52649 3065 52652
rect 3099 52649 3111 52683
rect 3053 52643 3111 52649
rect 3234 52476 3240 52488
rect 3195 52448 3240 52476
rect 3234 52436 3240 52448
rect 3292 52436 3298 52488
rect 5813 52479 5871 52485
rect 5813 52445 5825 52479
rect 5859 52476 5871 52479
rect 6454 52476 6460 52488
rect 5859 52448 6460 52476
rect 5859 52445 5871 52448
rect 5813 52439 5871 52445
rect 6454 52436 6460 52448
rect 6512 52436 6518 52488
rect 5994 52340 6000 52352
rect 5955 52312 6000 52340
rect 5994 52300 6000 52312
rect 6052 52300 6058 52352
rect 1104 52250 6808 52272
rect 1104 52198 2880 52250
rect 2932 52198 2944 52250
rect 2996 52198 3008 52250
rect 3060 52198 3072 52250
rect 3124 52198 3136 52250
rect 3188 52198 4811 52250
rect 4863 52198 4875 52250
rect 4927 52198 4939 52250
rect 4991 52198 5003 52250
rect 5055 52198 5067 52250
rect 5119 52198 6808 52250
rect 1104 52176 6808 52198
rect 3513 52139 3571 52145
rect 3513 52105 3525 52139
rect 3559 52136 3571 52139
rect 6917 52139 6975 52145
rect 6917 52136 6929 52139
rect 3559 52108 6929 52136
rect 3559 52105 3571 52108
rect 3513 52099 3571 52105
rect 6917 52105 6929 52108
rect 6963 52105 6975 52139
rect 6917 52099 6975 52105
rect 1397 52003 1455 52009
rect 1397 51969 1409 52003
rect 1443 52000 1455 52003
rect 1670 52000 1676 52012
rect 1443 51972 1676 52000
rect 1443 51969 1455 51972
rect 1397 51963 1455 51969
rect 1670 51960 1676 51972
rect 1728 51960 1734 52012
rect 3694 52000 3700 52012
rect 3655 51972 3700 52000
rect 3694 51960 3700 51972
rect 3752 51960 3758 52012
rect 5537 52003 5595 52009
rect 5537 51969 5549 52003
rect 5583 52000 5595 52003
rect 7193 52003 7251 52009
rect 7193 52000 7205 52003
rect 5583 51972 7205 52000
rect 5583 51969 5595 51972
rect 5537 51963 5595 51969
rect 7193 51969 7205 51972
rect 7239 51969 7251 52003
rect 7193 51963 7251 51969
rect 1578 51864 1584 51876
rect 1539 51836 1584 51864
rect 1578 51824 1584 51836
rect 1636 51824 1642 51876
rect 5721 51799 5779 51805
rect 5721 51765 5733 51799
rect 5767 51796 5779 51799
rect 6178 51796 6184 51808
rect 5767 51768 6184 51796
rect 5767 51765 5779 51768
rect 5721 51759 5779 51765
rect 6178 51756 6184 51768
rect 6236 51756 6242 51808
rect 1104 51706 6808 51728
rect 1104 51654 1915 51706
rect 1967 51654 1979 51706
rect 2031 51654 2043 51706
rect 2095 51654 2107 51706
rect 2159 51654 2171 51706
rect 2223 51654 3846 51706
rect 3898 51654 3910 51706
rect 3962 51654 3974 51706
rect 4026 51654 4038 51706
rect 4090 51654 4102 51706
rect 4154 51654 5776 51706
rect 5828 51654 5840 51706
rect 5892 51654 5904 51706
rect 5956 51654 5968 51706
rect 6020 51654 6032 51706
rect 6084 51654 6808 51706
rect 1104 51632 6808 51654
rect 1394 51388 1400 51400
rect 1355 51360 1400 51388
rect 1394 51348 1400 51360
rect 1452 51348 1458 51400
rect 5721 51391 5779 51397
rect 5721 51357 5733 51391
rect 5767 51388 5779 51391
rect 5813 51391 5871 51397
rect 5813 51388 5825 51391
rect 5767 51360 5825 51388
rect 5767 51357 5779 51360
rect 5721 51351 5779 51357
rect 5813 51357 5825 51360
rect 5859 51388 5871 51391
rect 6917 51391 6975 51397
rect 6917 51388 6929 51391
rect 5859 51360 6929 51388
rect 5859 51357 5871 51360
rect 5813 51351 5871 51357
rect 6917 51357 6929 51360
rect 6963 51357 6975 51391
rect 6917 51351 6975 51357
rect 1578 51252 1584 51264
rect 1539 51224 1584 51252
rect 1578 51212 1584 51224
rect 1636 51212 1642 51264
rect 5994 51252 6000 51264
rect 5955 51224 6000 51252
rect 5994 51212 6000 51224
rect 6052 51212 6058 51264
rect 1104 51162 6808 51184
rect 1104 51110 2880 51162
rect 2932 51110 2944 51162
rect 2996 51110 3008 51162
rect 3060 51110 3072 51162
rect 3124 51110 3136 51162
rect 3188 51110 4811 51162
rect 4863 51110 4875 51162
rect 4927 51110 4939 51162
rect 4991 51110 5003 51162
rect 5055 51110 5067 51162
rect 5119 51110 6808 51162
rect 1104 51088 6808 51110
rect 1394 51008 1400 51060
rect 1452 51048 1458 51060
rect 2133 51051 2191 51057
rect 2133 51048 2145 51051
rect 1452 51020 2145 51048
rect 1452 51008 1458 51020
rect 2133 51017 2145 51020
rect 2179 51017 2191 51051
rect 2133 51011 2191 51017
rect 2774 51008 2780 51060
rect 2832 51048 2838 51060
rect 2832 51020 2877 51048
rect 2832 51008 2838 51020
rect 1394 50912 1400 50924
rect 1355 50884 1400 50912
rect 1394 50872 1400 50884
rect 1452 50872 1458 50924
rect 2314 50912 2320 50924
rect 2275 50884 2320 50912
rect 2314 50872 2320 50884
rect 2372 50872 2378 50924
rect 2774 50872 2780 50924
rect 2832 50912 2838 50924
rect 2961 50915 3019 50921
rect 2961 50912 2973 50915
rect 2832 50884 2973 50912
rect 2832 50872 2838 50884
rect 2961 50881 2973 50884
rect 3007 50881 3019 50915
rect 2961 50875 3019 50881
rect 5537 50915 5595 50921
rect 5537 50881 5549 50915
rect 5583 50912 5595 50915
rect 7101 50915 7159 50921
rect 7101 50912 7113 50915
rect 5583 50884 7113 50912
rect 5583 50881 5595 50884
rect 5537 50875 5595 50881
rect 7101 50881 7113 50884
rect 7147 50881 7159 50915
rect 7101 50875 7159 50881
rect 1578 50708 1584 50720
rect 1539 50680 1584 50708
rect 1578 50668 1584 50680
rect 1636 50668 1642 50720
rect 5721 50711 5779 50717
rect 5721 50677 5733 50711
rect 5767 50708 5779 50711
rect 6362 50708 6368 50720
rect 5767 50680 6368 50708
rect 5767 50677 5779 50680
rect 5721 50671 5779 50677
rect 6362 50668 6368 50680
rect 6420 50668 6426 50720
rect 1104 50618 6808 50640
rect 1104 50566 1915 50618
rect 1967 50566 1979 50618
rect 2031 50566 2043 50618
rect 2095 50566 2107 50618
rect 2159 50566 2171 50618
rect 2223 50566 3846 50618
rect 3898 50566 3910 50618
rect 3962 50566 3974 50618
rect 4026 50566 4038 50618
rect 4090 50566 4102 50618
rect 4154 50566 5776 50618
rect 5828 50566 5840 50618
rect 5892 50566 5904 50618
rect 5956 50566 5968 50618
rect 6020 50566 6032 50618
rect 6084 50566 6808 50618
rect 1104 50544 6808 50566
rect 1394 50464 1400 50516
rect 1452 50504 1458 50516
rect 1581 50507 1639 50513
rect 1581 50504 1593 50507
rect 1452 50476 1593 50504
rect 1452 50464 1458 50476
rect 1581 50473 1593 50476
rect 1627 50473 1639 50507
rect 1581 50467 1639 50473
rect 1765 50303 1823 50309
rect 1765 50269 1777 50303
rect 1811 50300 1823 50303
rect 1811 50272 2774 50300
rect 1811 50269 1823 50272
rect 1765 50263 1823 50269
rect 2746 50232 2774 50272
rect 5534 50260 5540 50312
rect 5592 50300 5598 50312
rect 5813 50303 5871 50309
rect 5813 50300 5825 50303
rect 5592 50272 5825 50300
rect 5592 50260 5598 50272
rect 5813 50269 5825 50272
rect 5859 50269 5871 50303
rect 5813 50263 5871 50269
rect 7377 50235 7435 50241
rect 7377 50232 7389 50235
rect 2746 50204 7389 50232
rect 7377 50201 7389 50204
rect 7423 50201 7435 50235
rect 7377 50195 7435 50201
rect 5994 50164 6000 50176
rect 5955 50136 6000 50164
rect 5994 50124 6000 50136
rect 6052 50124 6058 50176
rect 1104 50074 6808 50096
rect 1104 50022 2880 50074
rect 2932 50022 2944 50074
rect 2996 50022 3008 50074
rect 3060 50022 3072 50074
rect 3124 50022 3136 50074
rect 3188 50022 4811 50074
rect 4863 50022 4875 50074
rect 4927 50022 4939 50074
rect 4991 50022 5003 50074
rect 5055 50022 5067 50074
rect 5119 50022 6808 50074
rect 1104 50000 6808 50022
rect 1670 49920 1676 49972
rect 1728 49960 1734 49972
rect 2133 49963 2191 49969
rect 2133 49960 2145 49963
rect 1728 49932 2145 49960
rect 1728 49920 1734 49932
rect 2133 49929 2145 49932
rect 2179 49929 2191 49963
rect 2133 49923 2191 49929
rect 7745 49895 7803 49901
rect 7745 49892 7757 49895
rect 2746 49864 7757 49892
rect 1397 49827 1455 49833
rect 1397 49793 1409 49827
rect 1443 49793 1455 49827
rect 1397 49787 1455 49793
rect 2317 49827 2375 49833
rect 2317 49793 2329 49827
rect 2363 49824 2375 49827
rect 2746 49824 2774 49864
rect 7745 49861 7757 49864
rect 7791 49861 7803 49895
rect 7745 49855 7803 49861
rect 2363 49796 2774 49824
rect 5537 49827 5595 49833
rect 2363 49793 2375 49796
rect 2317 49787 2375 49793
rect 5537 49793 5549 49827
rect 5583 49793 5595 49827
rect 5537 49787 5595 49793
rect 1412 49756 1440 49787
rect 3418 49756 3424 49768
rect 1412 49728 3424 49756
rect 3418 49716 3424 49728
rect 3476 49716 3482 49768
rect 4706 49716 4712 49768
rect 4764 49756 4770 49768
rect 5353 49759 5411 49765
rect 5353 49756 5365 49759
rect 4764 49728 5365 49756
rect 4764 49716 4770 49728
rect 5353 49725 5365 49728
rect 5399 49756 5411 49759
rect 5552 49756 5580 49787
rect 5399 49728 5580 49756
rect 5399 49725 5411 49728
rect 5353 49719 5411 49725
rect 1578 49620 1584 49632
rect 1539 49592 1584 49620
rect 1578 49580 1584 49592
rect 1636 49580 1642 49632
rect 5721 49623 5779 49629
rect 5721 49589 5733 49623
rect 5767 49620 5779 49623
rect 6178 49620 6184 49632
rect 5767 49592 6184 49620
rect 5767 49589 5779 49592
rect 5721 49583 5779 49589
rect 6178 49580 6184 49592
rect 6236 49580 6242 49632
rect 1104 49530 6808 49552
rect 1104 49478 1915 49530
rect 1967 49478 1979 49530
rect 2031 49478 2043 49530
rect 2095 49478 2107 49530
rect 2159 49478 2171 49530
rect 2223 49478 3846 49530
rect 3898 49478 3910 49530
rect 3962 49478 3974 49530
rect 4026 49478 4038 49530
rect 4090 49478 4102 49530
rect 4154 49478 5776 49530
rect 5828 49478 5840 49530
rect 5892 49478 5904 49530
rect 5956 49478 5968 49530
rect 6020 49478 6032 49530
rect 6084 49478 6808 49530
rect 1104 49456 6808 49478
rect 1397 49215 1455 49221
rect 1397 49181 1409 49215
rect 1443 49212 1455 49215
rect 3326 49212 3332 49224
rect 1443 49184 3332 49212
rect 1443 49181 1455 49184
rect 1397 49175 1455 49181
rect 3326 49172 3332 49184
rect 3384 49172 3390 49224
rect 4338 49172 4344 49224
rect 4396 49212 4402 49224
rect 5813 49215 5871 49221
rect 5813 49212 5825 49215
rect 4396 49184 5825 49212
rect 4396 49172 4402 49184
rect 5813 49181 5825 49184
rect 5859 49181 5871 49215
rect 5813 49175 5871 49181
rect 1578 49076 1584 49088
rect 1539 49048 1584 49076
rect 1578 49036 1584 49048
rect 1636 49036 1642 49088
rect 5994 49076 6000 49088
rect 5955 49048 6000 49076
rect 5994 49036 6000 49048
rect 6052 49036 6058 49088
rect 1104 48986 6808 49008
rect 1104 48934 2880 48986
rect 2932 48934 2944 48986
rect 2996 48934 3008 48986
rect 3060 48934 3072 48986
rect 3124 48934 3136 48986
rect 3188 48934 4811 48986
rect 4863 48934 4875 48986
rect 4927 48934 4939 48986
rect 4991 48934 5003 48986
rect 5055 48934 5067 48986
rect 5119 48934 6808 48986
rect 1104 48912 6808 48934
rect 4614 48764 4620 48816
rect 4672 48804 4678 48816
rect 5350 48804 5356 48816
rect 4672 48776 5356 48804
rect 4672 48764 4678 48776
rect 5350 48764 5356 48776
rect 5408 48764 5414 48816
rect 5537 48739 5595 48745
rect 5537 48736 5549 48739
rect 5368 48708 5549 48736
rect 4614 48492 4620 48544
rect 4672 48532 4678 48544
rect 5368 48541 5396 48708
rect 5537 48705 5549 48708
rect 5583 48705 5595 48739
rect 5537 48699 5595 48705
rect 5353 48535 5411 48541
rect 5353 48532 5365 48535
rect 4672 48504 5365 48532
rect 4672 48492 4678 48504
rect 5353 48501 5365 48504
rect 5399 48501 5411 48535
rect 5353 48495 5411 48501
rect 5721 48535 5779 48541
rect 5721 48501 5733 48535
rect 5767 48532 5779 48535
rect 6178 48532 6184 48544
rect 5767 48504 6184 48532
rect 5767 48501 5779 48504
rect 5721 48495 5779 48501
rect 6178 48492 6184 48504
rect 6236 48492 6242 48544
rect 1104 48442 6808 48464
rect 1104 48390 1915 48442
rect 1967 48390 1979 48442
rect 2031 48390 2043 48442
rect 2095 48390 2107 48442
rect 2159 48390 2171 48442
rect 2223 48390 3846 48442
rect 3898 48390 3910 48442
rect 3962 48390 3974 48442
rect 4026 48390 4038 48442
rect 4090 48390 4102 48442
rect 4154 48390 5776 48442
rect 5828 48390 5840 48442
rect 5892 48390 5904 48442
rect 5956 48390 5968 48442
rect 6020 48390 6032 48442
rect 6084 48390 6808 48442
rect 1104 48368 6808 48390
rect 4798 48288 4804 48340
rect 4856 48328 4862 48340
rect 5534 48328 5540 48340
rect 4856 48300 5540 48328
rect 4856 48288 4862 48300
rect 5534 48288 5540 48300
rect 5592 48288 5598 48340
rect 3789 48263 3847 48269
rect 3789 48260 3801 48263
rect 2746 48232 3801 48260
rect 1397 48127 1455 48133
rect 1397 48093 1409 48127
rect 1443 48124 1455 48127
rect 2746 48124 2774 48232
rect 3789 48229 3801 48232
rect 3835 48229 3847 48263
rect 3789 48223 3847 48229
rect 1443 48096 2774 48124
rect 1443 48093 1455 48096
rect 1397 48087 1455 48093
rect 2866 48084 2872 48136
rect 2924 48124 2930 48136
rect 3237 48127 3295 48133
rect 3237 48124 3249 48127
rect 2924 48096 3249 48124
rect 2924 48084 2930 48096
rect 3237 48093 3249 48096
rect 3283 48093 3295 48127
rect 3237 48087 3295 48093
rect 3510 48084 3516 48136
rect 3568 48124 3574 48136
rect 3973 48127 4031 48133
rect 3973 48124 3985 48127
rect 3568 48096 3985 48124
rect 3568 48084 3574 48096
rect 3973 48093 3985 48096
rect 4019 48093 4031 48127
rect 3973 48087 4031 48093
rect 5813 48127 5871 48133
rect 5813 48093 5825 48127
rect 5859 48124 5871 48127
rect 6638 48124 6644 48136
rect 5859 48096 6644 48124
rect 5859 48093 5871 48096
rect 5813 48087 5871 48093
rect 6638 48084 6644 48096
rect 6696 48084 6702 48136
rect 1578 47988 1584 48000
rect 1539 47960 1584 47988
rect 1578 47948 1584 47960
rect 1636 47948 1642 48000
rect 3053 47991 3111 47997
rect 3053 47957 3065 47991
rect 3099 47988 3111 47991
rect 3418 47988 3424 48000
rect 3099 47960 3424 47988
rect 3099 47957 3111 47960
rect 3053 47951 3111 47957
rect 3418 47948 3424 47960
rect 3476 47948 3482 48000
rect 5994 47988 6000 48000
rect 5955 47960 6000 47988
rect 5994 47948 6000 47960
rect 6052 47948 6058 48000
rect 1104 47898 6808 47920
rect 1104 47846 2880 47898
rect 2932 47846 2944 47898
rect 2996 47846 3008 47898
rect 3060 47846 3072 47898
rect 3124 47846 3136 47898
rect 3188 47846 4811 47898
rect 4863 47846 4875 47898
rect 4927 47846 4939 47898
rect 4991 47846 5003 47898
rect 5055 47846 5067 47898
rect 5119 47846 6808 47898
rect 1104 47824 6808 47846
rect 1397 47651 1455 47657
rect 1397 47617 1409 47651
rect 1443 47648 1455 47651
rect 4338 47648 4344 47660
rect 1443 47620 4344 47648
rect 1443 47617 1455 47620
rect 1397 47611 1455 47617
rect 4338 47608 4344 47620
rect 4396 47608 4402 47660
rect 5537 47651 5595 47657
rect 5537 47617 5549 47651
rect 5583 47617 5595 47651
rect 5537 47611 5595 47617
rect 5445 47515 5503 47521
rect 5445 47481 5457 47515
rect 5491 47512 5503 47515
rect 5552 47512 5580 47611
rect 6546 47512 6552 47524
rect 5491 47484 6552 47512
rect 5491 47481 5503 47484
rect 5445 47475 5503 47481
rect 6546 47472 6552 47484
rect 6604 47472 6610 47524
rect 1578 47444 1584 47456
rect 1539 47416 1584 47444
rect 1578 47404 1584 47416
rect 1636 47404 1642 47456
rect 5721 47447 5779 47453
rect 5721 47413 5733 47447
rect 5767 47444 5779 47447
rect 6178 47444 6184 47456
rect 5767 47416 6184 47444
rect 5767 47413 5779 47416
rect 5721 47407 5779 47413
rect 6178 47404 6184 47416
rect 6236 47404 6242 47456
rect 1104 47354 6808 47376
rect 1104 47302 1915 47354
rect 1967 47302 1979 47354
rect 2031 47302 2043 47354
rect 2095 47302 2107 47354
rect 2159 47302 2171 47354
rect 2223 47302 3846 47354
rect 3898 47302 3910 47354
rect 3962 47302 3974 47354
rect 4026 47302 4038 47354
rect 4090 47302 4102 47354
rect 4154 47302 5776 47354
rect 5828 47302 5840 47354
rect 5892 47302 5904 47354
rect 5956 47302 5968 47354
rect 6020 47302 6032 47354
rect 6084 47302 6808 47354
rect 1104 47280 6808 47302
rect 3789 47243 3847 47249
rect 3789 47209 3801 47243
rect 3835 47240 3847 47243
rect 7469 47243 7527 47249
rect 7469 47240 7481 47243
rect 3835 47212 7481 47240
rect 3835 47209 3847 47212
rect 3789 47203 3847 47209
rect 7469 47209 7481 47212
rect 7515 47209 7527 47243
rect 7469 47203 7527 47209
rect 1394 47036 1400 47048
rect 1355 47008 1400 47036
rect 1394 46996 1400 47008
rect 1452 46996 1458 47048
rect 3418 46996 3424 47048
rect 3476 47036 3482 47048
rect 3973 47039 4031 47045
rect 3973 47036 3985 47039
rect 3476 47008 3985 47036
rect 3476 46996 3482 47008
rect 3973 47005 3985 47008
rect 4019 47005 4031 47039
rect 3973 46999 4031 47005
rect 5721 47039 5779 47045
rect 5721 47005 5733 47039
rect 5767 47036 5779 47039
rect 5813 47039 5871 47045
rect 5813 47036 5825 47039
rect 5767 47008 5825 47036
rect 5767 47005 5779 47008
rect 5721 46999 5779 47005
rect 5813 47005 5825 47008
rect 5859 47036 5871 47039
rect 7377 47039 7435 47045
rect 7377 47036 7389 47039
rect 5859 47008 7389 47036
rect 5859 47005 5871 47008
rect 5813 46999 5871 47005
rect 7377 47005 7389 47008
rect 7423 47005 7435 47039
rect 7377 46999 7435 47005
rect 1578 46900 1584 46912
rect 1539 46872 1584 46900
rect 1578 46860 1584 46872
rect 1636 46860 1642 46912
rect 5994 46900 6000 46912
rect 5955 46872 6000 46900
rect 5994 46860 6000 46872
rect 6052 46860 6058 46912
rect 1104 46810 6808 46832
rect 1104 46758 2880 46810
rect 2932 46758 2944 46810
rect 2996 46758 3008 46810
rect 3060 46758 3072 46810
rect 3124 46758 3136 46810
rect 3188 46758 4811 46810
rect 4863 46758 4875 46810
rect 4927 46758 4939 46810
rect 4991 46758 5003 46810
rect 5055 46758 5067 46810
rect 5119 46758 6808 46810
rect 7742 46764 7748 46776
rect 1104 46736 6808 46758
rect 7703 46736 7748 46764
rect 7742 46724 7748 46736
rect 7800 46724 7806 46776
rect 2777 46699 2835 46705
rect 2777 46665 2789 46699
rect 2823 46696 2835 46699
rect 3326 46696 3332 46708
rect 2823 46668 3332 46696
rect 2823 46665 2835 46668
rect 2777 46659 2835 46665
rect 3326 46656 3332 46668
rect 3384 46656 3390 46708
rect 4157 46699 4215 46705
rect 4157 46665 4169 46699
rect 4203 46696 4215 46699
rect 4338 46696 4344 46708
rect 4203 46668 4344 46696
rect 4203 46665 4215 46668
rect 4157 46659 4215 46665
rect 4338 46656 4344 46668
rect 4396 46656 4402 46708
rect 7745 46631 7803 46637
rect 7745 46628 7757 46631
rect 2976 46600 7757 46628
rect 2976 46569 3004 46600
rect 7745 46597 7757 46600
rect 7791 46597 7803 46631
rect 7745 46591 7803 46597
rect 2961 46563 3019 46569
rect 2961 46529 2973 46563
rect 3007 46529 3019 46563
rect 2961 46523 3019 46529
rect 4341 46563 4399 46569
rect 4341 46529 4353 46563
rect 4387 46529 4399 46563
rect 4341 46523 4399 46529
rect 5537 46563 5595 46569
rect 5537 46529 5549 46563
rect 5583 46560 5595 46563
rect 6270 46560 6276 46572
rect 5583 46532 6276 46560
rect 5583 46529 5595 46532
rect 5537 46523 5595 46529
rect 4356 46492 4384 46523
rect 6270 46520 6276 46532
rect 6328 46520 6334 46572
rect 7561 46495 7619 46501
rect 7561 46492 7573 46495
rect 4356 46464 7573 46492
rect 7561 46461 7573 46464
rect 7607 46461 7619 46495
rect 7561 46455 7619 46461
rect 5074 46316 5080 46368
rect 5132 46356 5138 46368
rect 5258 46356 5264 46368
rect 5132 46328 5264 46356
rect 5132 46316 5138 46328
rect 5258 46316 5264 46328
rect 5316 46316 5322 46368
rect 5721 46359 5779 46365
rect 5721 46325 5733 46359
rect 5767 46356 5779 46359
rect 6178 46356 6184 46368
rect 5767 46328 6184 46356
rect 5767 46325 5779 46328
rect 5721 46319 5779 46325
rect 6178 46316 6184 46328
rect 6236 46316 6242 46368
rect 1104 46266 6808 46288
rect 1104 46214 1915 46266
rect 1967 46214 1979 46266
rect 2031 46214 2043 46266
rect 2095 46214 2107 46266
rect 2159 46214 2171 46266
rect 2223 46214 3846 46266
rect 3898 46214 3910 46266
rect 3962 46214 3974 46266
rect 4026 46214 4038 46266
rect 4090 46214 4102 46266
rect 4154 46214 5776 46266
rect 5828 46214 5840 46266
rect 5892 46214 5904 46266
rect 5956 46214 5968 46266
rect 6020 46214 6032 46266
rect 6084 46214 6808 46266
rect 1104 46192 6808 46214
rect 5350 46152 5356 46164
rect 5276 46124 5356 46152
rect 4246 46044 4252 46096
rect 4304 46084 4310 46096
rect 4706 46084 4712 46096
rect 4304 46056 4712 46084
rect 4304 46044 4310 46056
rect 4706 46044 4712 46056
rect 4764 46044 4770 46096
rect 5276 46028 5304 46124
rect 5350 46112 5356 46124
rect 5408 46112 5414 46164
rect 3234 45976 3240 46028
rect 3292 45976 3298 46028
rect 5258 45976 5264 46028
rect 5316 45976 5322 46028
rect 1397 45951 1455 45957
rect 1397 45917 1409 45951
rect 1443 45948 1455 45951
rect 2682 45948 2688 45960
rect 1443 45920 2688 45948
rect 1443 45917 1455 45920
rect 1397 45911 1455 45917
rect 2682 45908 2688 45920
rect 2740 45908 2746 45960
rect 3252 45824 3280 45976
rect 5810 45948 5816 45960
rect 5771 45920 5816 45948
rect 5810 45908 5816 45920
rect 5868 45908 5874 45960
rect 5074 45840 5080 45892
rect 5132 45840 5138 45892
rect 1578 45812 1584 45824
rect 1539 45784 1584 45812
rect 1578 45772 1584 45784
rect 1636 45772 1642 45824
rect 3234 45772 3240 45824
rect 3292 45772 3298 45824
rect 5092 45812 5120 45840
rect 5350 45812 5356 45824
rect 5092 45784 5356 45812
rect 5350 45772 5356 45784
rect 5408 45772 5414 45824
rect 5994 45812 6000 45824
rect 5955 45784 6000 45812
rect 5994 45772 6000 45784
rect 6052 45772 6058 45824
rect 1104 45722 6808 45744
rect 1104 45670 2880 45722
rect 2932 45670 2944 45722
rect 2996 45670 3008 45722
rect 3060 45670 3072 45722
rect 3124 45670 3136 45722
rect 3188 45670 4811 45722
rect 4863 45670 4875 45722
rect 4927 45670 4939 45722
rect 4991 45670 5003 45722
rect 5055 45670 5067 45722
rect 5119 45670 6808 45722
rect 1104 45648 6808 45670
rect 1397 45475 1455 45481
rect 1397 45441 1409 45475
rect 1443 45472 1455 45475
rect 1486 45472 1492 45484
rect 1443 45444 1492 45472
rect 1443 45441 1455 45444
rect 1397 45435 1455 45441
rect 1486 45432 1492 45444
rect 1544 45432 1550 45484
rect 5537 45475 5595 45481
rect 5537 45472 5549 45475
rect 5368 45444 5549 45472
rect 1578 45268 1584 45280
rect 1539 45240 1584 45268
rect 1578 45228 1584 45240
rect 1636 45228 1642 45280
rect 4706 45228 4712 45280
rect 4764 45268 4770 45280
rect 5368 45277 5396 45444
rect 5537 45441 5549 45444
rect 5583 45441 5595 45475
rect 5537 45435 5595 45441
rect 5353 45271 5411 45277
rect 5353 45268 5365 45271
rect 4764 45240 5365 45268
rect 4764 45228 4770 45240
rect 5353 45237 5365 45240
rect 5399 45237 5411 45271
rect 5353 45231 5411 45237
rect 5721 45271 5779 45277
rect 5721 45237 5733 45271
rect 5767 45268 5779 45271
rect 6178 45268 6184 45280
rect 5767 45240 6184 45268
rect 5767 45237 5779 45240
rect 5721 45231 5779 45237
rect 6178 45228 6184 45240
rect 6236 45228 6242 45280
rect 1104 45178 6808 45200
rect 1104 45126 1915 45178
rect 1967 45126 1979 45178
rect 2031 45126 2043 45178
rect 2095 45126 2107 45178
rect 2159 45126 2171 45178
rect 2223 45126 3846 45178
rect 3898 45126 3910 45178
rect 3962 45126 3974 45178
rect 4026 45126 4038 45178
rect 4090 45126 4102 45178
rect 4154 45126 5776 45178
rect 5828 45126 5840 45178
rect 5892 45126 5904 45178
rect 5956 45126 5968 45178
rect 6020 45126 6032 45178
rect 6084 45126 6808 45178
rect 1104 45104 6808 45126
rect 1394 45024 1400 45076
rect 1452 45064 1458 45076
rect 2317 45067 2375 45073
rect 2317 45064 2329 45067
rect 1452 45036 2329 45064
rect 1452 45024 1458 45036
rect 2317 45033 2329 45036
rect 2363 45033 2375 45067
rect 2317 45027 2375 45033
rect 2406 44820 2412 44872
rect 2464 44860 2470 44872
rect 2501 44863 2559 44869
rect 2501 44860 2513 44863
rect 2464 44832 2513 44860
rect 2464 44820 2470 44832
rect 2501 44829 2513 44832
rect 2547 44829 2559 44863
rect 2501 44823 2559 44829
rect 5813 44863 5871 44869
rect 5813 44829 5825 44863
rect 5859 44860 5871 44863
rect 6822 44860 6828 44872
rect 5859 44832 6828 44860
rect 5859 44829 5871 44832
rect 5813 44823 5871 44829
rect 6822 44820 6828 44832
rect 6880 44820 6886 44872
rect 5994 44724 6000 44736
rect 5955 44696 6000 44724
rect 5994 44684 6000 44696
rect 6052 44684 6058 44736
rect 1104 44634 6808 44656
rect 1104 44582 2880 44634
rect 2932 44582 2944 44634
rect 2996 44582 3008 44634
rect 3060 44582 3072 44634
rect 3124 44582 3136 44634
rect 3188 44582 4811 44634
rect 4863 44582 4875 44634
rect 4927 44582 4939 44634
rect 4991 44582 5003 44634
rect 5055 44582 5067 44634
rect 5119 44582 6808 44634
rect 1104 44560 6808 44582
rect 1397 44387 1455 44393
rect 1397 44353 1409 44387
rect 1443 44384 1455 44387
rect 3142 44384 3148 44396
rect 1443 44356 3148 44384
rect 1443 44353 1455 44356
rect 1397 44347 1455 44353
rect 3142 44344 3148 44356
rect 3200 44344 3206 44396
rect 5534 44384 5540 44396
rect 5495 44356 5540 44384
rect 5534 44344 5540 44356
rect 5592 44344 5598 44396
rect 1578 44248 1584 44260
rect 1539 44220 1584 44248
rect 1578 44208 1584 44220
rect 1636 44208 1642 44260
rect 5626 44140 5632 44192
rect 5684 44180 5690 44192
rect 5721 44183 5779 44189
rect 5721 44180 5733 44183
rect 5684 44152 5733 44180
rect 5684 44140 5690 44152
rect 5721 44149 5733 44152
rect 5767 44149 5779 44183
rect 5721 44143 5779 44149
rect 1104 44090 6808 44112
rect 1104 44038 1915 44090
rect 1967 44038 1979 44090
rect 2031 44038 2043 44090
rect 2095 44038 2107 44090
rect 2159 44038 2171 44090
rect 2223 44038 3846 44090
rect 3898 44038 3910 44090
rect 3962 44038 3974 44090
rect 4026 44038 4038 44090
rect 4090 44038 4102 44090
rect 4154 44038 5776 44090
rect 5828 44038 5840 44090
rect 5892 44038 5904 44090
rect 5956 44038 5968 44090
rect 6020 44038 6032 44090
rect 6084 44038 6808 44090
rect 1104 44016 6808 44038
rect 1210 43868 1216 43920
rect 1268 43908 1274 43920
rect 2498 43908 2504 43920
rect 1268 43880 2504 43908
rect 1268 43868 1274 43880
rect 2498 43868 2504 43880
rect 2556 43868 2562 43920
rect 1397 43775 1455 43781
rect 1397 43741 1409 43775
rect 1443 43772 1455 43775
rect 2498 43772 2504 43784
rect 1443 43744 2504 43772
rect 1443 43741 1455 43744
rect 1397 43735 1455 43741
rect 2498 43732 2504 43744
rect 2556 43732 2562 43784
rect 5813 43775 5871 43781
rect 5813 43741 5825 43775
rect 5859 43772 5871 43775
rect 6270 43772 6276 43784
rect 5859 43744 6276 43772
rect 5859 43741 5871 43744
rect 5813 43735 5871 43741
rect 6270 43732 6276 43744
rect 6328 43732 6334 43784
rect 1578 43636 1584 43648
rect 1539 43608 1584 43636
rect 1578 43596 1584 43608
rect 1636 43596 1642 43648
rect 5994 43636 6000 43648
rect 5955 43608 6000 43636
rect 5994 43596 6000 43608
rect 6052 43596 6058 43648
rect 1104 43546 6808 43568
rect 1104 43494 2880 43546
rect 2932 43494 2944 43546
rect 2996 43494 3008 43546
rect 3060 43494 3072 43546
rect 3124 43494 3136 43546
rect 3188 43494 4811 43546
rect 4863 43494 4875 43546
rect 4927 43494 4939 43546
rect 4991 43494 5003 43546
rect 5055 43494 5067 43546
rect 5119 43494 6808 43546
rect 1104 43472 6808 43494
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 5537 43299 5595 43305
rect 5537 43265 5549 43299
rect 5583 43296 5595 43299
rect 6362 43296 6368 43308
rect 5583 43268 6368 43296
rect 5583 43265 5595 43268
rect 5537 43259 5595 43265
rect 6362 43256 6368 43268
rect 6420 43256 6426 43308
rect 1578 43092 1584 43104
rect 1539 43064 1584 43092
rect 1578 43052 1584 43064
rect 1636 43052 1642 43104
rect 5626 43052 5632 43104
rect 5684 43092 5690 43104
rect 5721 43095 5779 43101
rect 5721 43092 5733 43095
rect 5684 43064 5733 43092
rect 5684 43052 5690 43064
rect 5721 43061 5733 43064
rect 5767 43061 5779 43095
rect 5721 43055 5779 43061
rect 1104 43002 6808 43024
rect 1104 42950 1915 43002
rect 1967 42950 1979 43002
rect 2031 42950 2043 43002
rect 2095 42950 2107 43002
rect 2159 42950 2171 43002
rect 2223 42950 3846 43002
rect 3898 42950 3910 43002
rect 3962 42950 3974 43002
rect 4026 42950 4038 43002
rect 4090 42950 4102 43002
rect 4154 42950 5776 43002
rect 5828 42950 5840 43002
rect 5892 42950 5904 43002
rect 5956 42950 5968 43002
rect 6020 42950 6032 43002
rect 6084 42950 6808 43002
rect 1104 42928 6808 42950
rect 1104 42458 6808 42480
rect 1104 42406 2880 42458
rect 2932 42406 2944 42458
rect 2996 42406 3008 42458
rect 3060 42406 3072 42458
rect 3124 42406 3136 42458
rect 3188 42406 4811 42458
rect 4863 42406 4875 42458
rect 4927 42406 4939 42458
rect 4991 42406 5003 42458
rect 5055 42406 5067 42458
rect 5119 42406 6808 42458
rect 1104 42384 6808 42406
rect 1394 42304 1400 42356
rect 1452 42344 1458 42356
rect 2133 42347 2191 42353
rect 2133 42344 2145 42347
rect 1452 42316 2145 42344
rect 1452 42304 1458 42316
rect 2133 42313 2145 42316
rect 2179 42313 2191 42347
rect 5442 42344 5448 42356
rect 2133 42307 2191 42313
rect 5092 42316 5448 42344
rect 5092 42288 5120 42316
rect 5442 42304 5448 42316
rect 5500 42304 5506 42356
rect 5074 42236 5080 42288
rect 5132 42236 5138 42288
rect 7466 42276 7472 42288
rect 7427 42248 7472 42276
rect 7466 42236 7472 42248
rect 7524 42236 7530 42288
rect 1397 42211 1455 42217
rect 1397 42177 1409 42211
rect 1443 42177 1455 42211
rect 1397 42171 1455 42177
rect 2317 42211 2375 42217
rect 2317 42177 2329 42211
rect 2363 42208 2375 42211
rect 2363 42180 5212 42208
rect 2363 42177 2375 42180
rect 2317 42171 2375 42177
rect 1412 42004 1440 42171
rect 5184 42140 5212 42180
rect 5442 42168 5448 42220
rect 5500 42208 5506 42220
rect 5537 42211 5595 42217
rect 5537 42208 5549 42211
rect 5500 42180 5549 42208
rect 5500 42168 5506 42180
rect 5537 42177 5549 42180
rect 5583 42177 5595 42211
rect 5537 42171 5595 42177
rect 7469 42143 7527 42149
rect 7469 42140 7481 42143
rect 5184 42112 7481 42140
rect 7469 42109 7481 42112
rect 7515 42109 7527 42143
rect 7469 42103 7527 42109
rect 1578 42072 1584 42084
rect 1539 42044 1584 42072
rect 1578 42032 1584 42044
rect 1636 42032 1642 42084
rect 5718 42072 5724 42084
rect 5679 42044 5724 42072
rect 5718 42032 5724 42044
rect 5776 42032 5782 42084
rect 5442 42004 5448 42016
rect 1044 41976 1440 42004
rect 5403 41976 5448 42004
rect 1044 41800 1072 41976
rect 5442 41964 5448 41976
rect 5500 41964 5506 42016
rect 1104 41914 6808 41936
rect 1104 41862 1915 41914
rect 1967 41862 1979 41914
rect 2031 41862 2043 41914
rect 2095 41862 2107 41914
rect 2159 41862 2171 41914
rect 2223 41862 3846 41914
rect 3898 41862 3910 41914
rect 3962 41862 3974 41914
rect 4026 41862 4038 41914
rect 4090 41862 4102 41914
rect 4154 41862 5776 41914
rect 5828 41862 5840 41914
rect 5892 41862 5904 41914
rect 5956 41862 5968 41914
rect 6020 41862 6032 41914
rect 6084 41862 6808 41914
rect 1104 41840 6808 41862
rect 3053 41803 3111 41809
rect 3053 41800 3065 41803
rect 1044 41772 3065 41800
rect 3053 41769 3065 41772
rect 3099 41769 3111 41803
rect 3053 41763 3111 41769
rect 4341 41803 4399 41809
rect 4341 41769 4353 41803
rect 4387 41800 4399 41803
rect 5166 41800 5172 41812
rect 4387 41772 5172 41800
rect 4387 41769 4399 41772
rect 4341 41763 4399 41769
rect 5166 41760 5172 41772
rect 5224 41760 5230 41812
rect 4246 41624 4252 41676
rect 4304 41664 4310 41676
rect 4522 41664 4528 41676
rect 4304 41636 4528 41664
rect 4304 41624 4310 41636
rect 4522 41624 4528 41636
rect 4580 41624 4586 41676
rect 5537 41667 5595 41673
rect 5537 41633 5549 41667
rect 5583 41664 5595 41667
rect 7929 41667 7987 41673
rect 7929 41664 7941 41667
rect 5583 41636 7941 41664
rect 5583 41633 5595 41636
rect 5537 41627 5595 41633
rect 7929 41633 7941 41636
rect 7975 41633 7987 41667
rect 7929 41627 7987 41633
rect 1397 41599 1455 41605
rect 1397 41565 1409 41599
rect 1443 41596 1455 41599
rect 2222 41596 2228 41608
rect 1443 41568 2228 41596
rect 1443 41565 1455 41568
rect 1397 41559 1455 41565
rect 2222 41556 2228 41568
rect 2280 41556 2286 41608
rect 3237 41599 3295 41605
rect 3237 41565 3249 41599
rect 3283 41596 3295 41599
rect 3326 41596 3332 41608
rect 3283 41568 3332 41596
rect 3283 41565 3295 41568
rect 3237 41559 3295 41565
rect 3326 41556 3332 41568
rect 3384 41556 3390 41608
rect 5258 41596 5264 41608
rect 5219 41568 5264 41596
rect 5258 41556 5264 41568
rect 5316 41556 5322 41608
rect 1302 41488 1308 41540
rect 1360 41528 1366 41540
rect 1670 41528 1676 41540
rect 1360 41500 1676 41528
rect 1360 41488 1366 41500
rect 1670 41488 1676 41500
rect 1728 41488 1734 41540
rect 4249 41531 4307 41537
rect 4249 41497 4261 41531
rect 4295 41497 4307 41531
rect 4249 41491 4307 41497
rect 7469 41531 7527 41537
rect 7469 41497 7481 41531
rect 7515 41528 7527 41531
rect 7650 41528 7656 41540
rect 7515 41500 7656 41528
rect 7515 41497 7527 41500
rect 7469 41491 7527 41497
rect 1578 41460 1584 41472
rect 1539 41432 1584 41460
rect 1578 41420 1584 41432
rect 1636 41420 1642 41472
rect 4264 41460 4292 41491
rect 7650 41488 7656 41500
rect 7708 41488 7714 41540
rect 7745 41531 7803 41537
rect 7745 41497 7757 41531
rect 7791 41528 7803 41531
rect 7929 41531 7987 41537
rect 7929 41528 7941 41531
rect 7791 41500 7941 41528
rect 7791 41497 7803 41500
rect 7745 41491 7803 41497
rect 7929 41497 7941 41500
rect 7975 41497 7987 41531
rect 7929 41491 7987 41497
rect 5534 41460 5540 41472
rect 4264 41432 5540 41460
rect 5534 41420 5540 41432
rect 5592 41420 5598 41472
rect 7466 41414 7472 41426
rect 1104 41370 6808 41392
rect 7427 41386 7472 41414
rect 7466 41374 7472 41386
rect 7524 41374 7530 41426
rect 7926 41392 7932 41404
rect 1104 41318 2880 41370
rect 2932 41318 2944 41370
rect 2996 41318 3008 41370
rect 3060 41318 3072 41370
rect 3124 41318 3136 41370
rect 3188 41318 4811 41370
rect 4863 41318 4875 41370
rect 4927 41318 4939 41370
rect 4991 41318 5003 41370
rect 5055 41318 5067 41370
rect 5119 41318 6808 41370
rect 7887 41364 7932 41392
rect 7926 41352 7932 41364
rect 7984 41352 7990 41404
rect 1104 41296 6808 41318
rect 3234 41216 3240 41268
rect 3292 41256 3298 41268
rect 3418 41256 3424 41268
rect 3292 41228 3424 41256
rect 3292 41216 3298 41228
rect 3418 41216 3424 41228
rect 3476 41216 3482 41268
rect 7561 41259 7619 41265
rect 7561 41225 7573 41259
rect 7607 41256 7619 41259
rect 7929 41259 7987 41265
rect 7929 41256 7941 41259
rect 7607 41228 7941 41256
rect 7607 41225 7619 41228
rect 7561 41219 7619 41225
rect 7929 41225 7941 41228
rect 7975 41225 7987 41259
rect 7929 41219 7987 41225
rect 7650 41148 7656 41200
rect 7708 41188 7714 41200
rect 7837 41191 7895 41197
rect 7837 41188 7849 41191
rect 7708 41160 7849 41188
rect 7708 41148 7714 41160
rect 7837 41157 7849 41160
rect 7883 41157 7895 41191
rect 7837 41151 7895 41157
rect 1118 41080 1124 41132
rect 1176 41120 1182 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 1176 41092 1409 41120
rect 1176 41080 1182 41092
rect 1397 41089 1409 41092
rect 1443 41089 1455 41123
rect 1397 41083 1455 41089
rect 2406 41080 2412 41132
rect 2464 41080 2470 41132
rect 2590 41080 2596 41132
rect 2648 41120 2654 41132
rect 5261 41123 5319 41129
rect 5261 41120 5273 41123
rect 2648 41092 5273 41120
rect 2648 41080 2654 41092
rect 5261 41089 5273 41092
rect 5307 41089 5319 41123
rect 5261 41083 5319 41089
rect 2424 41052 2452 41080
rect 4982 41052 4988 41064
rect 2424 41024 2636 41052
rect 4943 41024 4988 41052
rect 2608 40996 2636 41024
rect 4982 41012 4988 41024
rect 5040 41012 5046 41064
rect 5166 41012 5172 41064
rect 5224 41052 5230 41064
rect 6546 41052 6552 41064
rect 5224 41024 6552 41052
rect 5224 41012 5230 41024
rect 6546 41012 6552 41024
rect 6604 41012 6610 41064
rect 2222 40944 2228 40996
rect 2280 40984 2286 40996
rect 2406 40984 2412 40996
rect 2280 40956 2412 40984
rect 2280 40944 2286 40956
rect 2406 40944 2412 40956
rect 2464 40944 2470 40996
rect 2590 40944 2596 40996
rect 2648 40944 2654 40996
rect 1578 40916 1584 40928
rect 1539 40888 1584 40916
rect 1578 40876 1584 40888
rect 1636 40876 1642 40928
rect 1104 40826 6808 40848
rect 1104 40774 1915 40826
rect 1967 40774 1979 40826
rect 2031 40774 2043 40826
rect 2095 40774 2107 40826
rect 2159 40774 2171 40826
rect 2223 40774 3846 40826
rect 3898 40774 3910 40826
rect 3962 40774 3974 40826
rect 4026 40774 4038 40826
rect 4090 40774 4102 40826
rect 4154 40774 5776 40826
rect 5828 40774 5840 40826
rect 5892 40774 5904 40826
rect 5956 40774 5968 40826
rect 6020 40774 6032 40826
rect 6084 40774 6808 40826
rect 1104 40752 6808 40774
rect 5537 40579 5595 40585
rect 5537 40545 5549 40579
rect 5583 40576 5595 40579
rect 7653 40579 7711 40585
rect 7653 40576 7665 40579
rect 5583 40548 7665 40576
rect 5583 40545 5595 40548
rect 5537 40539 5595 40545
rect 7653 40545 7665 40548
rect 7699 40545 7711 40579
rect 7653 40539 7711 40545
rect 1394 40508 1400 40520
rect 1355 40480 1400 40508
rect 1394 40468 1400 40480
rect 1452 40468 1458 40520
rect 5261 40511 5319 40517
rect 5261 40477 5273 40511
rect 5307 40508 5319 40511
rect 5718 40508 5724 40520
rect 5307 40480 5724 40508
rect 5307 40477 5319 40480
rect 5261 40471 5319 40477
rect 5718 40468 5724 40480
rect 5776 40468 5782 40520
rect 7653 40443 7711 40449
rect 7653 40409 7665 40443
rect 7699 40440 7711 40443
rect 7742 40440 7748 40452
rect 7699 40412 7748 40440
rect 7699 40409 7711 40412
rect 7653 40403 7711 40409
rect 7742 40400 7748 40412
rect 7800 40400 7806 40452
rect 1578 40372 1584 40384
rect 1539 40344 1584 40372
rect 1578 40332 1584 40344
rect 1636 40332 1642 40384
rect 1104 40282 6808 40304
rect 1104 40230 2880 40282
rect 2932 40230 2944 40282
rect 2996 40230 3008 40282
rect 3060 40230 3072 40282
rect 3124 40230 3136 40282
rect 3188 40230 4811 40282
rect 4863 40230 4875 40282
rect 4927 40230 4939 40282
rect 4991 40230 5003 40282
rect 5055 40230 5067 40282
rect 5119 40230 6808 40282
rect 1104 40208 6808 40230
rect 5534 40128 5540 40180
rect 5592 40168 5598 40180
rect 5629 40171 5687 40177
rect 5629 40168 5641 40171
rect 5592 40140 5641 40168
rect 5592 40128 5598 40140
rect 5629 40137 5641 40140
rect 5675 40137 5687 40171
rect 5629 40131 5687 40137
rect 1857 40103 1915 40109
rect 1857 40069 1869 40103
rect 1903 40100 1915 40103
rect 1903 40072 5672 40100
rect 1903 40069 1915 40072
rect 1857 40063 1915 40069
rect 1670 39992 1676 40044
rect 1728 40032 1734 40044
rect 2041 40035 2099 40041
rect 2041 40032 2053 40035
rect 1728 40004 2053 40032
rect 1728 39992 1734 40004
rect 2041 40001 2053 40004
rect 2087 40001 2099 40035
rect 2041 39995 2099 40001
rect 5644 39976 5672 40072
rect 5810 40032 5816 40044
rect 5771 40004 5816 40032
rect 5810 39992 5816 40004
rect 5868 39992 5874 40044
rect 5626 39924 5632 39976
rect 5684 39924 5690 39976
rect 1210 39856 1216 39908
rect 1268 39896 1274 39908
rect 1670 39896 1676 39908
rect 1268 39868 1676 39896
rect 1268 39856 1274 39868
rect 1670 39856 1676 39868
rect 1728 39856 1734 39908
rect 1104 39738 6808 39760
rect 1104 39686 1915 39738
rect 1967 39686 1979 39738
rect 2031 39686 2043 39738
rect 2095 39686 2107 39738
rect 2159 39686 2171 39738
rect 2223 39686 3846 39738
rect 3898 39686 3910 39738
rect 3962 39686 3974 39738
rect 4026 39686 4038 39738
rect 4090 39686 4102 39738
rect 4154 39686 5776 39738
rect 5828 39686 5840 39738
rect 5892 39686 5904 39738
rect 5956 39686 5968 39738
rect 6020 39686 6032 39738
rect 6084 39686 6808 39738
rect 1104 39664 6808 39686
rect 5626 39584 5632 39636
rect 5684 39624 5690 39636
rect 5905 39627 5963 39633
rect 5905 39624 5917 39627
rect 5684 39596 5917 39624
rect 5684 39584 5690 39596
rect 5905 39593 5917 39596
rect 5951 39593 5963 39627
rect 5905 39587 5963 39593
rect 1210 39380 1216 39432
rect 1268 39420 1274 39432
rect 1397 39423 1455 39429
rect 1397 39420 1409 39423
rect 1268 39392 1409 39420
rect 1268 39380 1274 39392
rect 1397 39389 1409 39392
rect 1443 39389 1455 39423
rect 6086 39420 6092 39432
rect 6047 39392 6092 39420
rect 1397 39383 1455 39389
rect 6086 39380 6092 39392
rect 6144 39380 6150 39432
rect 1578 39284 1584 39296
rect 1539 39256 1584 39284
rect 1578 39244 1584 39256
rect 1636 39244 1642 39296
rect 1104 39194 6808 39216
rect 1104 39142 2880 39194
rect 2932 39142 2944 39194
rect 2996 39142 3008 39194
rect 3060 39142 3072 39194
rect 3124 39142 3136 39194
rect 3188 39142 4811 39194
rect 4863 39142 4875 39194
rect 4927 39142 4939 39194
rect 4991 39142 5003 39194
rect 5055 39142 5067 39194
rect 5119 39142 6808 39194
rect 1104 39120 6808 39142
rect 5629 39083 5687 39089
rect 5629 39080 5641 39083
rect 3988 39052 5641 39080
rect 1670 38972 1676 39024
rect 1728 39012 1734 39024
rect 3988 39021 4016 39052
rect 5629 39049 5641 39052
rect 5675 39049 5687 39083
rect 5629 39043 5687 39049
rect 6178 39040 6184 39092
rect 6236 39080 6242 39092
rect 6730 39080 6736 39092
rect 6236 39052 6736 39080
rect 6236 39040 6242 39052
rect 6730 39040 6736 39052
rect 6788 39040 6794 39092
rect 3973 39015 4031 39021
rect 1728 38984 2774 39012
rect 1728 38972 1734 38984
rect 2746 38944 2774 38984
rect 3973 38981 3985 39015
rect 4019 38981 4031 39015
rect 3973 38975 4031 38981
rect 4157 38947 4215 38953
rect 4157 38944 4169 38947
rect 2746 38916 4169 38944
rect 4157 38913 4169 38916
rect 4203 38913 4215 38947
rect 4157 38907 4215 38913
rect 5813 38947 5871 38953
rect 5813 38913 5825 38947
rect 5859 38944 5871 38947
rect 6178 38944 6184 38956
rect 5859 38916 6184 38944
rect 5859 38913 5871 38916
rect 5813 38907 5871 38913
rect 6178 38904 6184 38916
rect 6236 38904 6242 38956
rect 1394 38836 1400 38888
rect 1452 38876 1458 38888
rect 1670 38876 1676 38888
rect 1452 38848 1676 38876
rect 1452 38836 1458 38848
rect 1670 38836 1676 38848
rect 1728 38836 1734 38888
rect 1394 38700 1400 38752
rect 1452 38740 1458 38752
rect 2498 38740 2504 38752
rect 1452 38712 2504 38740
rect 1452 38700 1458 38712
rect 2498 38700 2504 38712
rect 2556 38700 2562 38752
rect 7285 38743 7343 38749
rect 7285 38709 7297 38743
rect 7331 38740 7343 38743
rect 7469 38743 7527 38749
rect 7469 38740 7481 38743
rect 7331 38712 7481 38740
rect 7331 38709 7343 38712
rect 7285 38703 7343 38709
rect 7469 38709 7481 38712
rect 7515 38709 7527 38743
rect 7469 38703 7527 38709
rect 1104 38650 6808 38672
rect 1104 38598 1915 38650
rect 1967 38598 1979 38650
rect 2031 38598 2043 38650
rect 2095 38598 2107 38650
rect 2159 38598 2171 38650
rect 2223 38598 3846 38650
rect 3898 38598 3910 38650
rect 3962 38598 3974 38650
rect 4026 38598 4038 38650
rect 4090 38598 4102 38650
rect 4154 38598 5776 38650
rect 5828 38598 5840 38650
rect 5892 38598 5904 38650
rect 5956 38598 5968 38650
rect 6020 38598 6032 38650
rect 6084 38598 6808 38650
rect 1104 38576 6808 38598
rect 3050 38496 3056 38548
rect 3108 38536 3114 38548
rect 3326 38536 3332 38548
rect 3108 38508 3332 38536
rect 3108 38496 3114 38508
rect 3326 38496 3332 38508
rect 3384 38496 3390 38548
rect 3418 38496 3424 38548
rect 3476 38496 3482 38548
rect 1302 38360 1308 38412
rect 1360 38400 1366 38412
rect 3142 38400 3148 38412
rect 1360 38372 3148 38400
rect 1360 38360 1366 38372
rect 3142 38360 3148 38372
rect 3200 38360 3206 38412
rect 3436 38400 3464 38496
rect 3878 38400 3884 38412
rect 3436 38372 3884 38400
rect 3878 38360 3884 38372
rect 3936 38360 3942 38412
rect 1397 38335 1455 38341
rect 1397 38301 1409 38335
rect 1443 38332 1455 38335
rect 2590 38332 2596 38344
rect 1443 38304 2596 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 2590 38292 2596 38304
rect 2648 38292 2654 38344
rect 2958 38292 2964 38344
rect 3016 38332 3022 38344
rect 3510 38332 3516 38344
rect 3016 38304 3516 38332
rect 3016 38292 3022 38304
rect 3510 38292 3516 38304
rect 3568 38292 3574 38344
rect 6086 38332 6092 38344
rect 6047 38304 6092 38332
rect 6086 38292 6092 38304
rect 6144 38292 6150 38344
rect 3050 38224 3056 38276
rect 3108 38224 3114 38276
rect 3142 38224 3148 38276
rect 3200 38264 3206 38276
rect 4249 38267 4307 38273
rect 3200 38236 3464 38264
rect 3200 38224 3206 38236
rect 1578 38196 1584 38208
rect 1539 38168 1584 38196
rect 1578 38156 1584 38168
rect 1636 38156 1642 38208
rect 3068 38196 3096 38224
rect 3326 38196 3332 38208
rect 3068 38168 3332 38196
rect 3326 38156 3332 38168
rect 3384 38156 3390 38208
rect 3436 38196 3464 38236
rect 4249 38233 4261 38267
rect 4295 38264 4307 38267
rect 4295 38236 5948 38264
rect 4295 38233 4307 38236
rect 4249 38227 4307 38233
rect 5920 38205 5948 38236
rect 4341 38199 4399 38205
rect 4341 38196 4353 38199
rect 3436 38168 4353 38196
rect 4341 38165 4353 38168
rect 4387 38165 4399 38199
rect 4341 38159 4399 38165
rect 5905 38199 5963 38205
rect 5905 38165 5917 38199
rect 5951 38165 5963 38199
rect 5905 38159 5963 38165
rect 1104 38106 6808 38128
rect 1104 38054 2880 38106
rect 2932 38054 2944 38106
rect 2996 38054 3008 38106
rect 3060 38054 3072 38106
rect 3124 38054 3136 38106
rect 3188 38054 4811 38106
rect 4863 38054 4875 38106
rect 4927 38054 4939 38106
rect 4991 38054 5003 38106
rect 5055 38054 5067 38106
rect 5119 38054 6808 38106
rect 1104 38032 6808 38054
rect 1762 37884 1768 37936
rect 1820 37924 1826 37936
rect 2406 37924 2412 37936
rect 1820 37896 2412 37924
rect 1820 37884 1826 37896
rect 2406 37884 2412 37896
rect 2464 37884 2470 37936
rect 1397 37859 1455 37865
rect 1397 37825 1409 37859
rect 1443 37856 1455 37859
rect 2314 37856 2320 37868
rect 1443 37828 2320 37856
rect 1443 37825 1455 37828
rect 1397 37819 1455 37825
rect 2314 37816 2320 37828
rect 2372 37816 2378 37868
rect 3878 37816 3884 37868
rect 3936 37856 3942 37868
rect 5261 37859 5319 37865
rect 5261 37856 5273 37859
rect 3936 37828 5273 37856
rect 3936 37816 3942 37828
rect 5261 37825 5273 37828
rect 5307 37825 5319 37859
rect 5261 37819 5319 37825
rect 4982 37788 4988 37800
rect 4943 37760 4988 37788
rect 4982 37748 4988 37760
rect 5040 37748 5046 37800
rect 1578 37652 1584 37664
rect 1539 37624 1584 37652
rect 1578 37612 1584 37624
rect 1636 37612 1642 37664
rect 1104 37562 6808 37584
rect 1104 37510 1915 37562
rect 1967 37510 1979 37562
rect 2031 37510 2043 37562
rect 2095 37510 2107 37562
rect 2159 37510 2171 37562
rect 2223 37510 3846 37562
rect 3898 37510 3910 37562
rect 3962 37510 3974 37562
rect 4026 37510 4038 37562
rect 4090 37510 4102 37562
rect 4154 37510 5776 37562
rect 5828 37510 5840 37562
rect 5892 37510 5904 37562
rect 5956 37510 5968 37562
rect 6020 37510 6032 37562
rect 6084 37510 6808 37562
rect 1104 37488 6808 37510
rect 5258 37408 5264 37460
rect 5316 37408 5322 37460
rect 3878 37340 3884 37392
rect 3936 37380 3942 37392
rect 5276 37380 5304 37408
rect 3936 37352 5304 37380
rect 3936 37340 3942 37352
rect 5258 37312 5264 37324
rect 5219 37284 5264 37312
rect 5258 37272 5264 37284
rect 5316 37272 5322 37324
rect 5537 37315 5595 37321
rect 5537 37281 5549 37315
rect 5583 37312 5595 37315
rect 7745 37315 7803 37321
rect 7745 37312 7757 37315
rect 5583 37284 7757 37312
rect 5583 37281 5595 37284
rect 5537 37275 5595 37281
rect 7745 37281 7757 37284
rect 7791 37281 7803 37315
rect 7745 37275 7803 37281
rect 2041 37247 2099 37253
rect 2041 37213 2053 37247
rect 2087 37244 2099 37247
rect 2087 37216 2774 37244
rect 2087 37213 2099 37216
rect 2041 37207 2099 37213
rect 2746 37176 2774 37216
rect 7285 37179 7343 37185
rect 7285 37176 7297 37179
rect 2746 37148 7297 37176
rect 7285 37145 7297 37148
rect 7331 37145 7343 37179
rect 7285 37139 7343 37145
rect 7745 37179 7803 37185
rect 7745 37145 7757 37179
rect 7791 37176 7803 37179
rect 7929 37179 7987 37185
rect 7929 37176 7941 37179
rect 7791 37148 7941 37176
rect 7791 37145 7803 37148
rect 7745 37139 7803 37145
rect 7929 37145 7941 37148
rect 7975 37145 7987 37179
rect 7929 37139 7987 37145
rect 1857 37111 1915 37117
rect 1857 37077 1869 37111
rect 1903 37108 1915 37111
rect 2682 37108 2688 37120
rect 1903 37080 2688 37108
rect 1903 37077 1915 37080
rect 1857 37071 1915 37077
rect 2682 37068 2688 37080
rect 2740 37068 2746 37120
rect 1104 37018 6808 37040
rect 1104 36966 2880 37018
rect 2932 36966 2944 37018
rect 2996 36966 3008 37018
rect 3060 36966 3072 37018
rect 3124 36966 3136 37018
rect 3188 36966 4811 37018
rect 4863 36966 4875 37018
rect 4927 36966 4939 37018
rect 4991 36966 5003 37018
rect 5055 36966 5067 37018
rect 5119 36966 6808 37018
rect 1104 36944 6808 36966
rect 1486 36864 1492 36916
rect 1544 36904 1550 36916
rect 1762 36904 1768 36916
rect 1544 36876 1768 36904
rect 1544 36864 1550 36876
rect 1762 36864 1768 36876
rect 1820 36864 1826 36916
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1670 36768 1676 36780
rect 1443 36740 1676 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 1670 36728 1676 36740
rect 1728 36728 1734 36780
rect 2774 36728 2780 36780
rect 2832 36768 2838 36780
rect 5261 36771 5319 36777
rect 5261 36768 5273 36771
rect 2832 36740 5273 36768
rect 2832 36728 2838 36740
rect 5261 36737 5273 36740
rect 5307 36737 5319 36771
rect 5261 36731 5319 36737
rect 2866 36660 2872 36712
rect 2924 36700 2930 36712
rect 3878 36700 3884 36712
rect 2924 36672 3884 36700
rect 2924 36660 2930 36672
rect 3878 36660 3884 36672
rect 3936 36660 3942 36712
rect 4982 36700 4988 36712
rect 4943 36672 4988 36700
rect 4982 36660 4988 36672
rect 5040 36660 5046 36712
rect 1578 36632 1584 36644
rect 1539 36604 1584 36632
rect 1578 36592 1584 36604
rect 1636 36592 1642 36644
rect 2774 36592 2780 36644
rect 2832 36632 2838 36644
rect 3602 36632 3608 36644
rect 2832 36604 3608 36632
rect 2832 36592 2838 36604
rect 3602 36592 3608 36604
rect 3660 36592 3666 36644
rect 4614 36592 4620 36644
rect 4672 36632 4678 36644
rect 4798 36632 4804 36644
rect 4672 36604 4804 36632
rect 4672 36592 4678 36604
rect 4798 36592 4804 36604
rect 4856 36592 4862 36644
rect 7009 36635 7067 36641
rect 7009 36601 7021 36635
rect 7055 36632 7067 36635
rect 7929 36635 7987 36641
rect 7929 36632 7941 36635
rect 7055 36604 7941 36632
rect 7055 36601 7067 36604
rect 7009 36595 7067 36601
rect 7929 36601 7941 36604
rect 7975 36601 7987 36635
rect 7929 36595 7987 36601
rect 6917 36499 6975 36505
rect 1104 36474 6808 36496
rect 1104 36422 1915 36474
rect 1967 36422 1979 36474
rect 2031 36422 2043 36474
rect 2095 36422 2107 36474
rect 2159 36422 2171 36474
rect 2223 36422 3846 36474
rect 3898 36422 3910 36474
rect 3962 36422 3974 36474
rect 4026 36422 4038 36474
rect 4090 36422 4102 36474
rect 4154 36422 5776 36474
rect 5828 36422 5840 36474
rect 5892 36422 5904 36474
rect 5956 36422 5968 36474
rect 6020 36422 6032 36474
rect 6084 36422 6808 36474
rect 6917 36465 6929 36499
rect 6963 36496 6975 36499
rect 7926 36496 7932 36508
rect 6963 36468 7932 36496
rect 6963 36465 6975 36468
rect 6917 36459 6975 36465
rect 7926 36456 7932 36468
rect 7984 36456 7990 36508
rect 1104 36400 6808 36422
rect 5534 36320 5540 36372
rect 5592 36360 5598 36372
rect 6638 36360 6644 36372
rect 5592 36332 6644 36360
rect 5592 36320 5598 36332
rect 6638 36320 6644 36332
rect 6696 36320 6702 36372
rect 5537 36227 5595 36233
rect 5537 36193 5549 36227
rect 5583 36224 5595 36227
rect 7653 36227 7711 36233
rect 7653 36224 7665 36227
rect 5583 36196 7665 36224
rect 5583 36193 5595 36196
rect 5537 36187 5595 36193
rect 7653 36193 7665 36196
rect 7699 36193 7711 36227
rect 7653 36187 7711 36193
rect 1397 36159 1455 36165
rect 1397 36125 1409 36159
rect 1443 36156 1455 36159
rect 1486 36156 1492 36168
rect 1443 36128 1492 36156
rect 1443 36125 1455 36128
rect 1397 36119 1455 36125
rect 1486 36116 1492 36128
rect 1544 36116 1550 36168
rect 5258 36156 5264 36168
rect 5219 36128 5264 36156
rect 5258 36116 5264 36128
rect 5316 36116 5322 36168
rect 2038 36048 2044 36100
rect 2096 36088 2102 36100
rect 2866 36088 2872 36100
rect 2096 36060 2872 36088
rect 2096 36048 2102 36060
rect 2866 36048 2872 36060
rect 2924 36048 2930 36100
rect 1302 35980 1308 36032
rect 1360 36020 1366 36032
rect 1581 36023 1639 36029
rect 1581 36020 1593 36023
rect 1360 35992 1593 36020
rect 1360 35980 1366 35992
rect 1581 35989 1593 35992
rect 1627 35989 1639 36023
rect 1581 35983 1639 35989
rect 1104 35930 6808 35952
rect 1104 35878 2880 35930
rect 2932 35878 2944 35930
rect 2996 35878 3008 35930
rect 3060 35878 3072 35930
rect 3124 35878 3136 35930
rect 3188 35878 4811 35930
rect 4863 35878 4875 35930
rect 4927 35878 4939 35930
rect 4991 35878 5003 35930
rect 5055 35878 5067 35930
rect 5119 35878 6808 35930
rect 1104 35856 6808 35878
rect 3234 35776 3240 35828
rect 3292 35816 3298 35828
rect 4341 35819 4399 35825
rect 4341 35816 4353 35819
rect 3292 35788 4353 35816
rect 3292 35776 3298 35788
rect 4341 35785 4353 35788
rect 4387 35785 4399 35819
rect 4341 35779 4399 35785
rect 2038 35748 2044 35760
rect 1999 35720 2044 35748
rect 2038 35708 2044 35720
rect 2096 35708 2102 35760
rect 5166 35748 5172 35760
rect 4540 35720 5172 35748
rect 1394 35640 1400 35692
rect 1452 35680 1458 35692
rect 4540 35689 4568 35720
rect 5166 35708 5172 35720
rect 5224 35708 5230 35760
rect 1857 35683 1915 35689
rect 1857 35680 1869 35683
rect 1452 35652 1869 35680
rect 1452 35640 1458 35652
rect 1857 35649 1869 35652
rect 1903 35649 1915 35683
rect 1857 35643 1915 35649
rect 4525 35683 4583 35689
rect 4525 35649 4537 35683
rect 4571 35649 4583 35683
rect 5261 35683 5319 35689
rect 5261 35680 5273 35683
rect 4525 35643 4583 35649
rect 4632 35652 5273 35680
rect 2498 35572 2504 35624
rect 2556 35612 2562 35624
rect 4632 35612 4660 35652
rect 5261 35649 5273 35652
rect 5307 35649 5319 35683
rect 5261 35643 5319 35649
rect 4982 35612 4988 35624
rect 2556 35584 4660 35612
rect 4943 35584 4988 35612
rect 2556 35572 2562 35584
rect 4982 35572 4988 35584
rect 5040 35572 5046 35624
rect 1104 35386 6808 35408
rect 1104 35334 1915 35386
rect 1967 35334 1979 35386
rect 2031 35334 2043 35386
rect 2095 35334 2107 35386
rect 2159 35334 2171 35386
rect 2223 35334 3846 35386
rect 3898 35334 3910 35386
rect 3962 35334 3974 35386
rect 4026 35334 4038 35386
rect 4090 35334 4102 35386
rect 4154 35334 5776 35386
rect 5828 35334 5840 35386
rect 5892 35334 5904 35386
rect 5956 35334 5968 35386
rect 6020 35334 6032 35386
rect 6084 35334 6808 35386
rect 1104 35312 6808 35334
rect 5258 35164 5264 35216
rect 5316 35204 5322 35216
rect 5534 35204 5540 35216
rect 5316 35176 5540 35204
rect 5316 35164 5322 35176
rect 5534 35164 5540 35176
rect 5592 35164 5598 35216
rect 5258 35068 5264 35080
rect 5219 35040 5264 35068
rect 5258 35028 5264 35040
rect 5316 35028 5322 35080
rect 5537 35071 5595 35077
rect 5537 35037 5549 35071
rect 5583 35068 5595 35071
rect 7561 35071 7619 35077
rect 7561 35068 7573 35071
rect 5583 35040 7573 35068
rect 5583 35037 5595 35040
rect 5537 35031 5595 35037
rect 7561 35037 7573 35040
rect 7607 35037 7619 35071
rect 7561 35031 7619 35037
rect 1104 34842 6808 34864
rect 1104 34790 2880 34842
rect 2932 34790 2944 34842
rect 2996 34790 3008 34842
rect 3060 34790 3072 34842
rect 3124 34790 3136 34842
rect 3188 34790 4811 34842
rect 4863 34790 4875 34842
rect 4927 34790 4939 34842
rect 4991 34790 5003 34842
rect 5055 34790 5067 34842
rect 5119 34790 6808 34842
rect 1104 34768 6808 34790
rect 2501 34731 2559 34737
rect 2501 34697 2513 34731
rect 2547 34728 2559 34731
rect 2590 34728 2596 34740
rect 2547 34700 2596 34728
rect 2547 34697 2559 34700
rect 2501 34691 2559 34697
rect 2590 34688 2596 34700
rect 2648 34688 2654 34740
rect 2041 34663 2099 34669
rect 2041 34629 2053 34663
rect 2087 34660 2099 34663
rect 4338 34660 4344 34672
rect 2087 34632 4344 34660
rect 2087 34629 2099 34632
rect 2041 34623 2099 34629
rect 4338 34620 4344 34632
rect 4396 34620 4402 34672
rect 1854 34592 1860 34604
rect 1815 34564 1860 34592
rect 1854 34552 1860 34564
rect 1912 34552 1918 34604
rect 2685 34595 2743 34601
rect 2685 34561 2697 34595
rect 2731 34561 2743 34595
rect 2685 34555 2743 34561
rect 1210 34484 1216 34536
rect 1268 34524 1274 34536
rect 2590 34524 2596 34536
rect 1268 34496 2596 34524
rect 1268 34484 1274 34496
rect 2590 34484 2596 34496
rect 2648 34484 2654 34536
rect 2700 34524 2728 34555
rect 3418 34552 3424 34604
rect 3476 34592 3482 34604
rect 5261 34595 5319 34601
rect 5261 34592 5273 34595
rect 3476 34564 5273 34592
rect 3476 34552 3482 34564
rect 5261 34561 5273 34564
rect 5307 34561 5319 34595
rect 5261 34555 5319 34561
rect 4982 34524 4988 34536
rect 2700 34496 4844 34524
rect 4943 34496 4988 34524
rect 4816 34456 4844 34496
rect 4982 34484 4988 34496
rect 5040 34484 5046 34536
rect 7653 34527 7711 34533
rect 7653 34524 7665 34527
rect 5092 34496 7665 34524
rect 5092 34456 5120 34496
rect 7653 34493 7665 34496
rect 7699 34493 7711 34527
rect 7653 34487 7711 34493
rect 4816 34428 5120 34456
rect 1104 34298 6808 34320
rect 1104 34246 1915 34298
rect 1967 34246 1979 34298
rect 2031 34246 2043 34298
rect 2095 34246 2107 34298
rect 2159 34246 2171 34298
rect 2223 34246 3846 34298
rect 3898 34246 3910 34298
rect 3962 34246 3974 34298
rect 4026 34246 4038 34298
rect 4090 34246 4102 34298
rect 4154 34246 5776 34298
rect 5828 34246 5840 34298
rect 5892 34246 5904 34298
rect 5956 34246 5968 34298
rect 6020 34246 6032 34298
rect 6084 34246 6808 34298
rect 1104 34224 6808 34246
rect 2682 34144 2688 34196
rect 2740 34184 2746 34196
rect 3053 34187 3111 34193
rect 3053 34184 3065 34187
rect 2740 34156 3065 34184
rect 2740 34144 2746 34156
rect 3053 34153 3065 34156
rect 3099 34153 3111 34187
rect 3053 34147 3111 34153
rect 1394 34076 1400 34128
rect 1452 34116 1458 34128
rect 3789 34119 3847 34125
rect 3789 34116 3801 34119
rect 1452 34088 3801 34116
rect 1452 34076 1458 34088
rect 3789 34085 3801 34088
rect 3835 34085 3847 34119
rect 3789 34079 3847 34085
rect 2041 34051 2099 34057
rect 2041 34017 2053 34051
rect 2087 34048 2099 34051
rect 2774 34048 2780 34060
rect 2087 34020 2780 34048
rect 2087 34017 2099 34020
rect 2041 34011 2099 34017
rect 2774 34008 2780 34020
rect 2832 34008 2838 34060
rect 5537 34051 5595 34057
rect 5537 34017 5549 34051
rect 5583 34048 5595 34051
rect 6917 34051 6975 34057
rect 6917 34048 6929 34051
rect 5583 34020 6929 34048
rect 5583 34017 5595 34020
rect 5537 34011 5595 34017
rect 6917 34017 6929 34020
rect 6963 34017 6975 34051
rect 6917 34011 6975 34017
rect 3237 33983 3295 33989
rect 3237 33949 3249 33983
rect 3283 33949 3295 33983
rect 3237 33943 3295 33949
rect 3973 33983 4031 33989
rect 3973 33949 3985 33983
rect 4019 33949 4031 33983
rect 5258 33980 5264 33992
rect 5219 33952 5264 33980
rect 3973 33943 4031 33949
rect 1854 33912 1860 33924
rect 1815 33884 1860 33912
rect 1854 33872 1860 33884
rect 1912 33872 1918 33924
rect 3252 33844 3280 33943
rect 3988 33912 4016 33943
rect 5258 33940 5264 33952
rect 5316 33940 5322 33992
rect 6917 33915 6975 33921
rect 6917 33912 6929 33915
rect 3988 33884 6929 33912
rect 6917 33881 6929 33884
rect 6963 33881 6975 33915
rect 6917 33875 6975 33881
rect 7561 33847 7619 33853
rect 7561 33844 7573 33847
rect 3252 33816 7573 33844
rect 7561 33813 7573 33816
rect 7607 33813 7619 33847
rect 7561 33807 7619 33813
rect 1104 33754 6808 33776
rect 1104 33702 2880 33754
rect 2932 33702 2944 33754
rect 2996 33702 3008 33754
rect 3060 33702 3072 33754
rect 3124 33702 3136 33754
rect 3188 33702 4811 33754
rect 4863 33702 4875 33754
rect 4927 33702 4939 33754
rect 4991 33702 5003 33754
rect 5055 33702 5067 33754
rect 5119 33702 6808 33754
rect 1104 33680 6808 33702
rect 2682 33600 2688 33652
rect 2740 33640 2746 33652
rect 5350 33640 5356 33652
rect 2740 33612 5356 33640
rect 2740 33600 2746 33612
rect 5350 33600 5356 33612
rect 5408 33600 5414 33652
rect 2041 33575 2099 33581
rect 2041 33541 2053 33575
rect 2087 33572 2099 33575
rect 2406 33572 2412 33584
rect 2087 33544 2412 33572
rect 2087 33541 2099 33544
rect 2041 33535 2099 33541
rect 2406 33532 2412 33544
rect 2464 33532 2470 33584
rect 1394 33464 1400 33516
rect 1452 33504 1458 33516
rect 1857 33507 1915 33513
rect 1857 33504 1869 33507
rect 1452 33476 1869 33504
rect 1452 33464 1458 33476
rect 1857 33473 1869 33476
rect 1903 33473 1915 33507
rect 1857 33467 1915 33473
rect 3510 33464 3516 33516
rect 3568 33504 3574 33516
rect 5261 33507 5319 33513
rect 5261 33504 5273 33507
rect 3568 33476 5273 33504
rect 3568 33464 3574 33476
rect 5261 33473 5273 33476
rect 5307 33473 5319 33507
rect 5261 33467 5319 33473
rect 1118 33396 1124 33448
rect 1176 33436 1182 33448
rect 2406 33436 2412 33448
rect 1176 33408 2412 33436
rect 1176 33396 1182 33408
rect 2406 33396 2412 33408
rect 2464 33396 2470 33448
rect 4982 33436 4988 33448
rect 4943 33408 4988 33436
rect 4982 33396 4988 33408
rect 5040 33396 5046 33448
rect 1104 33210 6808 33232
rect 1104 33158 1915 33210
rect 1967 33158 1979 33210
rect 2031 33158 2043 33210
rect 2095 33158 2107 33210
rect 2159 33158 2171 33210
rect 2223 33158 3846 33210
rect 3898 33158 3910 33210
rect 3962 33158 3974 33210
rect 4026 33158 4038 33210
rect 4090 33158 4102 33210
rect 4154 33158 5776 33210
rect 5828 33158 5840 33210
rect 5892 33158 5904 33210
rect 5956 33158 5968 33210
rect 6020 33158 6032 33210
rect 6084 33158 6808 33210
rect 1104 33136 6808 33158
rect 5537 32963 5595 32969
rect 5537 32929 5549 32963
rect 5583 32960 5595 32963
rect 7745 32963 7803 32969
rect 7745 32960 7757 32963
rect 5583 32932 7757 32960
rect 5583 32929 5595 32932
rect 5537 32923 5595 32929
rect 7745 32929 7757 32932
rect 7791 32929 7803 32963
rect 7745 32923 7803 32929
rect 5258 32892 5264 32904
rect 5219 32864 5264 32892
rect 5258 32852 5264 32864
rect 5316 32852 5322 32904
rect 1104 32666 6808 32688
rect 1104 32614 2880 32666
rect 2932 32614 2944 32666
rect 2996 32614 3008 32666
rect 3060 32614 3072 32666
rect 3124 32614 3136 32666
rect 3188 32614 4811 32666
rect 4863 32614 4875 32666
rect 4927 32614 4939 32666
rect 4991 32614 5003 32666
rect 5055 32614 5067 32666
rect 5119 32614 6808 32666
rect 1104 32592 6808 32614
rect 2038 32484 2044 32496
rect 1999 32456 2044 32484
rect 2038 32444 2044 32456
rect 2096 32444 2102 32496
rect 1394 32376 1400 32428
rect 1452 32416 1458 32428
rect 1857 32419 1915 32425
rect 1857 32416 1869 32419
rect 1452 32388 1869 32416
rect 1452 32376 1458 32388
rect 1857 32385 1869 32388
rect 1903 32385 1915 32419
rect 1857 32379 1915 32385
rect 5261 32419 5319 32425
rect 5261 32385 5273 32419
rect 5307 32416 5319 32419
rect 5626 32416 5632 32428
rect 5307 32388 5632 32416
rect 5307 32385 5319 32388
rect 5261 32379 5319 32385
rect 5626 32376 5632 32388
rect 5684 32376 5690 32428
rect 4982 32348 4988 32360
rect 4943 32320 4988 32348
rect 4982 32308 4988 32320
rect 5040 32308 5046 32360
rect 5166 32308 5172 32360
rect 5224 32348 5230 32360
rect 5442 32348 5448 32360
rect 5224 32320 5448 32348
rect 5224 32308 5230 32320
rect 5442 32308 5448 32320
rect 5500 32308 5506 32360
rect 1104 32122 6808 32144
rect 1104 32070 1915 32122
rect 1967 32070 1979 32122
rect 2031 32070 2043 32122
rect 2095 32070 2107 32122
rect 2159 32070 2171 32122
rect 2223 32070 3846 32122
rect 3898 32070 3910 32122
rect 3962 32070 3974 32122
rect 4026 32070 4038 32122
rect 4090 32070 4102 32122
rect 4154 32070 5776 32122
rect 5828 32070 5840 32122
rect 5892 32070 5904 32122
rect 5956 32070 5968 32122
rect 6020 32070 6032 32122
rect 6084 32070 6808 32122
rect 1104 32048 6808 32070
rect 1394 31968 1400 32020
rect 1452 32008 1458 32020
rect 1762 32008 1768 32020
rect 1452 31980 1768 32008
rect 1452 31968 1458 31980
rect 1762 31968 1768 31980
rect 1820 31968 1826 32020
rect 2501 32011 2559 32017
rect 2501 31977 2513 32011
rect 2547 32008 2559 32011
rect 2590 32008 2596 32020
rect 2547 31980 2596 32008
rect 2547 31977 2559 31980
rect 2501 31971 2559 31977
rect 2590 31968 2596 31980
rect 2648 31968 2654 32020
rect 5905 32011 5963 32017
rect 5905 31977 5917 32011
rect 5951 32008 5963 32011
rect 7285 32011 7343 32017
rect 7285 32008 7297 32011
rect 5951 31980 7297 32008
rect 5951 31977 5963 31980
rect 5905 31971 5963 31977
rect 7285 31977 7297 31980
rect 7331 31977 7343 32011
rect 7285 31971 7343 31977
rect 2041 31875 2099 31881
rect 2041 31841 2053 31875
rect 2087 31872 2099 31875
rect 4338 31872 4344 31884
rect 2087 31844 4344 31872
rect 2087 31841 2099 31844
rect 2041 31835 2099 31841
rect 4338 31832 4344 31844
rect 4396 31832 4402 31884
rect 6822 31872 6828 31884
rect 4448 31844 6828 31872
rect 1854 31804 1860 31816
rect 1815 31776 1860 31804
rect 1854 31764 1860 31776
rect 1912 31764 1918 31816
rect 2685 31807 2743 31813
rect 2685 31773 2697 31807
rect 2731 31804 2743 31807
rect 3418 31804 3424 31816
rect 2731 31776 3424 31804
rect 2731 31773 2743 31776
rect 2685 31767 2743 31773
rect 3418 31764 3424 31776
rect 3476 31764 3482 31816
rect 4448 31804 4476 31844
rect 6822 31832 6828 31844
rect 6880 31832 6886 31884
rect 7285 31875 7343 31881
rect 7285 31841 7297 31875
rect 7331 31872 7343 31875
rect 7561 31875 7619 31881
rect 7561 31872 7573 31875
rect 7331 31844 7573 31872
rect 7331 31841 7343 31844
rect 7285 31835 7343 31841
rect 7561 31841 7573 31844
rect 7607 31841 7619 31875
rect 7561 31835 7619 31841
rect 4356 31792 4476 31804
rect 4338 31740 4344 31792
rect 4396 31776 4476 31792
rect 6089 31807 6147 31813
rect 4396 31740 4402 31776
rect 6089 31773 6101 31807
rect 6135 31804 6147 31807
rect 6135 31776 6169 31804
rect 6135 31773 6147 31776
rect 6089 31767 6147 31773
rect 6104 31736 6132 31767
rect 6822 31736 6828 31748
rect 6104 31708 6828 31736
rect 6822 31696 6828 31708
rect 6880 31696 6886 31748
rect 1104 31578 6808 31600
rect 1104 31526 2880 31578
rect 2932 31526 2944 31578
rect 2996 31526 3008 31578
rect 3060 31526 3072 31578
rect 3124 31526 3136 31578
rect 3188 31526 4811 31578
rect 4863 31526 4875 31578
rect 4927 31526 4939 31578
rect 4991 31526 5003 31578
rect 5055 31526 5067 31578
rect 5119 31526 6808 31578
rect 1104 31504 6808 31526
rect 5629 31467 5687 31473
rect 5629 31464 5641 31467
rect 4632 31436 5641 31464
rect 4632 31405 4660 31436
rect 5629 31433 5641 31436
rect 5675 31433 5687 31467
rect 5629 31427 5687 31433
rect 4617 31399 4675 31405
rect 4617 31365 4629 31399
rect 4663 31365 4675 31399
rect 4617 31359 4675 31365
rect 1394 31288 1400 31340
rect 1452 31328 1458 31340
rect 4801 31331 4859 31337
rect 4801 31328 4813 31331
rect 1452 31300 4813 31328
rect 1452 31288 1458 31300
rect 4801 31297 4813 31300
rect 4847 31297 4859 31331
rect 4801 31291 4859 31297
rect 5813 31331 5871 31337
rect 5813 31297 5825 31331
rect 5859 31328 5871 31331
rect 6178 31328 6184 31340
rect 5859 31300 6184 31328
rect 5859 31297 5871 31300
rect 5813 31291 5871 31297
rect 6178 31288 6184 31300
rect 6236 31288 6242 31340
rect 1104 31034 6808 31056
rect 1104 30982 1915 31034
rect 1967 30982 1979 31034
rect 2031 30982 2043 31034
rect 2095 30982 2107 31034
rect 2159 30982 2171 31034
rect 2223 30982 3846 31034
rect 3898 30982 3910 31034
rect 3962 30982 3974 31034
rect 4026 30982 4038 31034
rect 4090 30982 4102 31034
rect 4154 30982 5776 31034
rect 5828 30982 5840 31034
rect 5892 30982 5904 31034
rect 5956 30982 5968 31034
rect 6020 30982 6032 31034
rect 6084 30982 6808 31034
rect 1104 30960 6808 30982
rect 5258 30920 5264 30932
rect 5219 30892 5264 30920
rect 5258 30880 5264 30892
rect 5316 30880 5322 30932
rect 5905 30923 5963 30929
rect 5905 30889 5917 30923
rect 5951 30920 5963 30923
rect 6917 30923 6975 30929
rect 6917 30920 6929 30923
rect 5951 30892 6929 30920
rect 5951 30889 5963 30892
rect 5905 30883 5963 30889
rect 6917 30889 6929 30892
rect 6963 30889 6975 30923
rect 6917 30883 6975 30889
rect 5166 30812 5172 30864
rect 5224 30852 5230 30864
rect 5442 30852 5448 30864
rect 5224 30824 5448 30852
rect 5224 30812 5230 30824
rect 5442 30812 5448 30824
rect 5500 30812 5506 30864
rect 1673 30787 1731 30793
rect 1673 30753 1685 30787
rect 1719 30784 1731 30787
rect 2406 30784 2412 30796
rect 1719 30756 2412 30784
rect 1719 30753 1731 30756
rect 1673 30747 1731 30753
rect 2406 30744 2412 30756
rect 2464 30744 2470 30796
rect 1394 30716 1400 30728
rect 1355 30688 1400 30716
rect 1394 30676 1400 30688
rect 1452 30676 1458 30728
rect 5442 30716 5448 30728
rect 5403 30688 5448 30716
rect 5442 30676 5448 30688
rect 5500 30676 5506 30728
rect 6089 30719 6147 30725
rect 6089 30685 6101 30719
rect 6135 30716 6147 30719
rect 6178 30716 6184 30728
rect 6135 30688 6184 30716
rect 6135 30685 6147 30688
rect 6089 30679 6147 30685
rect 6178 30676 6184 30688
rect 6236 30676 6242 30728
rect 5074 30608 5080 30660
rect 5132 30648 5138 30660
rect 5534 30648 5540 30660
rect 5132 30620 5540 30648
rect 5132 30608 5138 30620
rect 5534 30608 5540 30620
rect 5592 30608 5598 30660
rect 1104 30490 6808 30512
rect 1104 30438 2880 30490
rect 2932 30438 2944 30490
rect 2996 30438 3008 30490
rect 3060 30438 3072 30490
rect 3124 30438 3136 30490
rect 3188 30438 4811 30490
rect 4863 30438 4875 30490
rect 4927 30438 4939 30490
rect 4991 30438 5003 30490
rect 5055 30438 5067 30490
rect 5119 30438 6808 30490
rect 1104 30416 6808 30438
rect 2041 30311 2099 30317
rect 2041 30277 2053 30311
rect 2087 30308 2099 30311
rect 3694 30308 3700 30320
rect 2087 30280 3700 30308
rect 2087 30277 2099 30280
rect 2041 30271 2099 30277
rect 3694 30268 3700 30280
rect 3752 30268 3758 30320
rect 5537 30311 5595 30317
rect 5537 30277 5549 30311
rect 5583 30308 5595 30311
rect 7469 30311 7527 30317
rect 7469 30308 7481 30311
rect 5583 30280 7481 30308
rect 5583 30277 5595 30280
rect 5537 30271 5595 30277
rect 7469 30277 7481 30280
rect 7515 30277 7527 30311
rect 7469 30271 7527 30277
rect 1394 30200 1400 30252
rect 1452 30240 1458 30252
rect 1857 30243 1915 30249
rect 1857 30240 1869 30243
rect 1452 30212 1869 30240
rect 1452 30200 1458 30212
rect 1857 30209 1869 30212
rect 1903 30209 1915 30243
rect 1857 30203 1915 30209
rect 2685 30243 2743 30249
rect 2685 30209 2697 30243
rect 2731 30209 2743 30243
rect 5350 30240 5356 30252
rect 5311 30212 5356 30240
rect 2685 30203 2743 30209
rect 2700 30172 2728 30203
rect 5350 30200 5356 30212
rect 5408 30200 5414 30252
rect 7561 30175 7619 30181
rect 7561 30172 7573 30175
rect 2700 30144 7573 30172
rect 7561 30141 7573 30144
rect 7607 30141 7619 30175
rect 7561 30135 7619 30141
rect 1762 30064 1768 30116
rect 1820 30104 1826 30116
rect 2501 30107 2559 30113
rect 2501 30104 2513 30107
rect 1820 30076 2513 30104
rect 1820 30064 1826 30076
rect 2501 30073 2513 30076
rect 2547 30073 2559 30107
rect 2501 30067 2559 30073
rect 1104 29946 6808 29968
rect 1104 29894 1915 29946
rect 1967 29894 1979 29946
rect 2031 29894 2043 29946
rect 2095 29894 2107 29946
rect 2159 29894 2171 29946
rect 2223 29894 3846 29946
rect 3898 29894 3910 29946
rect 3962 29894 3974 29946
rect 4026 29894 4038 29946
rect 4090 29894 4102 29946
rect 4154 29894 5776 29946
rect 5828 29894 5840 29946
rect 5892 29894 5904 29946
rect 5956 29894 5968 29946
rect 6020 29894 6032 29946
rect 6084 29894 6808 29946
rect 1104 29872 6808 29894
rect 1578 29724 1584 29776
rect 1636 29764 1642 29776
rect 1762 29764 1768 29776
rect 1636 29736 1768 29764
rect 1636 29724 1642 29736
rect 1762 29724 1768 29736
rect 1820 29724 1826 29776
rect 2866 29764 2872 29776
rect 2827 29736 2872 29764
rect 2866 29724 2872 29736
rect 2924 29724 2930 29776
rect 4154 29724 4160 29776
rect 4212 29764 4218 29776
rect 5258 29764 5264 29776
rect 4212 29736 5264 29764
rect 4212 29724 4218 29736
rect 5258 29724 5264 29736
rect 5316 29724 5322 29776
rect 5537 29699 5595 29705
rect 5537 29665 5549 29699
rect 5583 29696 5595 29699
rect 7837 29699 7895 29705
rect 7837 29696 7849 29699
rect 5583 29668 7849 29696
rect 5583 29665 5595 29668
rect 5537 29659 5595 29665
rect 7837 29665 7849 29668
rect 7883 29665 7895 29699
rect 7837 29659 7895 29665
rect 1578 29628 1584 29640
rect 1539 29600 1584 29628
rect 1578 29588 1584 29600
rect 1636 29588 1642 29640
rect 5258 29628 5264 29640
rect 5219 29600 5264 29628
rect 5258 29588 5264 29600
rect 5316 29588 5322 29640
rect 2314 29520 2320 29572
rect 2372 29560 2378 29572
rect 2685 29563 2743 29569
rect 2685 29560 2697 29563
rect 2372 29532 2697 29560
rect 2372 29520 2378 29532
rect 2685 29529 2697 29532
rect 2731 29529 2743 29563
rect 2685 29523 2743 29529
rect 1397 29495 1455 29501
rect 1397 29461 1409 29495
rect 1443 29492 1455 29495
rect 2590 29492 2596 29504
rect 1443 29464 2596 29492
rect 1443 29461 1455 29464
rect 1397 29455 1455 29461
rect 2590 29452 2596 29464
rect 2648 29452 2654 29504
rect 1104 29402 6808 29424
rect 1104 29350 2880 29402
rect 2932 29350 2944 29402
rect 2996 29350 3008 29402
rect 3060 29350 3072 29402
rect 3124 29350 3136 29402
rect 3188 29350 4811 29402
rect 4863 29350 4875 29402
rect 4927 29350 4939 29402
rect 4991 29350 5003 29402
rect 5055 29350 5067 29402
rect 5119 29350 6808 29402
rect 1104 29328 6808 29350
rect 1397 29291 1455 29297
rect 1397 29257 1409 29291
rect 1443 29288 1455 29291
rect 5350 29288 5356 29300
rect 1443 29260 5356 29288
rect 1443 29257 1455 29260
rect 1397 29251 1455 29257
rect 5350 29248 5356 29260
rect 5408 29248 5414 29300
rect 2590 29180 2596 29232
rect 2648 29220 2654 29232
rect 2869 29223 2927 29229
rect 2869 29220 2881 29223
rect 2648 29192 2881 29220
rect 2648 29180 2654 29192
rect 2869 29189 2881 29192
rect 2915 29189 2927 29223
rect 2869 29183 2927 29189
rect 3053 29223 3111 29229
rect 3053 29189 3065 29223
rect 3099 29220 3111 29223
rect 4154 29220 4160 29232
rect 3099 29192 4160 29220
rect 3099 29189 3111 29192
rect 3053 29183 3111 29189
rect 4154 29180 4160 29192
rect 4212 29180 4218 29232
rect 1394 29112 1400 29164
rect 1452 29152 1458 29164
rect 1581 29155 1639 29161
rect 1581 29152 1593 29155
rect 1452 29124 1593 29152
rect 1452 29112 1458 29124
rect 1581 29121 1593 29124
rect 1627 29121 1639 29155
rect 1581 29115 1639 29121
rect 2133 29155 2191 29161
rect 2133 29121 2145 29155
rect 2179 29152 2191 29155
rect 2406 29152 2412 29164
rect 2179 29124 2412 29152
rect 2179 29121 2191 29124
rect 2133 29115 2191 29121
rect 2406 29112 2412 29124
rect 2464 29112 2470 29164
rect 3326 29112 3332 29164
rect 3384 29152 3390 29164
rect 5261 29155 5319 29161
rect 5261 29152 5273 29155
rect 3384 29124 5273 29152
rect 3384 29112 3390 29124
rect 5261 29121 5273 29124
rect 5307 29121 5319 29155
rect 5261 29115 5319 29121
rect 2317 29087 2375 29093
rect 2317 29053 2329 29087
rect 2363 29084 2375 29087
rect 2682 29084 2688 29096
rect 2363 29056 2688 29084
rect 2363 29053 2375 29056
rect 2317 29047 2375 29053
rect 2682 29044 2688 29056
rect 2740 29044 2746 29096
rect 4982 29084 4988 29096
rect 4943 29056 4988 29084
rect 4982 29044 4988 29056
rect 5040 29044 5046 29096
rect 3418 28976 3424 29028
rect 3476 29016 3482 29028
rect 5258 29016 5264 29028
rect 3476 28988 5264 29016
rect 3476 28976 3482 28988
rect 5258 28976 5264 28988
rect 5316 28976 5322 29028
rect 1104 28858 6808 28880
rect 1104 28806 1915 28858
rect 1967 28806 1979 28858
rect 2031 28806 2043 28858
rect 2095 28806 2107 28858
rect 2159 28806 2171 28858
rect 2223 28806 3846 28858
rect 3898 28806 3910 28858
rect 3962 28806 3974 28858
rect 4026 28806 4038 28858
rect 4090 28806 4102 28858
rect 4154 28806 5776 28858
rect 5828 28806 5840 28858
rect 5892 28806 5904 28858
rect 5956 28806 5968 28858
rect 6020 28806 6032 28858
rect 6084 28806 6808 28858
rect 1104 28784 6808 28806
rect 7377 28815 7435 28821
rect 7377 28781 7389 28815
rect 7423 28812 7435 28815
rect 7745 28815 7803 28821
rect 7745 28812 7757 28815
rect 7423 28784 7757 28812
rect 7423 28781 7435 28784
rect 7377 28775 7435 28781
rect 7745 28781 7757 28784
rect 7791 28781 7803 28815
rect 7745 28775 7803 28781
rect 1762 28744 1768 28756
rect 1723 28716 1768 28744
rect 1762 28704 1768 28716
rect 1820 28704 1826 28756
rect 5166 28744 5172 28756
rect 5127 28716 5172 28744
rect 5166 28704 5172 28716
rect 5224 28704 5230 28756
rect 5905 28747 5963 28753
rect 5905 28713 5917 28747
rect 5951 28744 5963 28747
rect 7285 28747 7343 28753
rect 7285 28744 7297 28747
rect 5951 28716 7297 28744
rect 5951 28713 5963 28716
rect 5905 28707 5963 28713
rect 7285 28713 7297 28716
rect 7331 28713 7343 28747
rect 7285 28707 7343 28713
rect 7101 28679 7159 28685
rect 7101 28645 7113 28679
rect 7147 28676 7159 28679
rect 7377 28679 7435 28685
rect 7377 28676 7389 28679
rect 7147 28648 7389 28676
rect 7147 28645 7159 28648
rect 7101 28639 7159 28645
rect 7377 28645 7389 28648
rect 7423 28645 7435 28679
rect 7377 28639 7435 28645
rect 1949 28543 2007 28549
rect 1949 28509 1961 28543
rect 1995 28509 2007 28543
rect 6086 28540 6092 28552
rect 6047 28512 6092 28540
rect 1949 28503 2007 28509
rect 1964 28404 1992 28503
rect 6086 28500 6092 28512
rect 6144 28500 6150 28552
rect 2222 28432 2228 28484
rect 2280 28472 2286 28484
rect 5077 28475 5135 28481
rect 5077 28472 5089 28475
rect 2280 28444 5089 28472
rect 2280 28432 2286 28444
rect 5077 28441 5089 28444
rect 5123 28441 5135 28475
rect 5077 28435 5135 28441
rect 7009 28475 7067 28481
rect 7009 28441 7021 28475
rect 7055 28472 7067 28475
rect 7469 28475 7527 28481
rect 7469 28472 7481 28475
rect 7055 28444 7481 28472
rect 7055 28441 7067 28444
rect 7009 28435 7067 28441
rect 7469 28441 7481 28444
rect 7515 28441 7527 28475
rect 7469 28435 7527 28441
rect 7101 28407 7159 28413
rect 7101 28404 7113 28407
rect 1964 28376 7113 28404
rect 7101 28373 7113 28376
rect 7147 28373 7159 28407
rect 7101 28367 7159 28373
rect 1104 28314 6808 28336
rect 1104 28262 2880 28314
rect 2932 28262 2944 28314
rect 2996 28262 3008 28314
rect 3060 28262 3072 28314
rect 3124 28262 3136 28314
rect 3188 28262 4811 28314
rect 4863 28262 4875 28314
rect 4927 28262 4939 28314
rect 4991 28262 5003 28314
rect 5055 28262 5067 28314
rect 5119 28262 6808 28314
rect 1104 28240 6808 28262
rect 1581 28203 1639 28209
rect 1581 28169 1593 28203
rect 1627 28200 1639 28203
rect 1670 28200 1676 28212
rect 1627 28172 1676 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 1670 28160 1676 28172
rect 1728 28160 1734 28212
rect 2222 28200 2228 28212
rect 2183 28172 2228 28200
rect 2222 28160 2228 28172
rect 2280 28160 2286 28212
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28033 1823 28067
rect 1765 28027 1823 28033
rect 2409 28067 2467 28073
rect 2409 28033 2421 28067
rect 2455 28064 2467 28067
rect 2774 28064 2780 28076
rect 2455 28036 2780 28064
rect 2455 28033 2467 28036
rect 2409 28027 2467 28033
rect 1780 27996 1808 28027
rect 2774 28024 2780 28036
rect 2832 28024 2838 28076
rect 5813 28067 5871 28073
rect 5813 28033 5825 28067
rect 5859 28064 5871 28067
rect 6178 28064 6184 28076
rect 5859 28036 6184 28064
rect 5859 28033 5871 28036
rect 5813 28027 5871 28033
rect 6178 28024 6184 28036
rect 6236 28024 6242 28076
rect 5166 27996 5172 28008
rect 1780 27968 5172 27996
rect 5166 27956 5172 27968
rect 5224 27956 5230 28008
rect 5534 27820 5540 27872
rect 5592 27860 5598 27872
rect 5629 27863 5687 27869
rect 5629 27860 5641 27863
rect 5592 27832 5641 27860
rect 5592 27820 5598 27832
rect 5629 27829 5641 27832
rect 5675 27829 5687 27863
rect 5629 27823 5687 27829
rect 1104 27770 6808 27792
rect 1104 27718 1915 27770
rect 1967 27718 1979 27770
rect 2031 27718 2043 27770
rect 2095 27718 2107 27770
rect 2159 27718 2171 27770
rect 2223 27718 3846 27770
rect 3898 27718 3910 27770
rect 3962 27718 3974 27770
rect 4026 27718 4038 27770
rect 4090 27718 4102 27770
rect 4154 27718 5776 27770
rect 5828 27718 5840 27770
rect 5892 27718 5904 27770
rect 5956 27718 5968 27770
rect 6020 27718 6032 27770
rect 6084 27718 6808 27770
rect 1104 27696 6808 27718
rect 5905 27659 5963 27665
rect 5905 27625 5917 27659
rect 5951 27656 5963 27659
rect 6917 27659 6975 27665
rect 6917 27656 6929 27659
rect 5951 27628 6929 27656
rect 5951 27625 5963 27628
rect 5905 27619 5963 27625
rect 6917 27625 6929 27628
rect 6963 27625 6975 27659
rect 6917 27619 6975 27625
rect 4433 27591 4491 27597
rect 4433 27557 4445 27591
rect 4479 27588 4491 27591
rect 7929 27591 7987 27597
rect 7929 27588 7941 27591
rect 4479 27560 7941 27588
rect 4479 27557 4491 27560
rect 4433 27551 4491 27557
rect 7929 27557 7941 27560
rect 7975 27557 7987 27591
rect 7929 27551 7987 27557
rect 2041 27523 2099 27529
rect 2041 27489 2053 27523
rect 2087 27520 2099 27523
rect 6454 27520 6460 27532
rect 2087 27492 6460 27520
rect 2087 27489 2099 27492
rect 2041 27483 2099 27489
rect 6454 27480 6460 27492
rect 6512 27480 6518 27532
rect 5537 27455 5595 27461
rect 5537 27421 5549 27455
rect 5583 27452 5595 27455
rect 5626 27452 5632 27464
rect 5583 27424 5632 27452
rect 5583 27421 5595 27424
rect 5537 27415 5595 27421
rect 5626 27412 5632 27424
rect 5684 27412 5690 27464
rect 5810 27452 5816 27464
rect 5771 27424 5816 27452
rect 5810 27412 5816 27424
rect 5868 27412 5874 27464
rect 1670 27344 1676 27396
rect 1728 27384 1734 27396
rect 1857 27387 1915 27393
rect 1857 27384 1869 27387
rect 1728 27356 1869 27384
rect 1728 27344 1734 27356
rect 1857 27353 1869 27356
rect 1903 27353 1915 27387
rect 1857 27347 1915 27353
rect 2038 27344 2044 27396
rect 2096 27384 2102 27396
rect 4249 27387 4307 27393
rect 4249 27384 4261 27387
rect 2096 27356 4261 27384
rect 2096 27344 2102 27356
rect 4249 27353 4261 27356
rect 4295 27353 4307 27387
rect 4249 27347 4307 27353
rect 6089 27319 6147 27325
rect 6089 27285 6101 27319
rect 6135 27316 6147 27319
rect 7009 27319 7067 27325
rect 7009 27316 7021 27319
rect 6135 27288 7021 27316
rect 6135 27285 6147 27288
rect 6089 27279 6147 27285
rect 7009 27285 7021 27288
rect 7055 27285 7067 27319
rect 7009 27279 7067 27285
rect 1104 27226 6808 27248
rect 1104 27174 2880 27226
rect 2932 27174 2944 27226
rect 2996 27174 3008 27226
rect 3060 27174 3072 27226
rect 3124 27174 3136 27226
rect 3188 27174 4811 27226
rect 4863 27174 4875 27226
rect 4927 27174 4939 27226
rect 4991 27174 5003 27226
rect 5055 27174 5067 27226
rect 5119 27174 6808 27226
rect 1104 27152 6808 27174
rect 1397 27115 1455 27121
rect 1397 27081 1409 27115
rect 1443 27112 1455 27115
rect 2038 27112 2044 27124
rect 1443 27084 2044 27112
rect 1443 27081 1455 27084
rect 1397 27075 1455 27081
rect 2038 27072 2044 27084
rect 2096 27072 2102 27124
rect 2498 27072 2504 27124
rect 2556 27112 2562 27124
rect 3237 27115 3295 27121
rect 3237 27112 3249 27115
rect 2556 27084 3249 27112
rect 2556 27072 2562 27084
rect 3237 27081 3249 27084
rect 3283 27081 3295 27115
rect 3237 27075 3295 27081
rect 4893 27115 4951 27121
rect 4893 27081 4905 27115
rect 4939 27112 4951 27115
rect 5166 27112 5172 27124
rect 4939 27084 5172 27112
rect 4939 27081 4951 27084
rect 4893 27075 4951 27081
rect 5166 27072 5172 27084
rect 5224 27072 5230 27124
rect 3145 27047 3203 27053
rect 3145 27013 3157 27047
rect 3191 27044 3203 27047
rect 5534 27044 5540 27056
rect 3191 27016 5540 27044
rect 3191 27013 3203 27016
rect 3145 27007 3203 27013
rect 5534 27004 5540 27016
rect 5592 27004 5598 27056
rect 5813 27047 5871 27053
rect 5813 27013 5825 27047
rect 5859 27044 5871 27047
rect 7193 27047 7251 27053
rect 7193 27044 7205 27047
rect 5859 27016 7205 27044
rect 5859 27013 5871 27016
rect 5813 27007 5871 27013
rect 7193 27013 7205 27016
rect 7239 27013 7251 27047
rect 7193 27007 7251 27013
rect 1578 26976 1584 26988
rect 1539 26948 1584 26976
rect 1578 26936 1584 26948
rect 1636 26936 1642 26988
rect 5074 26976 5080 26988
rect 5035 26948 5080 26976
rect 5074 26936 5080 26948
rect 5132 26936 5138 26988
rect 5629 26979 5687 26985
rect 5629 26945 5641 26979
rect 5675 26945 5687 26979
rect 5629 26939 5687 26945
rect 5534 26868 5540 26920
rect 5592 26908 5598 26920
rect 5644 26908 5672 26939
rect 5592 26880 5672 26908
rect 5592 26868 5598 26880
rect 5166 26800 5172 26852
rect 5224 26840 5230 26852
rect 5810 26840 5816 26852
rect 5224 26812 5816 26840
rect 5224 26800 5230 26812
rect 5810 26800 5816 26812
rect 5868 26800 5874 26852
rect 1104 26682 6808 26704
rect 1104 26630 1915 26682
rect 1967 26630 1979 26682
rect 2031 26630 2043 26682
rect 2095 26630 2107 26682
rect 2159 26630 2171 26682
rect 2223 26630 3846 26682
rect 3898 26630 3910 26682
rect 3962 26630 3974 26682
rect 4026 26630 4038 26682
rect 4090 26630 4102 26682
rect 4154 26630 5776 26682
rect 5828 26630 5840 26682
rect 5892 26630 5904 26682
rect 5956 26630 5968 26682
rect 6020 26630 6032 26682
rect 6084 26630 6808 26682
rect 1104 26608 6808 26630
rect 1397 26571 1455 26577
rect 1397 26537 1409 26571
rect 1443 26568 1455 26571
rect 2406 26568 2412 26580
rect 1443 26540 2412 26568
rect 1443 26537 1455 26540
rect 1397 26531 1455 26537
rect 2406 26528 2412 26540
rect 2464 26528 2470 26580
rect 5258 26568 5264 26580
rect 5219 26540 5264 26568
rect 5258 26528 5264 26540
rect 5316 26528 5322 26580
rect 6178 26528 6184 26580
rect 6236 26568 6242 26580
rect 6546 26568 6552 26580
rect 6236 26540 6552 26568
rect 6236 26528 6242 26540
rect 6546 26528 6552 26540
rect 6604 26528 6610 26580
rect 5442 26460 5448 26512
rect 5500 26460 5506 26512
rect 5905 26503 5963 26509
rect 5905 26469 5917 26503
rect 5951 26500 5963 26503
rect 7653 26503 7711 26509
rect 7653 26500 7665 26503
rect 5951 26472 7665 26500
rect 5951 26469 5963 26472
rect 5905 26463 5963 26469
rect 7653 26469 7665 26472
rect 7699 26469 7711 26503
rect 7653 26463 7711 26469
rect 5258 26392 5264 26444
rect 5316 26432 5322 26444
rect 5460 26432 5488 26460
rect 5316 26404 5488 26432
rect 5316 26392 5322 26404
rect 1578 26364 1584 26376
rect 1539 26336 1584 26364
rect 1578 26324 1584 26336
rect 1636 26324 1642 26376
rect 5442 26364 5448 26376
rect 5403 26336 5448 26364
rect 5442 26324 5448 26336
rect 5500 26324 5506 26376
rect 6089 26367 6147 26373
rect 6089 26333 6101 26367
rect 6135 26333 6147 26367
rect 6089 26327 6147 26333
rect 6104 26228 6132 26327
rect 6822 26228 6828 26240
rect 6104 26200 6828 26228
rect 6822 26188 6828 26200
rect 6880 26188 6886 26240
rect 1104 26138 6808 26160
rect 1104 26086 2880 26138
rect 2932 26086 2944 26138
rect 2996 26086 3008 26138
rect 3060 26086 3072 26138
rect 3124 26086 3136 26138
rect 3188 26086 4811 26138
rect 4863 26086 4875 26138
rect 4927 26086 4939 26138
rect 4991 26086 5003 26138
rect 5055 26086 5067 26138
rect 5119 26086 6808 26138
rect 1104 26064 6808 26086
rect 1397 26027 1455 26033
rect 1397 25993 1409 26027
rect 1443 26024 1455 26027
rect 1670 26024 1676 26036
rect 1443 25996 1676 26024
rect 1443 25993 1455 25996
rect 1397 25987 1455 25993
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 4706 26024 4712 26036
rect 4667 25996 4712 26024
rect 4706 25984 4712 25996
rect 4764 25984 4770 26036
rect 3694 25916 3700 25968
rect 3752 25956 3758 25968
rect 5353 25959 5411 25965
rect 5353 25956 5365 25959
rect 3752 25928 5365 25956
rect 3752 25916 3758 25928
rect 5353 25925 5365 25928
rect 5399 25925 5411 25959
rect 5353 25919 5411 25925
rect 5537 25959 5595 25965
rect 5537 25925 5549 25959
rect 5583 25956 5595 25959
rect 7377 25959 7435 25965
rect 7377 25956 7389 25959
rect 5583 25928 7389 25956
rect 5583 25925 5595 25928
rect 5537 25919 5595 25925
rect 7377 25925 7389 25928
rect 7423 25925 7435 25959
rect 7377 25919 7435 25925
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 3510 25848 3516 25900
rect 3568 25888 3574 25900
rect 4617 25891 4675 25897
rect 4617 25888 4629 25891
rect 3568 25860 4629 25888
rect 3568 25848 3574 25860
rect 4617 25857 4629 25860
rect 4663 25857 4675 25891
rect 4617 25851 4675 25857
rect 4430 25780 4436 25832
rect 4488 25820 4494 25832
rect 4706 25820 4712 25832
rect 4488 25792 4712 25820
rect 4488 25780 4494 25792
rect 4706 25780 4712 25792
rect 4764 25780 4770 25832
rect 1104 25594 6808 25616
rect 1104 25542 1915 25594
rect 1967 25542 1979 25594
rect 2031 25542 2043 25594
rect 2095 25542 2107 25594
rect 2159 25542 2171 25594
rect 2223 25542 3846 25594
rect 3898 25542 3910 25594
rect 3962 25542 3974 25594
rect 4026 25542 4038 25594
rect 4090 25542 4102 25594
rect 4154 25542 5776 25594
rect 5828 25542 5840 25594
rect 5892 25542 5904 25594
rect 5956 25542 5968 25594
rect 6020 25542 6032 25594
rect 6084 25542 6808 25594
rect 1104 25520 6808 25542
rect 5905 25483 5963 25489
rect 5905 25449 5917 25483
rect 5951 25480 5963 25483
rect 7561 25483 7619 25489
rect 7561 25480 7573 25483
rect 5951 25452 7573 25480
rect 5951 25449 5963 25452
rect 5905 25443 5963 25449
rect 7561 25449 7573 25452
rect 7607 25449 7619 25483
rect 7561 25443 7619 25449
rect 5353 25415 5411 25421
rect 5353 25381 5365 25415
rect 5399 25412 5411 25415
rect 7469 25415 7527 25421
rect 7469 25412 7481 25415
rect 5399 25384 7481 25412
rect 5399 25381 5411 25384
rect 5353 25375 5411 25381
rect 7469 25381 7481 25384
rect 7515 25381 7527 25415
rect 7469 25375 7527 25381
rect 5166 25304 5172 25356
rect 5224 25344 5230 25356
rect 5442 25344 5448 25356
rect 5224 25316 5448 25344
rect 5224 25304 5230 25316
rect 5442 25304 5448 25316
rect 5500 25304 5506 25356
rect 6086 25276 6092 25288
rect 6047 25248 6092 25276
rect 6086 25236 6092 25248
rect 6144 25236 6150 25288
rect 5166 25208 5172 25220
rect 5127 25180 5172 25208
rect 5166 25168 5172 25180
rect 5224 25168 5230 25220
rect 1104 25050 6808 25072
rect 1104 24998 2880 25050
rect 2932 24998 2944 25050
rect 2996 24998 3008 25050
rect 3060 24998 3072 25050
rect 3124 24998 3136 25050
rect 3188 24998 4811 25050
rect 4863 24998 4875 25050
rect 4927 24998 4939 25050
rect 4991 24998 5003 25050
rect 5055 24998 5067 25050
rect 5119 24998 6808 25050
rect 1104 24976 6808 24998
rect 5629 24939 5687 24945
rect 5629 24905 5641 24939
rect 5675 24936 5687 24939
rect 7101 24939 7159 24945
rect 7101 24936 7113 24939
rect 5675 24908 7113 24936
rect 5675 24905 5687 24908
rect 5629 24899 5687 24905
rect 7101 24905 7113 24908
rect 7147 24905 7159 24939
rect 7101 24899 7159 24905
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24800 5871 24803
rect 6178 24800 6184 24812
rect 5859 24772 6184 24800
rect 5859 24769 5871 24772
rect 5813 24763 5871 24769
rect 6178 24760 6184 24772
rect 6236 24760 6242 24812
rect 1397 24667 1455 24673
rect 1397 24633 1409 24667
rect 1443 24664 1455 24667
rect 5534 24664 5540 24676
rect 1443 24636 5540 24664
rect 1443 24633 1455 24636
rect 1397 24627 1455 24633
rect 5534 24624 5540 24636
rect 5592 24624 5598 24676
rect 1104 24506 6808 24528
rect 1104 24454 1915 24506
rect 1967 24454 1979 24506
rect 2031 24454 2043 24506
rect 2095 24454 2107 24506
rect 2159 24454 2171 24506
rect 2223 24454 3846 24506
rect 3898 24454 3910 24506
rect 3962 24454 3974 24506
rect 4026 24454 4038 24506
rect 4090 24454 4102 24506
rect 4154 24454 5776 24506
rect 5828 24454 5840 24506
rect 5892 24454 5904 24506
rect 5956 24454 5968 24506
rect 6020 24454 6032 24506
rect 6084 24454 6808 24506
rect 1104 24432 6808 24454
rect 1486 24392 1492 24404
rect 1447 24364 1492 24392
rect 1486 24352 1492 24364
rect 1544 24352 1550 24404
rect 4341 24395 4399 24401
rect 4341 24361 4353 24395
rect 4387 24392 4399 24395
rect 4522 24392 4528 24404
rect 4387 24364 4528 24392
rect 4387 24361 4399 24364
rect 4341 24355 4399 24361
rect 4522 24352 4528 24364
rect 4580 24352 4586 24404
rect 5905 24395 5963 24401
rect 5905 24361 5917 24395
rect 5951 24392 5963 24395
rect 6917 24395 6975 24401
rect 6917 24392 6929 24395
rect 5951 24364 6929 24392
rect 5951 24361 5963 24364
rect 5905 24355 5963 24361
rect 6917 24361 6929 24364
rect 6963 24361 6975 24395
rect 6917 24355 6975 24361
rect 5261 24327 5319 24333
rect 5261 24324 5273 24327
rect 2746 24296 5273 24324
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24188 1731 24191
rect 2746 24188 2774 24296
rect 5261 24293 5273 24296
rect 5307 24293 5319 24327
rect 5261 24287 5319 24293
rect 5442 24188 5448 24200
rect 1719 24160 2774 24188
rect 5403 24160 5448 24188
rect 1719 24157 1731 24160
rect 1673 24151 1731 24157
rect 5442 24148 5448 24160
rect 5500 24148 5506 24200
rect 6089 24191 6147 24197
rect 6089 24157 6101 24191
rect 6135 24188 6147 24191
rect 6178 24188 6184 24200
rect 6135 24160 6184 24188
rect 6135 24157 6147 24160
rect 6089 24151 6147 24157
rect 6178 24148 6184 24160
rect 6236 24148 6242 24200
rect 2774 24080 2780 24132
rect 2832 24120 2838 24132
rect 4249 24123 4307 24129
rect 4249 24120 4261 24123
rect 2832 24092 4261 24120
rect 2832 24080 2838 24092
rect 4249 24089 4261 24092
rect 4295 24089 4307 24123
rect 4249 24083 4307 24089
rect 1104 23962 6808 23984
rect 1104 23910 2880 23962
rect 2932 23910 2944 23962
rect 2996 23910 3008 23962
rect 3060 23910 3072 23962
rect 3124 23910 3136 23962
rect 3188 23910 4811 23962
rect 4863 23910 4875 23962
rect 4927 23910 4939 23962
rect 4991 23910 5003 23962
rect 5055 23910 5067 23962
rect 5119 23910 6808 23962
rect 1104 23888 6808 23910
rect 1397 23851 1455 23857
rect 1397 23817 1409 23851
rect 1443 23848 1455 23851
rect 5166 23848 5172 23860
rect 1443 23820 5172 23848
rect 1443 23817 1455 23820
rect 1397 23811 1455 23817
rect 5166 23808 5172 23820
rect 5224 23808 5230 23860
rect 1578 23712 1584 23724
rect 1539 23684 1584 23712
rect 1578 23672 1584 23684
rect 1636 23672 1642 23724
rect 5166 23712 5172 23724
rect 5127 23684 5172 23712
rect 5166 23672 5172 23684
rect 5224 23672 5230 23724
rect 5629 23715 5687 23721
rect 5629 23681 5641 23715
rect 5675 23712 5687 23715
rect 7193 23715 7251 23721
rect 7193 23712 7205 23715
rect 5675 23684 7205 23712
rect 5675 23681 5687 23684
rect 5629 23675 5687 23681
rect 7193 23681 7205 23684
rect 7239 23681 7251 23715
rect 7193 23675 7251 23681
rect 5537 23647 5595 23653
rect 5537 23613 5549 23647
rect 5583 23644 5595 23647
rect 7101 23647 7159 23653
rect 7101 23644 7113 23647
rect 5583 23616 7113 23644
rect 5583 23613 5595 23616
rect 5537 23607 5595 23613
rect 7101 23613 7113 23616
rect 7147 23613 7159 23647
rect 7101 23607 7159 23613
rect 5442 23508 5448 23520
rect 5403 23480 5448 23508
rect 5442 23468 5448 23480
rect 5500 23468 5506 23520
rect 5813 23511 5871 23517
rect 5813 23477 5825 23511
rect 5859 23508 5871 23511
rect 6822 23508 6828 23520
rect 5859 23480 6828 23508
rect 5859 23477 5871 23480
rect 5813 23471 5871 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 1104 23418 6808 23440
rect 1104 23366 1915 23418
rect 1967 23366 1979 23418
rect 2031 23366 2043 23418
rect 2095 23366 2107 23418
rect 2159 23366 2171 23418
rect 2223 23366 3846 23418
rect 3898 23366 3910 23418
rect 3962 23366 3974 23418
rect 4026 23366 4038 23418
rect 4090 23366 4102 23418
rect 4154 23366 5776 23418
rect 5828 23366 5840 23418
rect 5892 23366 5904 23418
rect 5956 23366 5968 23418
rect 6020 23366 6032 23418
rect 6084 23366 6808 23418
rect 1104 23344 6808 23366
rect 1397 23307 1455 23313
rect 1397 23273 1409 23307
rect 1443 23304 1455 23307
rect 3694 23304 3700 23316
rect 1443 23276 3700 23304
rect 1443 23273 1455 23276
rect 1397 23267 1455 23273
rect 3694 23264 3700 23276
rect 3752 23264 3758 23316
rect 4893 23307 4951 23313
rect 4893 23273 4905 23307
rect 4939 23304 4951 23307
rect 5534 23304 5540 23316
rect 4939 23276 5540 23304
rect 4939 23273 4951 23276
rect 4893 23267 4951 23273
rect 5534 23264 5540 23276
rect 5592 23264 5598 23316
rect 5813 23307 5871 23313
rect 5813 23273 5825 23307
rect 5859 23304 5871 23307
rect 6454 23304 6460 23316
rect 5859 23276 6460 23304
rect 5859 23273 5871 23276
rect 5813 23267 5871 23273
rect 6454 23264 6460 23276
rect 6512 23264 6518 23316
rect 3237 23239 3295 23245
rect 3237 23205 3249 23239
rect 3283 23236 3295 23239
rect 5258 23236 5264 23248
rect 3283 23208 5264 23236
rect 3283 23205 3295 23208
rect 3237 23199 3295 23205
rect 5258 23196 5264 23208
rect 5316 23196 5322 23248
rect 7745 23239 7803 23245
rect 7745 23236 7757 23239
rect 5460 23208 7757 23236
rect 4433 23171 4491 23177
rect 4433 23137 4445 23171
rect 4479 23168 4491 23171
rect 5460 23168 5488 23208
rect 7745 23205 7757 23208
rect 7791 23205 7803 23239
rect 7745 23199 7803 23205
rect 7377 23171 7435 23177
rect 7377 23168 7389 23171
rect 4479 23140 5488 23168
rect 5552 23140 7389 23168
rect 4479 23137 4491 23140
rect 4433 23131 4491 23137
rect 1578 23100 1584 23112
rect 1539 23072 1584 23100
rect 1578 23060 1584 23072
rect 1636 23060 1642 23112
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23100 5135 23103
rect 5258 23100 5264 23112
rect 5123 23072 5264 23100
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5552 23109 5580 23140
rect 7377 23137 7389 23140
rect 7423 23137 7435 23171
rect 7377 23131 7435 23137
rect 5537 23103 5595 23109
rect 5537 23069 5549 23103
rect 5583 23069 5595 23103
rect 5537 23063 5595 23069
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23069 5779 23103
rect 5721 23063 5779 23069
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23100 5871 23103
rect 6822 23100 6828 23112
rect 5859 23072 6828 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 3053 23035 3111 23041
rect 3053 23001 3065 23035
rect 3099 23032 3111 23035
rect 3234 23032 3240 23044
rect 3099 23004 3240 23032
rect 3099 23001 3111 23004
rect 3053 22995 3111 23001
rect 3234 22992 3240 23004
rect 3292 22992 3298 23044
rect 3418 22992 3424 23044
rect 3476 23032 3482 23044
rect 4249 23035 4307 23041
rect 4249 23032 4261 23035
rect 3476 23004 4261 23032
rect 3476 22992 3482 23004
rect 4249 23001 4261 23004
rect 4295 23001 4307 23035
rect 5736 23032 5764 23063
rect 6822 23060 6828 23072
rect 6880 23060 6886 23112
rect 6917 23035 6975 23041
rect 6917 23032 6929 23035
rect 5736 23004 6929 23032
rect 4249 22995 4307 23001
rect 6917 23001 6929 23004
rect 6963 23001 6975 23035
rect 6917 22995 6975 23001
rect 5997 22967 6055 22973
rect 5997 22933 6009 22967
rect 6043 22964 6055 22967
rect 7009 22967 7067 22973
rect 7009 22964 7021 22967
rect 6043 22936 7021 22964
rect 6043 22933 6055 22936
rect 5997 22927 6055 22933
rect 7009 22933 7021 22936
rect 7055 22933 7067 22967
rect 7009 22927 7067 22933
rect 1104 22874 6808 22896
rect 1104 22822 2880 22874
rect 2932 22822 2944 22874
rect 2996 22822 3008 22874
rect 3060 22822 3072 22874
rect 3124 22822 3136 22874
rect 3188 22822 4811 22874
rect 4863 22822 4875 22874
rect 4927 22822 4939 22874
rect 4991 22822 5003 22874
rect 5055 22822 5067 22874
rect 5119 22822 6808 22874
rect 1104 22800 6808 22822
rect 1397 22763 1455 22769
rect 1397 22729 1409 22763
rect 1443 22760 1455 22763
rect 3510 22760 3516 22772
rect 1443 22732 3516 22760
rect 1443 22729 1455 22732
rect 1397 22723 1455 22729
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 4985 22763 5043 22769
rect 4985 22729 4997 22763
rect 5031 22760 5043 22763
rect 5166 22760 5172 22772
rect 5031 22732 5172 22760
rect 5031 22729 5043 22732
rect 4985 22723 5043 22729
rect 5166 22720 5172 22732
rect 5224 22720 5230 22772
rect 5626 22760 5632 22772
rect 5587 22732 5632 22760
rect 5626 22720 5632 22732
rect 5684 22720 5690 22772
rect 1578 22624 1584 22636
rect 1539 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22584 1642 22636
rect 5166 22624 5172 22636
rect 5127 22596 5172 22624
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 6178 22624 6184 22636
rect 5859 22596 6184 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 6178 22584 6184 22596
rect 6236 22584 6242 22636
rect 1104 22330 6808 22352
rect 1104 22278 1915 22330
rect 1967 22278 1979 22330
rect 2031 22278 2043 22330
rect 2095 22278 2107 22330
rect 2159 22278 2171 22330
rect 2223 22278 3846 22330
rect 3898 22278 3910 22330
rect 3962 22278 3974 22330
rect 4026 22278 4038 22330
rect 4090 22278 4102 22330
rect 4154 22278 5776 22330
rect 5828 22278 5840 22330
rect 5892 22278 5904 22330
rect 5956 22278 5968 22330
rect 6020 22278 6032 22330
rect 6084 22278 6808 22330
rect 1104 22256 6808 22278
rect 5534 22176 5540 22228
rect 5592 22216 5598 22228
rect 5629 22219 5687 22225
rect 5629 22216 5641 22219
rect 5592 22188 5641 22216
rect 5592 22176 5598 22188
rect 5629 22185 5641 22188
rect 5675 22185 5687 22219
rect 5629 22179 5687 22185
rect 6089 22219 6147 22225
rect 6089 22185 6101 22219
rect 6135 22216 6147 22219
rect 6454 22216 6460 22228
rect 6135 22188 6460 22216
rect 6135 22185 6147 22188
rect 6089 22179 6147 22185
rect 6454 22176 6460 22188
rect 6512 22176 6518 22228
rect 4430 22040 4436 22092
rect 4488 22080 4494 22092
rect 4709 22083 4767 22089
rect 4709 22080 4721 22083
rect 4488 22052 4721 22080
rect 4488 22040 4494 22052
rect 4709 22049 4721 22052
rect 4755 22049 4767 22083
rect 4709 22043 4767 22049
rect 5813 22083 5871 22089
rect 5813 22049 5825 22083
rect 5859 22080 5871 22083
rect 6917 22083 6975 22089
rect 6917 22080 6929 22083
rect 5859 22052 6929 22080
rect 5859 22049 5871 22052
rect 5813 22043 5871 22049
rect 6917 22049 6929 22052
rect 6963 22049 6975 22083
rect 6917 22043 6975 22049
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 5905 22015 5963 22021
rect 5905 21981 5917 22015
rect 5951 22012 5963 22015
rect 7285 22015 7343 22021
rect 7285 22012 7297 22015
rect 5951 21984 7297 22012
rect 5951 21981 5963 21984
rect 5905 21975 5963 21981
rect 7285 21981 7297 21984
rect 7331 21981 7343 22015
rect 7285 21975 7343 21981
rect 4522 21944 4528 21956
rect 4483 21916 4528 21944
rect 4522 21904 4528 21916
rect 4580 21904 4586 21956
rect 5626 21944 5632 21956
rect 5587 21916 5632 21944
rect 5626 21904 5632 21916
rect 5684 21904 5690 21956
rect 1397 21879 1455 21885
rect 1397 21845 1409 21879
rect 1443 21876 1455 21879
rect 2774 21876 2780 21888
rect 1443 21848 2780 21876
rect 1443 21845 1455 21848
rect 1397 21839 1455 21845
rect 2774 21836 2780 21848
rect 2832 21836 2838 21888
rect 1104 21786 6808 21808
rect 1104 21734 2880 21786
rect 2932 21734 2944 21786
rect 2996 21734 3008 21786
rect 3060 21734 3072 21786
rect 3124 21734 3136 21786
rect 3188 21734 4811 21786
rect 4863 21734 4875 21786
rect 4927 21734 4939 21786
rect 4991 21734 5003 21786
rect 5055 21734 5067 21786
rect 5119 21734 6808 21786
rect 1104 21712 6808 21734
rect 5442 21632 5448 21684
rect 5500 21672 5506 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5500 21644 5641 21672
rect 5500 21632 5506 21644
rect 5629 21641 5641 21644
rect 5675 21641 5687 21675
rect 5629 21635 5687 21641
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 6178 21536 6184 21548
rect 5859 21508 6184 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 1104 21242 6808 21264
rect 1104 21190 1915 21242
rect 1967 21190 1979 21242
rect 2031 21190 2043 21242
rect 2095 21190 2107 21242
rect 2159 21190 2171 21242
rect 2223 21190 3846 21242
rect 3898 21190 3910 21242
rect 3962 21190 3974 21242
rect 4026 21190 4038 21242
rect 4090 21190 4102 21242
rect 4154 21190 5776 21242
rect 5828 21190 5840 21242
rect 5892 21190 5904 21242
rect 5956 21190 5968 21242
rect 6020 21190 6032 21242
rect 6084 21190 6808 21242
rect 1104 21168 6808 21190
rect 1397 21131 1455 21137
rect 1397 21097 1409 21131
rect 1443 21128 1455 21131
rect 4522 21128 4528 21140
rect 1443 21100 4528 21128
rect 1443 21097 1455 21100
rect 1397 21091 1455 21097
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 5905 21131 5963 21137
rect 5905 21097 5917 21131
rect 5951 21128 5963 21131
rect 7101 21131 7159 21137
rect 7101 21128 7113 21131
rect 5951 21100 7113 21128
rect 5951 21097 5963 21100
rect 5905 21091 5963 21097
rect 7101 21097 7113 21100
rect 7147 21097 7159 21131
rect 7101 21091 7159 21097
rect 1578 20924 1584 20936
rect 1539 20896 1584 20924
rect 1578 20884 1584 20896
rect 1636 20884 1642 20936
rect 6086 20924 6092 20936
rect 6047 20896 6092 20924
rect 6086 20884 6092 20896
rect 6144 20884 6150 20936
rect 1104 20698 6808 20720
rect 1104 20646 2880 20698
rect 2932 20646 2944 20698
rect 2996 20646 3008 20698
rect 3060 20646 3072 20698
rect 3124 20646 3136 20698
rect 3188 20646 4811 20698
rect 4863 20646 4875 20698
rect 4927 20646 4939 20698
rect 4991 20646 5003 20698
rect 5055 20646 5067 20698
rect 5119 20646 6808 20698
rect 1104 20624 6808 20646
rect 1397 20587 1455 20593
rect 1397 20553 1409 20587
rect 1443 20584 1455 20587
rect 1762 20584 1768 20596
rect 1443 20556 1768 20584
rect 1443 20553 1455 20556
rect 1397 20547 1455 20553
rect 1762 20544 1768 20556
rect 1820 20544 1826 20596
rect 5626 20584 5632 20596
rect 5587 20556 5632 20584
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 1578 20448 1584 20460
rect 1539 20420 1584 20448
rect 1578 20408 1584 20420
rect 1636 20408 1642 20460
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 6178 20448 6184 20460
rect 5859 20420 6184 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6178 20408 6184 20420
rect 6236 20408 6242 20460
rect 1104 20154 6808 20176
rect 1104 20102 1915 20154
rect 1967 20102 1979 20154
rect 2031 20102 2043 20154
rect 2095 20102 2107 20154
rect 2159 20102 2171 20154
rect 2223 20102 3846 20154
rect 3898 20102 3910 20154
rect 3962 20102 3974 20154
rect 4026 20102 4038 20154
rect 4090 20102 4102 20154
rect 4154 20102 5776 20154
rect 5828 20102 5840 20154
rect 5892 20102 5904 20154
rect 5956 20102 5968 20154
rect 6020 20102 6032 20154
rect 6084 20102 6808 20154
rect 1104 20080 6808 20102
rect 5905 20043 5963 20049
rect 5905 20009 5917 20043
rect 5951 20040 5963 20043
rect 7193 20043 7251 20049
rect 7193 20040 7205 20043
rect 5951 20012 7205 20040
rect 5951 20009 5963 20012
rect 5905 20003 5963 20009
rect 7193 20009 7205 20012
rect 7239 20009 7251 20043
rect 7193 20003 7251 20009
rect 2041 19975 2099 19981
rect 2041 19941 2053 19975
rect 2087 19972 2099 19975
rect 6730 19972 6736 19984
rect 2087 19944 6736 19972
rect 2087 19941 2099 19944
rect 2041 19935 2099 19941
rect 6730 19932 6736 19944
rect 6788 19932 6794 19984
rect 6086 19836 6092 19848
rect 6047 19808 6092 19836
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 1394 19728 1400 19780
rect 1452 19768 1458 19780
rect 1857 19771 1915 19777
rect 1857 19768 1869 19771
rect 1452 19740 1869 19768
rect 1452 19728 1458 19740
rect 1857 19737 1869 19740
rect 1903 19737 1915 19771
rect 1857 19731 1915 19737
rect 1104 19610 6808 19632
rect 1104 19558 2880 19610
rect 2932 19558 2944 19610
rect 2996 19558 3008 19610
rect 3060 19558 3072 19610
rect 3124 19558 3136 19610
rect 3188 19558 4811 19610
rect 4863 19558 4875 19610
rect 4927 19558 4939 19610
rect 4991 19558 5003 19610
rect 5055 19558 5067 19610
rect 5119 19558 6808 19610
rect 1104 19536 6808 19558
rect 1397 19499 1455 19505
rect 1397 19465 1409 19499
rect 1443 19496 1455 19499
rect 1443 19468 3372 19496
rect 1443 19465 1455 19468
rect 1397 19459 1455 19465
rect 3344 19437 3372 19468
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 5629 19499 5687 19505
rect 5629 19496 5641 19499
rect 5592 19468 5641 19496
rect 5592 19456 5598 19468
rect 5629 19465 5641 19468
rect 5675 19465 5687 19499
rect 5629 19459 5687 19465
rect 3329 19431 3387 19437
rect 3329 19397 3341 19431
rect 3375 19397 3387 19431
rect 3329 19391 3387 19397
rect 1578 19360 1584 19372
rect 1539 19332 1584 19360
rect 1578 19320 1584 19332
rect 1636 19320 1642 19372
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19329 5871 19363
rect 5813 19323 5871 19329
rect 5828 19292 5856 19323
rect 6454 19292 6460 19304
rect 5828 19264 6460 19292
rect 6454 19252 6460 19264
rect 6512 19252 6518 19304
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19224 3571 19227
rect 6362 19224 6368 19236
rect 3559 19196 6368 19224
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 1104 19066 6808 19088
rect 1104 19014 1915 19066
rect 1967 19014 1979 19066
rect 2031 19014 2043 19066
rect 2095 19014 2107 19066
rect 2159 19014 2171 19066
rect 2223 19014 3846 19066
rect 3898 19014 3910 19066
rect 3962 19014 3974 19066
rect 4026 19014 4038 19066
rect 4090 19014 4102 19066
rect 4154 19014 5776 19066
rect 5828 19014 5840 19066
rect 5892 19014 5904 19066
rect 5956 19014 5968 19066
rect 6020 19014 6032 19066
rect 6084 19014 6808 19066
rect 1104 18992 6808 19014
rect 1397 18955 1455 18961
rect 1397 18921 1409 18955
rect 1443 18952 1455 18955
rect 3234 18952 3240 18964
rect 1443 18924 3240 18952
rect 1443 18921 1455 18924
rect 1397 18915 1455 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 5905 18955 5963 18961
rect 5905 18921 5917 18955
rect 5951 18952 5963 18955
rect 6917 18955 6975 18961
rect 6917 18952 6929 18955
rect 5951 18924 6929 18952
rect 5951 18921 5963 18924
rect 5905 18915 5963 18921
rect 6917 18921 6929 18924
rect 6963 18921 6975 18955
rect 6917 18915 6975 18921
rect 1578 18748 1584 18760
rect 1539 18720 1584 18748
rect 1578 18708 1584 18720
rect 1636 18708 1642 18760
rect 6086 18748 6092 18760
rect 6047 18720 6092 18748
rect 6086 18708 6092 18720
rect 6144 18708 6150 18760
rect 1104 18522 6808 18544
rect 1104 18470 2880 18522
rect 2932 18470 2944 18522
rect 2996 18470 3008 18522
rect 3060 18470 3072 18522
rect 3124 18470 3136 18522
rect 3188 18470 4811 18522
rect 4863 18470 4875 18522
rect 4927 18470 4939 18522
rect 4991 18470 5003 18522
rect 5055 18470 5067 18522
rect 5119 18470 6808 18522
rect 1104 18448 6808 18470
rect 1397 18411 1455 18417
rect 1397 18377 1409 18411
rect 1443 18408 1455 18411
rect 3418 18408 3424 18420
rect 1443 18380 3424 18408
rect 1443 18377 1455 18380
rect 1397 18371 1455 18377
rect 3418 18368 3424 18380
rect 3476 18368 3482 18420
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 6178 18272 6184 18284
rect 5859 18244 6184 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 6178 18232 6184 18244
rect 6236 18232 6242 18284
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5592 18040 5641 18068
rect 5592 18028 5598 18040
rect 5629 18037 5641 18040
rect 5675 18037 5687 18071
rect 5629 18031 5687 18037
rect 1104 17978 6808 18000
rect 1104 17926 1915 17978
rect 1967 17926 1979 17978
rect 2031 17926 2043 17978
rect 2095 17926 2107 17978
rect 2159 17926 2171 17978
rect 2223 17926 3846 17978
rect 3898 17926 3910 17978
rect 3962 17926 3974 17978
rect 4026 17926 4038 17978
rect 4090 17926 4102 17978
rect 4154 17926 5776 17978
rect 5828 17926 5840 17978
rect 5892 17926 5904 17978
rect 5956 17926 5968 17978
rect 6020 17926 6032 17978
rect 6084 17926 6808 17978
rect 1104 17904 6808 17926
rect 4614 17864 4620 17876
rect 4575 17836 4620 17864
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5261 17867 5319 17873
rect 5261 17833 5273 17867
rect 5307 17864 5319 17867
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 5307 17836 7297 17864
rect 5307 17833 5319 17836
rect 5261 17827 5319 17833
rect 7285 17833 7297 17836
rect 7331 17833 7343 17867
rect 7285 17827 7343 17833
rect 5442 17660 5448 17672
rect 5403 17632 5448 17660
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 6089 17663 6147 17669
rect 6089 17629 6101 17663
rect 6135 17660 6147 17663
rect 6178 17660 6184 17672
rect 6135 17632 6184 17660
rect 6135 17629 6147 17632
rect 6089 17623 6147 17629
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 4522 17592 4528 17604
rect 4483 17564 4528 17592
rect 4522 17552 4528 17564
rect 4580 17552 4586 17604
rect 5905 17527 5963 17533
rect 5905 17493 5917 17527
rect 5951 17524 5963 17527
rect 6917 17527 6975 17533
rect 6917 17524 6929 17527
rect 5951 17496 6929 17524
rect 5951 17493 5963 17496
rect 5905 17487 5963 17493
rect 6917 17493 6929 17496
rect 6963 17493 6975 17527
rect 6917 17487 6975 17493
rect 1104 17434 6808 17456
rect 1104 17382 2880 17434
rect 2932 17382 2944 17434
rect 2996 17382 3008 17434
rect 3060 17382 3072 17434
rect 3124 17382 3136 17434
rect 3188 17382 4811 17434
rect 4863 17382 4875 17434
rect 4927 17382 4939 17434
rect 4991 17382 5003 17434
rect 5055 17382 5067 17434
rect 5119 17382 6808 17434
rect 1104 17360 6808 17382
rect 1394 17320 1400 17332
rect 1355 17292 1400 17320
rect 1394 17280 1400 17292
rect 1452 17280 1458 17332
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 4304 17292 4445 17320
rect 4304 17280 4310 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 4433 17283 4491 17289
rect 1578 17184 1584 17196
rect 1539 17156 1584 17184
rect 1578 17144 1584 17156
rect 1636 17144 1642 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4430 17184 4436 17196
rect 4387 17156 4436 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 4430 17144 4436 17156
rect 4488 17144 4494 17196
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6362 17184 6368 17196
rect 5859 17156 6368 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 5626 16980 5632 16992
rect 5587 16952 5632 16980
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 1104 16890 6808 16912
rect 1104 16838 1915 16890
rect 1967 16838 1979 16890
rect 2031 16838 2043 16890
rect 2095 16838 2107 16890
rect 2159 16838 2171 16890
rect 2223 16838 3846 16890
rect 3898 16838 3910 16890
rect 3962 16838 3974 16890
rect 4026 16838 4038 16890
rect 4090 16838 4102 16890
rect 4154 16838 5776 16890
rect 5828 16838 5840 16890
rect 5892 16838 5904 16890
rect 5956 16838 5968 16890
rect 6020 16838 6032 16890
rect 6084 16838 6808 16890
rect 1104 16816 6808 16838
rect 4338 16776 4344 16788
rect 4299 16748 4344 16776
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16776 5963 16779
rect 6917 16779 6975 16785
rect 6917 16776 6929 16779
rect 5951 16748 6929 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 6917 16745 6929 16748
rect 6963 16745 6975 16779
rect 6917 16739 6975 16745
rect 5810 16668 5816 16720
rect 5868 16708 5874 16720
rect 6638 16708 6644 16720
rect 5868 16680 6644 16708
rect 5868 16668 5874 16680
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 5626 16600 5632 16652
rect 5684 16640 5690 16652
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 5684 16612 5733 16640
rect 5684 16600 5690 16612
rect 5721 16609 5733 16612
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 1578 16572 1584 16584
rect 1539 16544 1584 16572
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 5258 16532 5264 16584
rect 5316 16572 5322 16584
rect 5905 16575 5963 16581
rect 5905 16572 5917 16575
rect 5316 16544 5917 16572
rect 5316 16532 5322 16544
rect 5905 16541 5917 16544
rect 5951 16541 5963 16575
rect 5905 16535 5963 16541
rect 4246 16504 4252 16516
rect 4207 16476 4252 16504
rect 4246 16464 4252 16476
rect 4304 16464 4310 16516
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 5629 16507 5687 16513
rect 5629 16504 5641 16507
rect 5592 16476 5641 16504
rect 5592 16464 5598 16476
rect 5629 16473 5641 16476
rect 5675 16473 5687 16507
rect 5629 16467 5687 16473
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 4430 16436 4436 16448
rect 1443 16408 4436 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 4430 16396 4436 16408
rect 4488 16396 4494 16448
rect 6089 16439 6147 16445
rect 6089 16405 6101 16439
rect 6135 16436 6147 16439
rect 6270 16436 6276 16448
rect 6135 16408 6276 16436
rect 6135 16405 6147 16408
rect 6089 16399 6147 16405
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 1104 16346 6808 16368
rect 1104 16294 2880 16346
rect 2932 16294 2944 16346
rect 2996 16294 3008 16346
rect 3060 16294 3072 16346
rect 3124 16294 3136 16346
rect 3188 16294 4811 16346
rect 4863 16294 4875 16346
rect 4927 16294 4939 16346
rect 4991 16294 5003 16346
rect 5055 16294 5067 16346
rect 5119 16294 6808 16346
rect 1104 16272 6808 16294
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5810 16232 5816 16244
rect 4939 16204 5816 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 4338 16056 4344 16108
rect 4396 16096 4402 16108
rect 4801 16099 4859 16105
rect 4801 16096 4813 16099
rect 4396 16068 4813 16096
rect 4396 16056 4402 16068
rect 4801 16065 4813 16068
rect 4847 16065 4859 16099
rect 4801 16059 4859 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6178 16096 6184 16108
rect 5859 16068 6184 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6178 16056 6184 16068
rect 6236 16056 6242 16108
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 1104 15802 6808 15824
rect 1104 15750 1915 15802
rect 1967 15750 1979 15802
rect 2031 15750 2043 15802
rect 2095 15750 2107 15802
rect 2159 15750 2171 15802
rect 2223 15750 3846 15802
rect 3898 15750 3910 15802
rect 3962 15750 3974 15802
rect 4026 15750 4038 15802
rect 4090 15750 4102 15802
rect 4154 15750 5776 15802
rect 5828 15750 5840 15802
rect 5892 15750 5904 15802
rect 5956 15750 5968 15802
rect 6020 15750 6032 15802
rect 6084 15750 6808 15802
rect 1104 15728 6808 15750
rect 1397 15691 1455 15697
rect 1397 15657 1409 15691
rect 1443 15688 1455 15691
rect 4522 15688 4528 15700
rect 1443 15660 4528 15688
rect 1443 15657 1455 15660
rect 1397 15651 1455 15657
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 5442 15484 5448 15496
rect 5403 15456 5448 15484
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15484 6147 15487
rect 6178 15484 6184 15496
rect 6135 15456 6184 15484
rect 6135 15453 6147 15456
rect 6089 15447 6147 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 5905 15351 5963 15357
rect 5905 15348 5917 15351
rect 5592 15320 5917 15348
rect 5592 15308 5598 15320
rect 5905 15317 5917 15320
rect 5951 15317 5963 15351
rect 5905 15311 5963 15317
rect 1104 15258 6808 15280
rect 1104 15206 2880 15258
rect 2932 15206 2944 15258
rect 2996 15206 3008 15258
rect 3060 15206 3072 15258
rect 3124 15206 3136 15258
rect 3188 15206 4811 15258
rect 4863 15206 4875 15258
rect 4927 15206 4939 15258
rect 4991 15206 5003 15258
rect 5055 15206 5067 15258
rect 5119 15206 6808 15258
rect 1104 15184 6808 15206
rect 1397 15147 1455 15153
rect 1397 15113 1409 15147
rect 1443 15144 1455 15147
rect 4246 15144 4252 15156
rect 1443 15116 4252 15144
rect 1443 15113 1455 15116
rect 1397 15107 1455 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 5813 15147 5871 15153
rect 5813 15113 5825 15147
rect 5859 15144 5871 15147
rect 7377 15147 7435 15153
rect 7377 15144 7389 15147
rect 5859 15116 7389 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 7377 15113 7389 15116
rect 7423 15113 7435 15147
rect 7377 15107 7435 15113
rect 1578 15008 1584 15020
rect 1539 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 5350 15008 5356 15020
rect 5311 14980 5356 15008
rect 5350 14968 5356 14980
rect 5408 14968 5414 15020
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 6917 15011 6975 15017
rect 6917 15008 6929 15011
rect 5675 14980 6929 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 6917 14977 6929 14980
rect 6963 14977 6975 15011
rect 6917 14971 6975 14977
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14940 5595 14943
rect 6270 14940 6276 14952
rect 5583 14912 6276 14940
rect 5583 14909 5595 14912
rect 5537 14903 5595 14909
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 5629 14807 5687 14813
rect 5629 14773 5641 14807
rect 5675 14804 5687 14807
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 5675 14776 7297 14804
rect 5675 14773 5687 14776
rect 5629 14767 5687 14773
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 1104 14714 6808 14736
rect 1104 14662 1915 14714
rect 1967 14662 1979 14714
rect 2031 14662 2043 14714
rect 2095 14662 2107 14714
rect 2159 14662 2171 14714
rect 2223 14662 3846 14714
rect 3898 14662 3910 14714
rect 3962 14662 3974 14714
rect 4026 14662 4038 14714
rect 4090 14662 4102 14714
rect 4154 14662 5776 14714
rect 5828 14662 5840 14714
rect 5892 14662 5904 14714
rect 5956 14662 5968 14714
rect 6020 14662 6032 14714
rect 6084 14662 6808 14714
rect 1104 14640 6808 14662
rect 1397 14603 1455 14609
rect 1397 14569 1409 14603
rect 1443 14600 1455 14603
rect 4338 14600 4344 14612
rect 1443 14572 4344 14600
rect 1443 14569 1455 14572
rect 1397 14563 1455 14569
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5592 14572 5641 14600
rect 5592 14560 5598 14572
rect 5629 14569 5641 14572
rect 5675 14569 5687 14603
rect 5629 14563 5687 14569
rect 5350 14492 5356 14544
rect 5408 14532 5414 14544
rect 6089 14535 6147 14541
rect 6089 14532 6101 14535
rect 5408 14504 6101 14532
rect 5408 14492 5414 14504
rect 6089 14501 6101 14504
rect 6135 14501 6147 14535
rect 6089 14495 6147 14501
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 5626 14396 5632 14408
rect 5587 14368 5632 14396
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 5810 14396 5816 14408
rect 5771 14368 5816 14396
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 5905 14359 5963 14365
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 5920 14260 5948 14359
rect 5684 14232 5948 14260
rect 5684 14220 5690 14232
rect 1104 14170 6808 14192
rect 1104 14118 2880 14170
rect 2932 14118 2944 14170
rect 2996 14118 3008 14170
rect 3060 14118 3072 14170
rect 3124 14118 3136 14170
rect 3188 14118 4811 14170
rect 4863 14118 4875 14170
rect 4927 14118 4939 14170
rect 4991 14118 5003 14170
rect 5055 14118 5067 14170
rect 5119 14118 6808 14170
rect 1104 14096 6808 14118
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 5810 14056 5816 14068
rect 5675 14028 5816 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 3329 13991 3387 13997
rect 3329 13957 3341 13991
rect 3375 13988 3387 13991
rect 6546 13988 6552 14000
rect 3375 13960 6552 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 3142 13920 3148 13932
rect 3103 13892 3148 13920
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 5810 13920 5816 13932
rect 5771 13892 5816 13920
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 1104 13626 6808 13648
rect 1104 13574 1915 13626
rect 1967 13574 1979 13626
rect 2031 13574 2043 13626
rect 2095 13574 2107 13626
rect 2159 13574 2171 13626
rect 2223 13574 3846 13626
rect 3898 13574 3910 13626
rect 3962 13574 3974 13626
rect 4026 13574 4038 13626
rect 4090 13574 4102 13626
rect 4154 13574 5776 13626
rect 5828 13574 5840 13626
rect 5892 13574 5904 13626
rect 5956 13574 5968 13626
rect 6020 13574 6032 13626
rect 6084 13574 6808 13626
rect 1104 13552 6808 13574
rect 1397 13515 1455 13521
rect 1397 13481 1409 13515
rect 1443 13512 1455 13515
rect 3142 13512 3148 13524
rect 1443 13484 3148 13512
rect 1443 13481 1455 13484
rect 1397 13475 1455 13481
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 4433 13447 4491 13453
rect 4433 13413 4445 13447
rect 4479 13444 4491 13447
rect 6454 13444 6460 13456
rect 4479 13416 6460 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 6454 13404 6460 13416
rect 6512 13404 6518 13456
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 6086 13308 6092 13320
rect 6047 13280 6092 13308
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 1452 13212 4261 13240
rect 1452 13200 1458 13212
rect 4249 13209 4261 13212
rect 4295 13209 4307 13243
rect 4249 13203 4307 13209
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 5905 13175 5963 13181
rect 5905 13172 5917 13175
rect 5592 13144 5917 13172
rect 5592 13132 5598 13144
rect 5905 13141 5917 13144
rect 5951 13141 5963 13175
rect 5905 13135 5963 13141
rect 1104 13082 6808 13104
rect 1104 13030 2880 13082
rect 2932 13030 2944 13082
rect 2996 13030 3008 13082
rect 3060 13030 3072 13082
rect 3124 13030 3136 13082
rect 3188 13030 4811 13082
rect 4863 13030 4875 13082
rect 4927 13030 4939 13082
rect 4991 13030 5003 13082
rect 5055 13030 5067 13082
rect 5119 13030 6808 13082
rect 1104 13008 6808 13030
rect 1394 12968 1400 12980
rect 1355 12940 1400 12968
rect 1394 12928 1400 12940
rect 1452 12928 1458 12980
rect 5626 12968 5632 12980
rect 5587 12940 5632 12968
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 5166 12900 5172 12912
rect 5127 12872 5172 12900
rect 5166 12860 5172 12872
rect 5224 12860 5230 12912
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 4304 12804 4997 12832
rect 4304 12792 4310 12804
rect 4985 12801 4997 12804
rect 5031 12801 5043 12835
rect 5810 12832 5816 12844
rect 5771 12804 5816 12832
rect 4985 12795 5043 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 1104 12538 6808 12560
rect 1104 12486 1915 12538
rect 1967 12486 1979 12538
rect 2031 12486 2043 12538
rect 2095 12486 2107 12538
rect 2159 12486 2171 12538
rect 2223 12486 3846 12538
rect 3898 12486 3910 12538
rect 3962 12486 3974 12538
rect 4026 12486 4038 12538
rect 4090 12486 4102 12538
rect 4154 12486 5776 12538
rect 5828 12486 5840 12538
rect 5892 12486 5904 12538
rect 5956 12486 5968 12538
rect 6020 12486 6032 12538
rect 6084 12486 6808 12538
rect 1104 12464 6808 12486
rect 6086 12220 6092 12232
rect 6047 12192 6092 12220
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 5905 12087 5963 12093
rect 5905 12084 5917 12087
rect 5684 12056 5917 12084
rect 5684 12044 5690 12056
rect 5905 12053 5917 12056
rect 5951 12053 5963 12087
rect 5905 12047 5963 12053
rect 1104 11994 6808 12016
rect 1104 11942 2880 11994
rect 2932 11942 2944 11994
rect 2996 11942 3008 11994
rect 3060 11942 3072 11994
rect 3124 11942 3136 11994
rect 3188 11942 4811 11994
rect 4863 11942 4875 11994
rect 4927 11942 4939 11994
rect 4991 11942 5003 11994
rect 5055 11942 5067 11994
rect 5119 11942 6808 11994
rect 1104 11920 6808 11942
rect 1397 11883 1455 11889
rect 1397 11849 1409 11883
rect 1443 11880 1455 11883
rect 4246 11880 4252 11892
rect 1443 11852 4252 11880
rect 1443 11849 1455 11852
rect 1397 11843 1455 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 6917 11883 6975 11889
rect 6917 11880 6929 11883
rect 5859 11852 6929 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 6917 11849 6929 11852
rect 6963 11849 6975 11883
rect 6917 11843 6975 11849
rect 5353 11815 5411 11821
rect 5353 11781 5365 11815
rect 5399 11812 5411 11815
rect 5534 11812 5540 11824
rect 5399 11784 5540 11812
rect 5399 11781 5411 11784
rect 5353 11775 5411 11781
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 5629 11747 5687 11753
rect 5629 11744 5641 11747
rect 5500 11716 5641 11744
rect 5500 11704 5506 11716
rect 5629 11713 5641 11716
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 5534 11676 5540 11688
rect 5495 11648 5540 11676
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 5626 11540 5632 11552
rect 5587 11512 5632 11540
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 1104 11450 6808 11472
rect 1104 11398 1915 11450
rect 1967 11398 1979 11450
rect 2031 11398 2043 11450
rect 2095 11398 2107 11450
rect 2159 11398 2171 11450
rect 2223 11398 3846 11450
rect 3898 11398 3910 11450
rect 3962 11398 3974 11450
rect 4026 11398 4038 11450
rect 4090 11398 4102 11450
rect 4154 11398 5776 11450
rect 5828 11398 5840 11450
rect 5892 11398 5904 11450
rect 5956 11398 5968 11450
rect 6020 11398 6032 11450
rect 6084 11398 6808 11450
rect 1104 11376 6808 11398
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5442 11336 5448 11348
rect 5307 11308 5448 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5905 11339 5963 11345
rect 5905 11336 5917 11339
rect 5592 11308 5917 11336
rect 5592 11296 5598 11308
rect 5905 11305 5917 11308
rect 5951 11305 5963 11339
rect 5905 11299 5963 11305
rect 4617 11271 4675 11277
rect 4617 11237 4629 11271
rect 4663 11268 4675 11271
rect 7193 11271 7251 11277
rect 7193 11268 7205 11271
rect 4663 11240 7205 11268
rect 4663 11237 4675 11240
rect 4617 11231 4675 11237
rect 7193 11237 7205 11240
rect 7239 11237 7251 11271
rect 7193 11231 7251 11237
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 4246 11132 4252 11144
rect 1443 11104 4252 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4798 11132 4804 11144
rect 4759 11104 4804 11132
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 5408 11104 5457 11132
rect 5408 11092 5414 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6178 11132 6184 11144
rect 6135 11104 6184 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 1104 10906 6808 10928
rect 1104 10854 2880 10906
rect 2932 10854 2944 10906
rect 2996 10854 3008 10906
rect 3060 10854 3072 10906
rect 3124 10854 3136 10906
rect 3188 10854 4811 10906
rect 4863 10854 4875 10906
rect 4927 10854 4939 10906
rect 4991 10854 5003 10906
rect 5055 10854 5067 10906
rect 5119 10854 6808 10906
rect 1104 10832 6808 10854
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10761 5319 10795
rect 5261 10755 5319 10761
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 5276 10656 5304 10755
rect 5442 10656 5448 10668
rect 4479 10628 5304 10656
rect 5403 10628 5448 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 1104 10362 6808 10384
rect 1104 10310 1915 10362
rect 1967 10310 1979 10362
rect 2031 10310 2043 10362
rect 2095 10310 2107 10362
rect 2159 10310 2171 10362
rect 2223 10310 3846 10362
rect 3898 10310 3910 10362
rect 3962 10310 3974 10362
rect 4026 10310 4038 10362
rect 4090 10310 4102 10362
rect 4154 10310 5776 10362
rect 5828 10310 5840 10362
rect 5892 10310 5904 10362
rect 5956 10310 5968 10362
rect 6020 10310 6032 10362
rect 6084 10310 6808 10362
rect 1104 10288 6808 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 1452 10220 3801 10248
rect 1452 10208 1458 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 5166 10044 5172 10056
rect 4019 10016 5028 10044
rect 5127 10016 5172 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 5000 9917 5028 10016
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 5859 10016 6929 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 4985 9911 5043 9917
rect 4985 9877 4997 9911
rect 5031 9877 5043 9911
rect 5626 9908 5632 9920
rect 5587 9880 5632 9908
rect 4985 9871 5043 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 1104 9818 6808 9840
rect 1104 9766 2880 9818
rect 2932 9766 2944 9818
rect 2996 9766 3008 9818
rect 3060 9766 3072 9818
rect 3124 9766 3136 9818
rect 3188 9766 4811 9818
rect 4863 9766 4875 9818
rect 4927 9766 4939 9818
rect 4991 9766 5003 9818
rect 5055 9766 5067 9818
rect 5119 9766 6808 9818
rect 1104 9744 6808 9766
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 5442 9568 5448 9580
rect 5403 9540 5448 9568
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 4304 9336 5273 9364
rect 4304 9324 4310 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5261 9327 5319 9333
rect 1104 9274 6808 9296
rect 1104 9222 1915 9274
rect 1967 9222 1979 9274
rect 2031 9222 2043 9274
rect 2095 9222 2107 9274
rect 2159 9222 2171 9274
rect 2223 9222 3846 9274
rect 3898 9222 3910 9274
rect 3962 9222 3974 9274
rect 4026 9222 4038 9274
rect 4090 9222 4102 9274
rect 4154 9222 5776 9274
rect 5828 9222 5840 9274
rect 5892 9222 5904 9274
rect 5956 9222 5968 9274
rect 6020 9222 6032 9274
rect 6084 9222 6808 9274
rect 1104 9200 6808 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 2133 9163 2191 9169
rect 2133 9160 2145 9163
rect 1452 9132 2145 9160
rect 1452 9120 1458 9132
rect 2133 9129 2145 9132
rect 2179 9129 2191 9163
rect 2133 9123 2191 9129
rect 5626 9024 5632 9036
rect 2332 8996 5632 9024
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 2332 8965 2360 8996
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5408 8928 5457 8956
rect 5408 8916 5414 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 6135 8928 7113 8956
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 4580 8792 5273 8820
rect 4580 8780 4586 8792
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 5261 8783 5319 8789
rect 5905 8823 5963 8829
rect 5905 8789 5917 8823
rect 5951 8820 5963 8823
rect 6178 8820 6184 8832
rect 5951 8792 6184 8820
rect 5951 8789 5963 8792
rect 5905 8783 5963 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 1104 8730 6808 8752
rect 1104 8678 2880 8730
rect 2932 8678 2944 8730
rect 2996 8678 3008 8730
rect 3060 8678 3072 8730
rect 3124 8678 3136 8730
rect 3188 8678 4811 8730
rect 4863 8678 4875 8730
rect 4927 8678 4939 8730
rect 4991 8678 5003 8730
rect 5055 8678 5067 8730
rect 5119 8678 6808 8730
rect 1104 8656 6808 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 3605 8619 3663 8625
rect 3605 8616 3617 8619
rect 1452 8588 3617 8616
rect 1452 8576 1458 8588
rect 3605 8585 3617 8588
rect 3651 8585 3663 8619
rect 3605 8579 3663 8585
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 4246 8480 4252 8492
rect 3835 8452 4252 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4700 8483 4758 8489
rect 4700 8449 4712 8483
rect 4746 8480 4758 8483
rect 5258 8480 5264 8492
rect 4746 8452 5264 8480
rect 4746 8449 4758 8452
rect 4700 8443 4758 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 4430 8412 4436 8424
rect 4391 8384 4436 8412
rect 4430 8372 4436 8384
rect 4488 8372 4494 8424
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 5813 8279 5871 8285
rect 5813 8276 5825 8279
rect 5500 8248 5825 8276
rect 5500 8236 5506 8248
rect 5813 8245 5825 8248
rect 5859 8245 5871 8279
rect 5813 8239 5871 8245
rect 1104 8186 6808 8208
rect 1104 8134 1915 8186
rect 1967 8134 1979 8186
rect 2031 8134 2043 8186
rect 2095 8134 2107 8186
rect 2159 8134 2171 8186
rect 2223 8134 3846 8186
rect 3898 8134 3910 8186
rect 3962 8134 3974 8186
rect 4026 8134 4038 8186
rect 4090 8134 4102 8186
rect 4154 8134 5776 8186
rect 5828 8134 5840 8186
rect 5892 8134 5904 8186
rect 5956 8134 5968 8186
rect 6020 8134 6032 8186
rect 6084 8134 6808 8186
rect 1104 8112 6808 8134
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 7009 8007 7067 8013
rect 7009 7973 7021 8007
rect 7055 7973 7067 8007
rect 7009 7967 7067 7973
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 5276 7908 6929 7936
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 5166 7868 5172 7880
rect 4847 7840 5172 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5276 7877 5304 7908
rect 6917 7905 6929 7908
rect 6963 7936 6975 7939
rect 7024 7936 7052 7967
rect 6963 7908 7052 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5442 7868 5448 7880
rect 5403 7840 5448 7868
rect 5261 7831 5319 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6135 7840 7021 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 4617 7735 4675 7741
rect 4617 7732 4629 7735
rect 4396 7704 4629 7732
rect 4396 7692 4402 7704
rect 4617 7701 4629 7704
rect 4663 7701 4675 7735
rect 4617 7695 4675 7701
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 6270 7732 6276 7744
rect 5951 7704 6276 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 1104 7642 6808 7664
rect 1104 7590 2880 7642
rect 2932 7590 2944 7642
rect 2996 7590 3008 7642
rect 3060 7590 3072 7642
rect 3124 7590 3136 7642
rect 3188 7590 4811 7642
rect 4863 7590 4875 7642
rect 4927 7590 4939 7642
rect 4991 7590 5003 7642
rect 5055 7590 5067 7642
rect 5119 7590 6808 7642
rect 1104 7568 6808 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 1452 7500 3157 7528
rect 1452 7488 1458 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4488 7500 4629 7528
rect 4488 7488 4494 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 4617 7491 4675 7497
rect 4522 7460 4528 7472
rect 3344 7432 4528 7460
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 3234 7392 3240 7404
rect 1443 7364 3240 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 3344 7401 3372 7432
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 4246 7392 4252 7404
rect 3835 7364 4252 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4430 7392 4436 7404
rect 4391 7364 4436 7392
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5442 7392 5448 7404
rect 5123 7364 5448 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 3752 7160 3893 7188
rect 3752 7148 3758 7160
rect 3881 7157 3893 7160
rect 3927 7157 3939 7191
rect 3881 7151 3939 7157
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7188 5227 7191
rect 5350 7188 5356 7200
rect 5215 7160 5356 7188
rect 5215 7157 5227 7160
rect 5169 7151 5227 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 1104 7098 6808 7120
rect 1104 7046 1915 7098
rect 1967 7046 1979 7098
rect 2031 7046 2043 7098
rect 2095 7046 2107 7098
rect 2159 7046 2171 7098
rect 2223 7046 3846 7098
rect 3898 7046 3910 7098
rect 3962 7046 3974 7098
rect 4026 7046 4038 7098
rect 4090 7046 4102 7098
rect 4154 7046 5776 7098
rect 5828 7046 5840 7098
rect 5892 7046 5904 7098
rect 5956 7046 5968 7098
rect 6020 7046 6032 7098
rect 6084 7046 6808 7098
rect 1104 7024 6808 7046
rect 7006 7012 7012 7064
rect 7064 7052 7070 7064
rect 7101 7055 7159 7061
rect 7101 7052 7113 7055
rect 7064 7024 7113 7052
rect 7064 7012 7070 7024
rect 7101 7021 7113 7024
rect 7147 7021 7159 7055
rect 7101 7015 7159 7021
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 3292 6956 3801 6984
rect 3292 6944 3298 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 3789 6947 3847 6953
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4985 6987 5043 6993
rect 4985 6984 4997 6987
rect 4304 6956 4997 6984
rect 4304 6944 4310 6956
rect 4985 6953 4997 6956
rect 5031 6953 5043 6987
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 4985 6947 5043 6953
rect 5460 6956 6929 6984
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 3988 6644 4016 6743
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 4893 6715 4951 6721
rect 4893 6712 4905 6715
rect 4764 6684 4905 6712
rect 4764 6672 4770 6684
rect 4893 6681 4905 6684
rect 4939 6681 4951 6715
rect 5460 6712 5488 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 5813 6919 5871 6925
rect 5813 6916 5825 6919
rect 5684 6888 5825 6916
rect 5684 6876 5690 6888
rect 5813 6885 5825 6888
rect 5859 6885 5871 6919
rect 5813 6879 5871 6885
rect 7101 6919 7159 6925
rect 7101 6885 7113 6919
rect 7147 6916 7159 6919
rect 7285 6919 7343 6925
rect 7285 6916 7297 6919
rect 7147 6888 7297 6916
rect 7147 6885 7159 6888
rect 7101 6879 7159 6885
rect 7285 6885 7297 6888
rect 7331 6885 7343 6919
rect 7285 6879 7343 6885
rect 5537 6715 5595 6721
rect 5537 6712 5549 6715
rect 5460 6684 5549 6712
rect 4893 6675 4951 6681
rect 5537 6681 5549 6684
rect 5583 6681 5595 6715
rect 6178 6712 6184 6724
rect 5537 6675 5595 6681
rect 5920 6684 6184 6712
rect 5920 6644 5948 6684
rect 6178 6672 6184 6684
rect 6236 6672 6242 6724
rect 3988 6616 5948 6644
rect 5997 6647 6055 6653
rect 5997 6613 6009 6647
rect 6043 6644 6055 6647
rect 6917 6647 6975 6653
rect 6917 6644 6929 6647
rect 6043 6616 6929 6644
rect 6043 6613 6055 6616
rect 5997 6607 6055 6613
rect 6917 6613 6929 6616
rect 6963 6613 6975 6647
rect 6917 6607 6975 6613
rect 1104 6554 6808 6576
rect 1104 6502 2880 6554
rect 2932 6502 2944 6554
rect 2996 6502 3008 6554
rect 3060 6502 3072 6554
rect 3124 6502 3136 6554
rect 3188 6502 4811 6554
rect 4863 6502 4875 6554
rect 4927 6502 4939 6554
rect 4991 6502 5003 6554
rect 5055 6502 5067 6554
rect 5119 6502 6808 6554
rect 1104 6480 6808 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 2869 6443 2927 6449
rect 2869 6440 2881 6443
rect 1452 6412 2881 6440
rect 1452 6400 1458 6412
rect 2869 6409 2881 6412
rect 2915 6409 2927 6443
rect 2869 6403 2927 6409
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4430 6440 4436 6452
rect 4203 6412 4436 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 4338 6372 4344 6384
rect 3068 6344 4344 6372
rect 3068 6313 3096 6344
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 3973 6307 4031 6313
rect 3973 6304 3985 6307
rect 3752 6276 3985 6304
rect 3752 6264 3758 6276
rect 3973 6273 3985 6276
rect 4019 6273 4031 6307
rect 4614 6304 4620 6316
rect 4575 6276 4620 6304
rect 3973 6267 4031 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 5442 6304 5448 6316
rect 5403 6276 5448 6304
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 4522 6128 4528 6180
rect 4580 6168 4586 6180
rect 5261 6171 5319 6177
rect 5261 6168 5273 6171
rect 4580 6140 5273 6168
rect 4580 6128 4586 6140
rect 5261 6137 5273 6140
rect 5307 6137 5319 6171
rect 5261 6131 5319 6137
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4488 6072 4721 6100
rect 4488 6060 4494 6072
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 4709 6063 4767 6069
rect 1104 6010 6808 6032
rect 1104 5958 1915 6010
rect 1967 5958 1979 6010
rect 2031 5958 2043 6010
rect 2095 5958 2107 6010
rect 2159 5958 2171 6010
rect 2223 5958 3846 6010
rect 3898 5958 3910 6010
rect 3962 5958 3974 6010
rect 4026 5958 4038 6010
rect 4090 5958 4102 6010
rect 4154 5958 5776 6010
rect 5828 5958 5840 6010
rect 5892 5958 5904 6010
rect 5956 5958 5968 6010
rect 6020 5958 6032 6010
rect 6084 5958 6808 6010
rect 7006 5964 7012 5976
rect 1104 5936 6808 5958
rect 6967 5936 7012 5964
rect 7006 5924 7012 5936
rect 7064 5924 7070 5976
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 3237 5695 3295 5701
rect 1443 5664 3096 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 3068 5565 3096 5664
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 6270 5692 6276 5704
rect 3283 5664 6276 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 4246 5624 4252 5636
rect 4203 5596 4252 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 3053 5559 3111 5565
rect 3053 5525 3065 5559
rect 3099 5525 3111 5559
rect 3053 5519 3111 5525
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 4764 5528 5457 5556
rect 4764 5516 4770 5528
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 5445 5519 5503 5525
rect 1104 5466 6808 5488
rect 1104 5414 2880 5466
rect 2932 5414 2944 5466
rect 2996 5414 3008 5466
rect 3060 5414 3072 5466
rect 3124 5414 3136 5466
rect 3188 5414 4811 5466
rect 4863 5414 4875 5466
rect 4927 5414 4939 5466
rect 4991 5414 5003 5466
rect 5055 5414 5067 5466
rect 5119 5414 6808 5466
rect 1104 5392 6808 5414
rect 2133 5355 2191 5361
rect 2133 5321 2145 5355
rect 2179 5321 2191 5355
rect 2133 5315 2191 5321
rect 3421 5355 3479 5361
rect 3421 5321 3433 5355
rect 3467 5321 3479 5355
rect 3421 5315 3479 5321
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 2148 5216 2176 5315
rect 1443 5188 2176 5216
rect 2317 5219 2375 5225
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 3436 5216 3464 5315
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5684 5324 5825 5352
rect 5684 5312 5690 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 4700 5287 4758 5293
rect 4700 5253 4712 5287
rect 4746 5284 4758 5287
rect 4798 5284 4804 5296
rect 4746 5256 4804 5284
rect 4746 5253 4758 5256
rect 4700 5247 4758 5253
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 3602 5216 3608 5228
rect 2363 5188 3464 5216
rect 3563 5188 3608 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4430 5216 4436 5228
rect 4391 5188 4436 5216
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 1104 4922 6808 4944
rect 1104 4870 1915 4922
rect 1967 4870 1979 4922
rect 2031 4870 2043 4922
rect 2095 4870 2107 4922
rect 2159 4870 2171 4922
rect 2223 4870 3846 4922
rect 3898 4870 3910 4922
rect 3962 4870 3974 4922
rect 4026 4870 4038 4922
rect 4090 4870 4102 4922
rect 4154 4870 5776 4922
rect 5828 4870 5840 4922
rect 5892 4870 5904 4922
rect 5956 4870 5968 4922
rect 6020 4870 6032 4922
rect 6084 4870 6808 4922
rect 1104 4848 6808 4870
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4808 4767 4811
rect 4798 4808 4804 4820
rect 4755 4780 4804 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5905 4811 5963 4817
rect 5905 4777 5917 4811
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 6089 4811 6147 4817
rect 6089 4777 6101 4811
rect 6135 4808 6147 4811
rect 7101 4811 7159 4817
rect 7101 4808 7113 4811
rect 6135 4780 7113 4808
rect 6135 4777 6147 4780
rect 6089 4771 6147 4777
rect 7101 4777 7113 4780
rect 7147 4777 7159 4811
rect 7101 4771 7159 4777
rect 5920 4740 5948 4771
rect 7193 4743 7251 4749
rect 7193 4740 7205 4743
rect 5920 4712 7205 4740
rect 7193 4709 7205 4712
rect 7239 4709 7251 4743
rect 7193 4703 7251 4709
rect 4430 4672 4436 4684
rect 2516 4644 4436 4672
rect 2516 4613 2544 4644
rect 4430 4632 4436 4644
rect 4488 4632 4494 4684
rect 5166 4672 5172 4684
rect 4724 4644 5172 4672
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4338 4604 4344 4616
rect 4295 4576 4344 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 1780 4536 1808 4567
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 4724 4613 4752 4644
rect 5166 4632 5172 4644
rect 5224 4672 5230 4684
rect 5350 4672 5356 4684
rect 5224 4644 5356 4672
rect 5224 4632 5230 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 5442 4604 5448 4616
rect 5403 4576 5448 4604
rect 4893 4567 4951 4573
rect 4614 4536 4620 4548
rect 1780 4508 4620 4536
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 4908 4536 4936 4567
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5905 4607 5963 4613
rect 5592 4576 5637 4604
rect 5592 4564 5598 4576
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 5350 4536 5356 4548
rect 4908 4508 5356 4536
rect 5350 4496 5356 4508
rect 5408 4536 5414 4548
rect 5920 4536 5948 4567
rect 5408 4508 5948 4536
rect 5408 4496 5414 4508
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 2314 4468 2320 4480
rect 1995 4440 2320 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2590 4468 2596 4480
rect 2551 4440 2596 4468
rect 2590 4428 2596 4440
rect 2648 4428 2654 4480
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 2832 4440 4077 4468
rect 2832 4428 2838 4440
rect 4065 4437 4077 4440
rect 4111 4437 4123 4471
rect 4065 4431 4123 4437
rect 1104 4378 6808 4400
rect 1104 4326 2880 4378
rect 2932 4326 2944 4378
rect 2996 4326 3008 4378
rect 3060 4326 3072 4378
rect 3124 4326 3136 4378
rect 3188 4326 4811 4378
rect 4863 4326 4875 4378
rect 4927 4326 4939 4378
rect 4991 4326 5003 4378
rect 5055 4326 5067 4378
rect 5119 4326 6808 4378
rect 1104 4304 6808 4326
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 4249 4131 4307 4137
rect 2179 4100 4108 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 1412 4060 1440 4091
rect 1412 4032 2452 4060
rect 1394 3952 1400 4004
rect 1452 3992 1458 4004
rect 2317 3995 2375 4001
rect 2317 3992 2329 3995
rect 1452 3964 2329 3992
rect 1452 3952 1458 3964
rect 2317 3961 2329 3964
rect 2363 3961 2375 3995
rect 2317 3955 2375 3961
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2424 3924 2452 4032
rect 4080 4001 4108 4100
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4522 4128 4528 4140
rect 4295 4100 4528 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4128 4951 4131
rect 4982 4128 4988 4140
rect 4939 4100 4988 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 5859 4100 6929 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 4065 3995 4123 4001
rect 4065 3961 4077 3995
rect 4111 3961 4123 3995
rect 4065 3955 4123 3961
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 2424 3896 4721 3924
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 5626 3924 5632 3936
rect 5587 3896 5632 3924
rect 4709 3887 4767 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 1104 3834 6808 3856
rect 1104 3782 1915 3834
rect 1967 3782 1979 3834
rect 2031 3782 2043 3834
rect 2095 3782 2107 3834
rect 2159 3782 2171 3834
rect 2223 3782 3846 3834
rect 3898 3782 3910 3834
rect 3962 3782 3974 3834
rect 4026 3782 4038 3834
rect 4090 3782 4102 3834
rect 4154 3782 5776 3834
rect 5828 3782 5840 3834
rect 5892 3782 5904 3834
rect 5956 3782 5968 3834
rect 6020 3782 6032 3834
rect 6084 3782 6808 3834
rect 1104 3760 6808 3782
rect 4338 3720 4344 3732
rect 4299 3692 4344 3720
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 4982 3720 4988 3732
rect 4943 3692 4988 3720
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3516 1455 3519
rect 2774 3516 2780 3528
rect 1443 3488 2780 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5258 3516 5264 3528
rect 5215 3488 5264 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5684 3488 5825 3516
rect 5684 3476 5690 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 1452 3352 1593 3380
rect 1452 3340 1458 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 5994 3380 6000 3392
rect 5955 3352 6000 3380
rect 1581 3343 1639 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 1104 3290 6808 3312
rect 1104 3238 2880 3290
rect 2932 3238 2944 3290
rect 2996 3238 3008 3290
rect 3060 3238 3072 3290
rect 3124 3238 3136 3290
rect 3188 3238 4811 3290
rect 4863 3238 4875 3290
rect 4927 3238 4939 3290
rect 4991 3238 5003 3290
rect 5055 3238 5067 3290
rect 5119 3238 6808 3290
rect 1104 3216 6808 3238
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4985 3179 5043 3185
rect 4985 3176 4997 3179
rect 4488 3148 4997 3176
rect 4488 3136 4494 3148
rect 4985 3145 4997 3148
rect 5031 3145 5043 3179
rect 4985 3139 5043 3145
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5592 3148 5641 3176
rect 5592 3136 5598 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 5629 3139 5687 3145
rect 3605 3111 3663 3117
rect 3605 3077 3617 3111
rect 3651 3108 3663 3111
rect 4614 3108 4620 3120
rect 3651 3080 4620 3108
rect 3651 3077 3663 3080
rect 3605 3071 3663 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 2590 3040 2596 3052
rect 1443 3012 2596 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3040 3479 3043
rect 4706 3040 4712 3052
rect 3467 3012 4712 3040
rect 3467 3009 3479 3012
rect 3421 3003 3479 3009
rect 4706 3000 4712 3012
rect 4764 3000 4770 3052
rect 5166 3040 5172 3052
rect 5127 3012 5172 3040
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6178 3040 6184 3052
rect 5859 3012 6184 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1544 2808 1593 2836
rect 1544 2796 1550 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 1104 2746 6808 2768
rect 1104 2694 1915 2746
rect 1967 2694 1979 2746
rect 2031 2694 2043 2746
rect 2095 2694 2107 2746
rect 2159 2694 2171 2746
rect 2223 2694 3846 2746
rect 3898 2694 3910 2746
rect 3962 2694 3974 2746
rect 4026 2694 4038 2746
rect 4090 2694 4102 2746
rect 4154 2694 5776 2746
rect 5828 2694 5840 2746
rect 5892 2694 5904 2746
rect 5956 2694 5968 2746
rect 6020 2694 6032 2746
rect 6084 2694 6808 2746
rect 1104 2672 6808 2694
rect 4985 2635 5043 2641
rect 4985 2601 4997 2635
rect 5031 2632 5043 2635
rect 5442 2632 5448 2644
rect 5031 2604 5448 2632
rect 5031 2601 5043 2604
rect 4985 2595 5043 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 5350 2524 5356 2576
rect 5408 2564 5414 2576
rect 5629 2567 5687 2573
rect 5629 2564 5641 2567
rect 5408 2536 5641 2564
rect 5408 2524 5414 2536
rect 5629 2533 5641 2536
rect 5675 2533 5687 2567
rect 5629 2527 5687 2533
rect 5258 2496 5264 2508
rect 1412 2468 5264 2496
rect 1412 2437 1440 2468
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 2314 2428 2320 2440
rect 2275 2400 2320 2428
rect 1397 2391 1455 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 2133 2295 2191 2301
rect 2133 2261 2145 2295
rect 2179 2292 2191 2295
rect 2774 2292 2780 2304
rect 2179 2264 2780 2292
rect 2179 2261 2191 2264
rect 2133 2255 2191 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 1104 2202 6808 2224
rect 1104 2150 2880 2202
rect 2932 2150 2944 2202
rect 2996 2150 3008 2202
rect 3060 2150 3072 2202
rect 3124 2150 3136 2202
rect 3188 2150 4811 2202
rect 4863 2150 4875 2202
rect 4927 2150 4939 2202
rect 4991 2150 5003 2202
rect 5055 2150 5067 2202
rect 5119 2150 6808 2202
rect 1104 2128 6808 2150
<< via1 >>
rect 2880 57638 2932 57690
rect 2944 57638 2996 57690
rect 3008 57638 3060 57690
rect 3072 57638 3124 57690
rect 3136 57638 3188 57690
rect 4811 57638 4863 57690
rect 4875 57638 4927 57690
rect 4939 57638 4991 57690
rect 5003 57638 5055 57690
rect 5067 57638 5119 57690
rect 2780 57536 2832 57588
rect 3240 57536 3292 57588
rect 4252 57579 4304 57588
rect 4252 57545 4261 57579
rect 4261 57545 4295 57579
rect 4295 57545 4304 57579
rect 4252 57536 4304 57545
rect 5448 57536 5500 57588
rect 2780 57400 2832 57452
rect 4252 57400 4304 57452
rect 5540 57443 5592 57452
rect 3240 57332 3292 57384
rect 3424 57332 3476 57384
rect 5540 57409 5549 57443
rect 5549 57409 5583 57443
rect 5583 57409 5592 57443
rect 5540 57400 5592 57409
rect 4712 57264 4764 57316
rect 1584 57239 1636 57248
rect 1584 57205 1593 57239
rect 1593 57205 1627 57239
rect 1627 57205 1636 57239
rect 1584 57196 1636 57205
rect 6184 57196 6236 57248
rect 1915 57094 1967 57146
rect 1979 57094 2031 57146
rect 2043 57094 2095 57146
rect 2107 57094 2159 57146
rect 2171 57094 2223 57146
rect 3846 57094 3898 57146
rect 3910 57094 3962 57146
rect 3974 57094 4026 57146
rect 4038 57094 4090 57146
rect 4102 57094 4154 57146
rect 5776 57094 5828 57146
rect 5840 57094 5892 57146
rect 5904 57094 5956 57146
rect 5968 57094 6020 57146
rect 6032 57094 6084 57146
rect 4528 57035 4580 57044
rect 4528 57001 4537 57035
rect 4537 57001 4571 57035
rect 4571 57001 4580 57035
rect 4528 56992 4580 57001
rect 5264 57035 5316 57044
rect 5264 57001 5273 57035
rect 5273 57001 5307 57035
rect 5307 57001 5316 57035
rect 5264 56992 5316 57001
rect 6276 56992 6328 57044
rect 1400 56831 1452 56840
rect 1400 56797 1409 56831
rect 1409 56797 1443 56831
rect 1443 56797 1452 56831
rect 1400 56788 1452 56797
rect 4344 56831 4396 56840
rect 4344 56797 4353 56831
rect 4353 56797 4387 56831
rect 4387 56797 4396 56831
rect 4344 56788 4396 56797
rect 4528 56788 4580 56840
rect 5632 56788 5684 56840
rect 1584 56695 1636 56704
rect 1584 56661 1593 56695
rect 1593 56661 1627 56695
rect 1627 56661 1636 56695
rect 1584 56652 1636 56661
rect 2880 56550 2932 56602
rect 2944 56550 2996 56602
rect 3008 56550 3060 56602
rect 3072 56550 3124 56602
rect 3136 56550 3188 56602
rect 4811 56550 4863 56602
rect 4875 56550 4927 56602
rect 4939 56550 4991 56602
rect 5003 56550 5055 56602
rect 5067 56550 5119 56602
rect 3332 56448 3384 56500
rect 3332 56312 3384 56364
rect 5724 56219 5776 56228
rect 5724 56185 5733 56219
rect 5733 56185 5767 56219
rect 5767 56185 5776 56219
rect 5724 56176 5776 56185
rect 1915 56006 1967 56058
rect 1979 56006 2031 56058
rect 2043 56006 2095 56058
rect 2107 56006 2159 56058
rect 2171 56006 2223 56058
rect 3846 56006 3898 56058
rect 3910 56006 3962 56058
rect 3974 56006 4026 56058
rect 4038 56006 4090 56058
rect 4102 56006 4154 56058
rect 5776 56006 5828 56058
rect 5840 56006 5892 56058
rect 5904 56006 5956 56058
rect 5968 56006 6020 56058
rect 6032 56006 6084 56058
rect 4252 55947 4304 55956
rect 4252 55913 4261 55947
rect 4261 55913 4295 55947
rect 4295 55913 4304 55947
rect 4252 55904 4304 55913
rect 1676 55700 1728 55752
rect 4436 55743 4488 55752
rect 4436 55709 4445 55743
rect 4445 55709 4479 55743
rect 4479 55709 4488 55743
rect 4436 55700 4488 55709
rect 4068 55632 4120 55684
rect 1584 55607 1636 55616
rect 1584 55573 1593 55607
rect 1593 55573 1627 55607
rect 1627 55573 1636 55607
rect 1584 55564 1636 55573
rect 6000 55607 6052 55616
rect 6000 55573 6009 55607
rect 6009 55573 6043 55607
rect 6043 55573 6052 55607
rect 6000 55564 6052 55573
rect 2880 55462 2932 55514
rect 2944 55462 2996 55514
rect 3008 55462 3060 55514
rect 3072 55462 3124 55514
rect 3136 55462 3188 55514
rect 4811 55462 4863 55514
rect 4875 55462 4927 55514
rect 4939 55462 4991 55514
rect 5003 55462 5055 55514
rect 5067 55462 5119 55514
rect 2780 55360 2832 55412
rect 3240 55360 3292 55412
rect 5540 55360 5592 55412
rect 5632 55292 5684 55344
rect 1492 55224 1544 55276
rect 2412 55224 2464 55276
rect 4068 55224 4120 55276
rect 4252 55267 4304 55276
rect 4252 55233 4261 55267
rect 4261 55233 4295 55267
rect 4295 55233 4304 55267
rect 4252 55224 4304 55233
rect 4252 55088 4304 55140
rect 5356 55267 5408 55276
rect 5356 55233 5365 55267
rect 5365 55233 5399 55267
rect 5399 55233 5408 55267
rect 5356 55224 5408 55233
rect 5724 55131 5776 55140
rect 5724 55097 5733 55131
rect 5733 55097 5767 55131
rect 5767 55097 5776 55131
rect 5724 55088 5776 55097
rect 1584 55063 1636 55072
rect 1584 55029 1593 55063
rect 1593 55029 1627 55063
rect 1627 55029 1636 55063
rect 1584 55020 1636 55029
rect 1915 54918 1967 54970
rect 1979 54918 2031 54970
rect 2043 54918 2095 54970
rect 2107 54918 2159 54970
rect 2171 54918 2223 54970
rect 3846 54918 3898 54970
rect 3910 54918 3962 54970
rect 3974 54918 4026 54970
rect 4038 54918 4090 54970
rect 4102 54918 4154 54970
rect 5776 54918 5828 54970
rect 5840 54918 5892 54970
rect 5904 54918 5956 54970
rect 5968 54918 6020 54970
rect 6032 54918 6084 54970
rect 3424 54816 3476 54868
rect 4528 54816 4580 54868
rect 1768 54612 1820 54664
rect 3516 54612 3568 54664
rect 2780 54544 2832 54596
rect 1584 54519 1636 54528
rect 1584 54485 1593 54519
rect 1593 54485 1627 54519
rect 1627 54485 1636 54519
rect 1584 54476 1636 54485
rect 4620 54476 4672 54528
rect 5356 54476 5408 54528
rect 6000 54519 6052 54528
rect 6000 54485 6009 54519
rect 6009 54485 6043 54519
rect 6043 54485 6052 54519
rect 6000 54476 6052 54485
rect 2880 54374 2932 54426
rect 2944 54374 2996 54426
rect 3008 54374 3060 54426
rect 3072 54374 3124 54426
rect 3136 54374 3188 54426
rect 4811 54374 4863 54426
rect 4875 54374 4927 54426
rect 4939 54374 4991 54426
rect 5003 54374 5055 54426
rect 5067 54374 5119 54426
rect 3332 54272 3384 54324
rect 4344 54272 4396 54324
rect 5356 54136 5408 54188
rect 4528 54068 4580 54120
rect 5724 54043 5776 54052
rect 5724 54009 5733 54043
rect 5733 54009 5767 54043
rect 5767 54009 5776 54043
rect 5724 54000 5776 54009
rect 1915 53830 1967 53882
rect 1979 53830 2031 53882
rect 2043 53830 2095 53882
rect 2107 53830 2159 53882
rect 2171 53830 2223 53882
rect 3846 53830 3898 53882
rect 3910 53830 3962 53882
rect 3974 53830 4026 53882
rect 4038 53830 4090 53882
rect 4102 53830 4154 53882
rect 5776 53830 5828 53882
rect 5840 53830 5892 53882
rect 5904 53830 5956 53882
rect 5968 53830 6020 53882
rect 6032 53830 6084 53882
rect 3424 53524 3476 53576
rect 1584 53431 1636 53440
rect 1584 53397 1593 53431
rect 1593 53397 1627 53431
rect 1627 53397 1636 53431
rect 1584 53388 1636 53397
rect 6000 53431 6052 53440
rect 6000 53397 6009 53431
rect 6009 53397 6043 53431
rect 6043 53397 6052 53431
rect 6000 53388 6052 53397
rect 2880 53286 2932 53338
rect 2944 53286 2996 53338
rect 3008 53286 3060 53338
rect 3072 53286 3124 53338
rect 3136 53286 3188 53338
rect 4811 53286 4863 53338
rect 4875 53286 4927 53338
rect 4939 53286 4991 53338
rect 5003 53286 5055 53338
rect 5067 53286 5119 53338
rect 3424 53227 3476 53236
rect 3424 53193 3433 53227
rect 3433 53193 3467 53227
rect 3467 53193 3476 53227
rect 3424 53184 3476 53193
rect 2872 53048 2924 53100
rect 1584 52887 1636 52896
rect 1584 52853 1593 52887
rect 1593 52853 1627 52887
rect 1627 52853 1636 52887
rect 1584 52844 1636 52853
rect 5264 52844 5316 52896
rect 6184 52844 6236 52896
rect 1915 52742 1967 52794
rect 1979 52742 2031 52794
rect 2043 52742 2095 52794
rect 2107 52742 2159 52794
rect 2171 52742 2223 52794
rect 3846 52742 3898 52794
rect 3910 52742 3962 52794
rect 3974 52742 4026 52794
rect 4038 52742 4090 52794
rect 4102 52742 4154 52794
rect 5776 52742 5828 52794
rect 5840 52742 5892 52794
rect 5904 52742 5956 52794
rect 5968 52742 6020 52794
rect 6032 52742 6084 52794
rect 2780 52640 2832 52692
rect 3240 52479 3292 52488
rect 3240 52445 3249 52479
rect 3249 52445 3283 52479
rect 3283 52445 3292 52479
rect 3240 52436 3292 52445
rect 6460 52436 6512 52488
rect 6000 52343 6052 52352
rect 6000 52309 6009 52343
rect 6009 52309 6043 52343
rect 6043 52309 6052 52343
rect 6000 52300 6052 52309
rect 2880 52198 2932 52250
rect 2944 52198 2996 52250
rect 3008 52198 3060 52250
rect 3072 52198 3124 52250
rect 3136 52198 3188 52250
rect 4811 52198 4863 52250
rect 4875 52198 4927 52250
rect 4939 52198 4991 52250
rect 5003 52198 5055 52250
rect 5067 52198 5119 52250
rect 1676 51960 1728 52012
rect 3700 52003 3752 52012
rect 3700 51969 3709 52003
rect 3709 51969 3743 52003
rect 3743 51969 3752 52003
rect 3700 51960 3752 51969
rect 1584 51867 1636 51876
rect 1584 51833 1593 51867
rect 1593 51833 1627 51867
rect 1627 51833 1636 51867
rect 1584 51824 1636 51833
rect 6184 51756 6236 51808
rect 1915 51654 1967 51706
rect 1979 51654 2031 51706
rect 2043 51654 2095 51706
rect 2107 51654 2159 51706
rect 2171 51654 2223 51706
rect 3846 51654 3898 51706
rect 3910 51654 3962 51706
rect 3974 51654 4026 51706
rect 4038 51654 4090 51706
rect 4102 51654 4154 51706
rect 5776 51654 5828 51706
rect 5840 51654 5892 51706
rect 5904 51654 5956 51706
rect 5968 51654 6020 51706
rect 6032 51654 6084 51706
rect 1400 51391 1452 51400
rect 1400 51357 1409 51391
rect 1409 51357 1443 51391
rect 1443 51357 1452 51391
rect 1400 51348 1452 51357
rect 1584 51255 1636 51264
rect 1584 51221 1593 51255
rect 1593 51221 1627 51255
rect 1627 51221 1636 51255
rect 1584 51212 1636 51221
rect 6000 51255 6052 51264
rect 6000 51221 6009 51255
rect 6009 51221 6043 51255
rect 6043 51221 6052 51255
rect 6000 51212 6052 51221
rect 2880 51110 2932 51162
rect 2944 51110 2996 51162
rect 3008 51110 3060 51162
rect 3072 51110 3124 51162
rect 3136 51110 3188 51162
rect 4811 51110 4863 51162
rect 4875 51110 4927 51162
rect 4939 51110 4991 51162
rect 5003 51110 5055 51162
rect 5067 51110 5119 51162
rect 1400 51008 1452 51060
rect 2780 51051 2832 51060
rect 2780 51017 2789 51051
rect 2789 51017 2823 51051
rect 2823 51017 2832 51051
rect 2780 51008 2832 51017
rect 1400 50915 1452 50924
rect 1400 50881 1409 50915
rect 1409 50881 1443 50915
rect 1443 50881 1452 50915
rect 1400 50872 1452 50881
rect 2320 50915 2372 50924
rect 2320 50881 2329 50915
rect 2329 50881 2363 50915
rect 2363 50881 2372 50915
rect 2320 50872 2372 50881
rect 2780 50872 2832 50924
rect 1584 50711 1636 50720
rect 1584 50677 1593 50711
rect 1593 50677 1627 50711
rect 1627 50677 1636 50711
rect 1584 50668 1636 50677
rect 6368 50668 6420 50720
rect 1915 50566 1967 50618
rect 1979 50566 2031 50618
rect 2043 50566 2095 50618
rect 2107 50566 2159 50618
rect 2171 50566 2223 50618
rect 3846 50566 3898 50618
rect 3910 50566 3962 50618
rect 3974 50566 4026 50618
rect 4038 50566 4090 50618
rect 4102 50566 4154 50618
rect 5776 50566 5828 50618
rect 5840 50566 5892 50618
rect 5904 50566 5956 50618
rect 5968 50566 6020 50618
rect 6032 50566 6084 50618
rect 1400 50464 1452 50516
rect 5540 50260 5592 50312
rect 6000 50167 6052 50176
rect 6000 50133 6009 50167
rect 6009 50133 6043 50167
rect 6043 50133 6052 50167
rect 6000 50124 6052 50133
rect 2880 50022 2932 50074
rect 2944 50022 2996 50074
rect 3008 50022 3060 50074
rect 3072 50022 3124 50074
rect 3136 50022 3188 50074
rect 4811 50022 4863 50074
rect 4875 50022 4927 50074
rect 4939 50022 4991 50074
rect 5003 50022 5055 50074
rect 5067 50022 5119 50074
rect 1676 49920 1728 49972
rect 3424 49716 3476 49768
rect 4712 49716 4764 49768
rect 1584 49623 1636 49632
rect 1584 49589 1593 49623
rect 1593 49589 1627 49623
rect 1627 49589 1636 49623
rect 1584 49580 1636 49589
rect 6184 49580 6236 49632
rect 1915 49478 1967 49530
rect 1979 49478 2031 49530
rect 2043 49478 2095 49530
rect 2107 49478 2159 49530
rect 2171 49478 2223 49530
rect 3846 49478 3898 49530
rect 3910 49478 3962 49530
rect 3974 49478 4026 49530
rect 4038 49478 4090 49530
rect 4102 49478 4154 49530
rect 5776 49478 5828 49530
rect 5840 49478 5892 49530
rect 5904 49478 5956 49530
rect 5968 49478 6020 49530
rect 6032 49478 6084 49530
rect 3332 49172 3384 49224
rect 4344 49172 4396 49224
rect 1584 49079 1636 49088
rect 1584 49045 1593 49079
rect 1593 49045 1627 49079
rect 1627 49045 1636 49079
rect 1584 49036 1636 49045
rect 6000 49079 6052 49088
rect 6000 49045 6009 49079
rect 6009 49045 6043 49079
rect 6043 49045 6052 49079
rect 6000 49036 6052 49045
rect 2880 48934 2932 48986
rect 2944 48934 2996 48986
rect 3008 48934 3060 48986
rect 3072 48934 3124 48986
rect 3136 48934 3188 48986
rect 4811 48934 4863 48986
rect 4875 48934 4927 48986
rect 4939 48934 4991 48986
rect 5003 48934 5055 48986
rect 5067 48934 5119 48986
rect 4620 48764 4672 48816
rect 5356 48764 5408 48816
rect 4620 48492 4672 48544
rect 6184 48492 6236 48544
rect 1915 48390 1967 48442
rect 1979 48390 2031 48442
rect 2043 48390 2095 48442
rect 2107 48390 2159 48442
rect 2171 48390 2223 48442
rect 3846 48390 3898 48442
rect 3910 48390 3962 48442
rect 3974 48390 4026 48442
rect 4038 48390 4090 48442
rect 4102 48390 4154 48442
rect 5776 48390 5828 48442
rect 5840 48390 5892 48442
rect 5904 48390 5956 48442
rect 5968 48390 6020 48442
rect 6032 48390 6084 48442
rect 4804 48288 4856 48340
rect 5540 48288 5592 48340
rect 2872 48084 2924 48136
rect 3516 48084 3568 48136
rect 6644 48084 6696 48136
rect 1584 47991 1636 48000
rect 1584 47957 1593 47991
rect 1593 47957 1627 47991
rect 1627 47957 1636 47991
rect 1584 47948 1636 47957
rect 3424 47948 3476 48000
rect 6000 47991 6052 48000
rect 6000 47957 6009 47991
rect 6009 47957 6043 47991
rect 6043 47957 6052 47991
rect 6000 47948 6052 47957
rect 2880 47846 2932 47898
rect 2944 47846 2996 47898
rect 3008 47846 3060 47898
rect 3072 47846 3124 47898
rect 3136 47846 3188 47898
rect 4811 47846 4863 47898
rect 4875 47846 4927 47898
rect 4939 47846 4991 47898
rect 5003 47846 5055 47898
rect 5067 47846 5119 47898
rect 4344 47608 4396 47660
rect 6552 47472 6604 47524
rect 1584 47447 1636 47456
rect 1584 47413 1593 47447
rect 1593 47413 1627 47447
rect 1627 47413 1636 47447
rect 1584 47404 1636 47413
rect 6184 47404 6236 47456
rect 1915 47302 1967 47354
rect 1979 47302 2031 47354
rect 2043 47302 2095 47354
rect 2107 47302 2159 47354
rect 2171 47302 2223 47354
rect 3846 47302 3898 47354
rect 3910 47302 3962 47354
rect 3974 47302 4026 47354
rect 4038 47302 4090 47354
rect 4102 47302 4154 47354
rect 5776 47302 5828 47354
rect 5840 47302 5892 47354
rect 5904 47302 5956 47354
rect 5968 47302 6020 47354
rect 6032 47302 6084 47354
rect 1400 47039 1452 47048
rect 1400 47005 1409 47039
rect 1409 47005 1443 47039
rect 1443 47005 1452 47039
rect 1400 46996 1452 47005
rect 3424 46996 3476 47048
rect 1584 46903 1636 46912
rect 1584 46869 1593 46903
rect 1593 46869 1627 46903
rect 1627 46869 1636 46903
rect 1584 46860 1636 46869
rect 6000 46903 6052 46912
rect 6000 46869 6009 46903
rect 6009 46869 6043 46903
rect 6043 46869 6052 46903
rect 6000 46860 6052 46869
rect 2880 46758 2932 46810
rect 2944 46758 2996 46810
rect 3008 46758 3060 46810
rect 3072 46758 3124 46810
rect 3136 46758 3188 46810
rect 4811 46758 4863 46810
rect 4875 46758 4927 46810
rect 4939 46758 4991 46810
rect 5003 46758 5055 46810
rect 5067 46758 5119 46810
rect 7748 46767 7800 46776
rect 7748 46733 7757 46767
rect 7757 46733 7791 46767
rect 7791 46733 7800 46767
rect 7748 46724 7800 46733
rect 3332 46656 3384 46708
rect 4344 46656 4396 46708
rect 6276 46520 6328 46572
rect 5080 46316 5132 46368
rect 5264 46316 5316 46368
rect 6184 46316 6236 46368
rect 1915 46214 1967 46266
rect 1979 46214 2031 46266
rect 2043 46214 2095 46266
rect 2107 46214 2159 46266
rect 2171 46214 2223 46266
rect 3846 46214 3898 46266
rect 3910 46214 3962 46266
rect 3974 46214 4026 46266
rect 4038 46214 4090 46266
rect 4102 46214 4154 46266
rect 5776 46214 5828 46266
rect 5840 46214 5892 46266
rect 5904 46214 5956 46266
rect 5968 46214 6020 46266
rect 6032 46214 6084 46266
rect 4252 46044 4304 46096
rect 4712 46044 4764 46096
rect 5356 46112 5408 46164
rect 3240 45976 3292 46028
rect 5264 45976 5316 46028
rect 2688 45908 2740 45960
rect 5816 45951 5868 45960
rect 5816 45917 5825 45951
rect 5825 45917 5859 45951
rect 5859 45917 5868 45951
rect 5816 45908 5868 45917
rect 5080 45840 5132 45892
rect 1584 45815 1636 45824
rect 1584 45781 1593 45815
rect 1593 45781 1627 45815
rect 1627 45781 1636 45815
rect 1584 45772 1636 45781
rect 3240 45772 3292 45824
rect 5356 45772 5408 45824
rect 6000 45815 6052 45824
rect 6000 45781 6009 45815
rect 6009 45781 6043 45815
rect 6043 45781 6052 45815
rect 6000 45772 6052 45781
rect 2880 45670 2932 45722
rect 2944 45670 2996 45722
rect 3008 45670 3060 45722
rect 3072 45670 3124 45722
rect 3136 45670 3188 45722
rect 4811 45670 4863 45722
rect 4875 45670 4927 45722
rect 4939 45670 4991 45722
rect 5003 45670 5055 45722
rect 5067 45670 5119 45722
rect 1492 45432 1544 45484
rect 1584 45271 1636 45280
rect 1584 45237 1593 45271
rect 1593 45237 1627 45271
rect 1627 45237 1636 45271
rect 1584 45228 1636 45237
rect 4712 45228 4764 45280
rect 6184 45228 6236 45280
rect 1915 45126 1967 45178
rect 1979 45126 2031 45178
rect 2043 45126 2095 45178
rect 2107 45126 2159 45178
rect 2171 45126 2223 45178
rect 3846 45126 3898 45178
rect 3910 45126 3962 45178
rect 3974 45126 4026 45178
rect 4038 45126 4090 45178
rect 4102 45126 4154 45178
rect 5776 45126 5828 45178
rect 5840 45126 5892 45178
rect 5904 45126 5956 45178
rect 5968 45126 6020 45178
rect 6032 45126 6084 45178
rect 1400 45024 1452 45076
rect 2412 44820 2464 44872
rect 6828 44820 6880 44872
rect 6000 44727 6052 44736
rect 6000 44693 6009 44727
rect 6009 44693 6043 44727
rect 6043 44693 6052 44727
rect 6000 44684 6052 44693
rect 2880 44582 2932 44634
rect 2944 44582 2996 44634
rect 3008 44582 3060 44634
rect 3072 44582 3124 44634
rect 3136 44582 3188 44634
rect 4811 44582 4863 44634
rect 4875 44582 4927 44634
rect 4939 44582 4991 44634
rect 5003 44582 5055 44634
rect 5067 44582 5119 44634
rect 3148 44344 3200 44396
rect 5540 44387 5592 44396
rect 5540 44353 5549 44387
rect 5549 44353 5583 44387
rect 5583 44353 5592 44387
rect 5540 44344 5592 44353
rect 1584 44251 1636 44260
rect 1584 44217 1593 44251
rect 1593 44217 1627 44251
rect 1627 44217 1636 44251
rect 1584 44208 1636 44217
rect 5632 44140 5684 44192
rect 1915 44038 1967 44090
rect 1979 44038 2031 44090
rect 2043 44038 2095 44090
rect 2107 44038 2159 44090
rect 2171 44038 2223 44090
rect 3846 44038 3898 44090
rect 3910 44038 3962 44090
rect 3974 44038 4026 44090
rect 4038 44038 4090 44090
rect 4102 44038 4154 44090
rect 5776 44038 5828 44090
rect 5840 44038 5892 44090
rect 5904 44038 5956 44090
rect 5968 44038 6020 44090
rect 6032 44038 6084 44090
rect 1216 43868 1268 43920
rect 2504 43868 2556 43920
rect 2504 43732 2556 43784
rect 6276 43732 6328 43784
rect 1584 43639 1636 43648
rect 1584 43605 1593 43639
rect 1593 43605 1627 43639
rect 1627 43605 1636 43639
rect 1584 43596 1636 43605
rect 6000 43639 6052 43648
rect 6000 43605 6009 43639
rect 6009 43605 6043 43639
rect 6043 43605 6052 43639
rect 6000 43596 6052 43605
rect 2880 43494 2932 43546
rect 2944 43494 2996 43546
rect 3008 43494 3060 43546
rect 3072 43494 3124 43546
rect 3136 43494 3188 43546
rect 4811 43494 4863 43546
rect 4875 43494 4927 43546
rect 4939 43494 4991 43546
rect 5003 43494 5055 43546
rect 5067 43494 5119 43546
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 6368 43256 6420 43308
rect 1584 43095 1636 43104
rect 1584 43061 1593 43095
rect 1593 43061 1627 43095
rect 1627 43061 1636 43095
rect 1584 43052 1636 43061
rect 5632 43052 5684 43104
rect 1915 42950 1967 43002
rect 1979 42950 2031 43002
rect 2043 42950 2095 43002
rect 2107 42950 2159 43002
rect 2171 42950 2223 43002
rect 3846 42950 3898 43002
rect 3910 42950 3962 43002
rect 3974 42950 4026 43002
rect 4038 42950 4090 43002
rect 4102 42950 4154 43002
rect 5776 42950 5828 43002
rect 5840 42950 5892 43002
rect 5904 42950 5956 43002
rect 5968 42950 6020 43002
rect 6032 42950 6084 43002
rect 2880 42406 2932 42458
rect 2944 42406 2996 42458
rect 3008 42406 3060 42458
rect 3072 42406 3124 42458
rect 3136 42406 3188 42458
rect 4811 42406 4863 42458
rect 4875 42406 4927 42458
rect 4939 42406 4991 42458
rect 5003 42406 5055 42458
rect 5067 42406 5119 42458
rect 1400 42304 1452 42356
rect 5448 42304 5500 42356
rect 5080 42236 5132 42288
rect 7472 42279 7524 42288
rect 7472 42245 7481 42279
rect 7481 42245 7515 42279
rect 7515 42245 7524 42279
rect 7472 42236 7524 42245
rect 5448 42168 5500 42220
rect 1584 42075 1636 42084
rect 1584 42041 1593 42075
rect 1593 42041 1627 42075
rect 1627 42041 1636 42075
rect 1584 42032 1636 42041
rect 5724 42075 5776 42084
rect 5724 42041 5733 42075
rect 5733 42041 5767 42075
rect 5767 42041 5776 42075
rect 5724 42032 5776 42041
rect 5448 42007 5500 42016
rect 5448 41973 5457 42007
rect 5457 41973 5491 42007
rect 5491 41973 5500 42007
rect 5448 41964 5500 41973
rect 1915 41862 1967 41914
rect 1979 41862 2031 41914
rect 2043 41862 2095 41914
rect 2107 41862 2159 41914
rect 2171 41862 2223 41914
rect 3846 41862 3898 41914
rect 3910 41862 3962 41914
rect 3974 41862 4026 41914
rect 4038 41862 4090 41914
rect 4102 41862 4154 41914
rect 5776 41862 5828 41914
rect 5840 41862 5892 41914
rect 5904 41862 5956 41914
rect 5968 41862 6020 41914
rect 6032 41862 6084 41914
rect 5172 41760 5224 41812
rect 4252 41624 4304 41676
rect 4528 41624 4580 41676
rect 2228 41556 2280 41608
rect 3332 41556 3384 41608
rect 5264 41599 5316 41608
rect 5264 41565 5273 41599
rect 5273 41565 5307 41599
rect 5307 41565 5316 41599
rect 5264 41556 5316 41565
rect 1308 41488 1360 41540
rect 1676 41488 1728 41540
rect 1584 41463 1636 41472
rect 1584 41429 1593 41463
rect 1593 41429 1627 41463
rect 1627 41429 1636 41463
rect 1584 41420 1636 41429
rect 7656 41488 7708 41540
rect 5540 41420 5592 41472
rect 7472 41417 7524 41426
rect 7472 41383 7481 41417
rect 7481 41383 7515 41417
rect 7515 41383 7524 41417
rect 7472 41374 7524 41383
rect 7932 41395 7984 41404
rect 2880 41318 2932 41370
rect 2944 41318 2996 41370
rect 3008 41318 3060 41370
rect 3072 41318 3124 41370
rect 3136 41318 3188 41370
rect 4811 41318 4863 41370
rect 4875 41318 4927 41370
rect 4939 41318 4991 41370
rect 5003 41318 5055 41370
rect 5067 41318 5119 41370
rect 7932 41361 7941 41395
rect 7941 41361 7975 41395
rect 7975 41361 7984 41395
rect 7932 41352 7984 41361
rect 3240 41216 3292 41268
rect 3424 41216 3476 41268
rect 7656 41148 7708 41200
rect 1124 41080 1176 41132
rect 2412 41080 2464 41132
rect 2596 41080 2648 41132
rect 4988 41055 5040 41064
rect 4988 41021 4997 41055
rect 4997 41021 5031 41055
rect 5031 41021 5040 41055
rect 4988 41012 5040 41021
rect 5172 41012 5224 41064
rect 6552 41012 6604 41064
rect 2228 40944 2280 40996
rect 2412 40944 2464 40996
rect 2596 40944 2648 40996
rect 1584 40919 1636 40928
rect 1584 40885 1593 40919
rect 1593 40885 1627 40919
rect 1627 40885 1636 40919
rect 1584 40876 1636 40885
rect 1915 40774 1967 40826
rect 1979 40774 2031 40826
rect 2043 40774 2095 40826
rect 2107 40774 2159 40826
rect 2171 40774 2223 40826
rect 3846 40774 3898 40826
rect 3910 40774 3962 40826
rect 3974 40774 4026 40826
rect 4038 40774 4090 40826
rect 4102 40774 4154 40826
rect 5776 40774 5828 40826
rect 5840 40774 5892 40826
rect 5904 40774 5956 40826
rect 5968 40774 6020 40826
rect 6032 40774 6084 40826
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 5724 40468 5776 40520
rect 7748 40400 7800 40452
rect 1584 40375 1636 40384
rect 1584 40341 1593 40375
rect 1593 40341 1627 40375
rect 1627 40341 1636 40375
rect 1584 40332 1636 40341
rect 2880 40230 2932 40282
rect 2944 40230 2996 40282
rect 3008 40230 3060 40282
rect 3072 40230 3124 40282
rect 3136 40230 3188 40282
rect 4811 40230 4863 40282
rect 4875 40230 4927 40282
rect 4939 40230 4991 40282
rect 5003 40230 5055 40282
rect 5067 40230 5119 40282
rect 5540 40128 5592 40180
rect 1676 39992 1728 40044
rect 5816 40035 5868 40044
rect 5816 40001 5825 40035
rect 5825 40001 5859 40035
rect 5859 40001 5868 40035
rect 5816 39992 5868 40001
rect 5632 39924 5684 39976
rect 1216 39856 1268 39908
rect 1676 39856 1728 39908
rect 1915 39686 1967 39738
rect 1979 39686 2031 39738
rect 2043 39686 2095 39738
rect 2107 39686 2159 39738
rect 2171 39686 2223 39738
rect 3846 39686 3898 39738
rect 3910 39686 3962 39738
rect 3974 39686 4026 39738
rect 4038 39686 4090 39738
rect 4102 39686 4154 39738
rect 5776 39686 5828 39738
rect 5840 39686 5892 39738
rect 5904 39686 5956 39738
rect 5968 39686 6020 39738
rect 6032 39686 6084 39738
rect 5632 39584 5684 39636
rect 1216 39380 1268 39432
rect 6092 39423 6144 39432
rect 6092 39389 6101 39423
rect 6101 39389 6135 39423
rect 6135 39389 6144 39423
rect 6092 39380 6144 39389
rect 1584 39287 1636 39296
rect 1584 39253 1593 39287
rect 1593 39253 1627 39287
rect 1627 39253 1636 39287
rect 1584 39244 1636 39253
rect 2880 39142 2932 39194
rect 2944 39142 2996 39194
rect 3008 39142 3060 39194
rect 3072 39142 3124 39194
rect 3136 39142 3188 39194
rect 4811 39142 4863 39194
rect 4875 39142 4927 39194
rect 4939 39142 4991 39194
rect 5003 39142 5055 39194
rect 5067 39142 5119 39194
rect 1676 38972 1728 39024
rect 6184 39040 6236 39092
rect 6736 39040 6788 39092
rect 6184 38904 6236 38956
rect 1400 38836 1452 38888
rect 1676 38836 1728 38888
rect 1400 38700 1452 38752
rect 2504 38700 2556 38752
rect 1915 38598 1967 38650
rect 1979 38598 2031 38650
rect 2043 38598 2095 38650
rect 2107 38598 2159 38650
rect 2171 38598 2223 38650
rect 3846 38598 3898 38650
rect 3910 38598 3962 38650
rect 3974 38598 4026 38650
rect 4038 38598 4090 38650
rect 4102 38598 4154 38650
rect 5776 38598 5828 38650
rect 5840 38598 5892 38650
rect 5904 38598 5956 38650
rect 5968 38598 6020 38650
rect 6032 38598 6084 38650
rect 3056 38496 3108 38548
rect 3332 38496 3384 38548
rect 3424 38496 3476 38548
rect 1308 38360 1360 38412
rect 3148 38360 3200 38412
rect 3884 38360 3936 38412
rect 2596 38292 2648 38344
rect 2964 38292 3016 38344
rect 3516 38292 3568 38344
rect 6092 38335 6144 38344
rect 6092 38301 6101 38335
rect 6101 38301 6135 38335
rect 6135 38301 6144 38335
rect 6092 38292 6144 38301
rect 3056 38224 3108 38276
rect 3148 38224 3200 38276
rect 1584 38199 1636 38208
rect 1584 38165 1593 38199
rect 1593 38165 1627 38199
rect 1627 38165 1636 38199
rect 1584 38156 1636 38165
rect 3332 38156 3384 38208
rect 2880 38054 2932 38106
rect 2944 38054 2996 38106
rect 3008 38054 3060 38106
rect 3072 38054 3124 38106
rect 3136 38054 3188 38106
rect 4811 38054 4863 38106
rect 4875 38054 4927 38106
rect 4939 38054 4991 38106
rect 5003 38054 5055 38106
rect 5067 38054 5119 38106
rect 1768 37884 1820 37936
rect 2412 37884 2464 37936
rect 2320 37816 2372 37868
rect 3884 37816 3936 37868
rect 4988 37791 5040 37800
rect 4988 37757 4997 37791
rect 4997 37757 5031 37791
rect 5031 37757 5040 37791
rect 4988 37748 5040 37757
rect 1584 37655 1636 37664
rect 1584 37621 1593 37655
rect 1593 37621 1627 37655
rect 1627 37621 1636 37655
rect 1584 37612 1636 37621
rect 1915 37510 1967 37562
rect 1979 37510 2031 37562
rect 2043 37510 2095 37562
rect 2107 37510 2159 37562
rect 2171 37510 2223 37562
rect 3846 37510 3898 37562
rect 3910 37510 3962 37562
rect 3974 37510 4026 37562
rect 4038 37510 4090 37562
rect 4102 37510 4154 37562
rect 5776 37510 5828 37562
rect 5840 37510 5892 37562
rect 5904 37510 5956 37562
rect 5968 37510 6020 37562
rect 6032 37510 6084 37562
rect 5264 37408 5316 37460
rect 3884 37340 3936 37392
rect 5264 37315 5316 37324
rect 5264 37281 5273 37315
rect 5273 37281 5307 37315
rect 5307 37281 5316 37315
rect 5264 37272 5316 37281
rect 2688 37068 2740 37120
rect 2880 36966 2932 37018
rect 2944 36966 2996 37018
rect 3008 36966 3060 37018
rect 3072 36966 3124 37018
rect 3136 36966 3188 37018
rect 4811 36966 4863 37018
rect 4875 36966 4927 37018
rect 4939 36966 4991 37018
rect 5003 36966 5055 37018
rect 5067 36966 5119 37018
rect 1492 36864 1544 36916
rect 1768 36864 1820 36916
rect 1676 36728 1728 36780
rect 2780 36728 2832 36780
rect 2872 36660 2924 36712
rect 3884 36660 3936 36712
rect 4988 36703 5040 36712
rect 4988 36669 4997 36703
rect 4997 36669 5031 36703
rect 5031 36669 5040 36703
rect 4988 36660 5040 36669
rect 1584 36635 1636 36644
rect 1584 36601 1593 36635
rect 1593 36601 1627 36635
rect 1627 36601 1636 36635
rect 1584 36592 1636 36601
rect 2780 36592 2832 36644
rect 3608 36592 3660 36644
rect 4620 36592 4672 36644
rect 4804 36592 4856 36644
rect 1915 36422 1967 36474
rect 1979 36422 2031 36474
rect 2043 36422 2095 36474
rect 2107 36422 2159 36474
rect 2171 36422 2223 36474
rect 3846 36422 3898 36474
rect 3910 36422 3962 36474
rect 3974 36422 4026 36474
rect 4038 36422 4090 36474
rect 4102 36422 4154 36474
rect 5776 36422 5828 36474
rect 5840 36422 5892 36474
rect 5904 36422 5956 36474
rect 5968 36422 6020 36474
rect 6032 36422 6084 36474
rect 7932 36456 7984 36508
rect 5540 36320 5592 36372
rect 6644 36320 6696 36372
rect 1492 36116 1544 36168
rect 5264 36159 5316 36168
rect 5264 36125 5273 36159
rect 5273 36125 5307 36159
rect 5307 36125 5316 36159
rect 5264 36116 5316 36125
rect 2044 36048 2096 36100
rect 2872 36048 2924 36100
rect 1308 35980 1360 36032
rect 2880 35878 2932 35930
rect 2944 35878 2996 35930
rect 3008 35878 3060 35930
rect 3072 35878 3124 35930
rect 3136 35878 3188 35930
rect 4811 35878 4863 35930
rect 4875 35878 4927 35930
rect 4939 35878 4991 35930
rect 5003 35878 5055 35930
rect 5067 35878 5119 35930
rect 3240 35776 3292 35828
rect 2044 35751 2096 35760
rect 2044 35717 2053 35751
rect 2053 35717 2087 35751
rect 2087 35717 2096 35751
rect 2044 35708 2096 35717
rect 1400 35640 1452 35692
rect 5172 35708 5224 35760
rect 2504 35572 2556 35624
rect 4988 35615 5040 35624
rect 4988 35581 4997 35615
rect 4997 35581 5031 35615
rect 5031 35581 5040 35615
rect 4988 35572 5040 35581
rect 1915 35334 1967 35386
rect 1979 35334 2031 35386
rect 2043 35334 2095 35386
rect 2107 35334 2159 35386
rect 2171 35334 2223 35386
rect 3846 35334 3898 35386
rect 3910 35334 3962 35386
rect 3974 35334 4026 35386
rect 4038 35334 4090 35386
rect 4102 35334 4154 35386
rect 5776 35334 5828 35386
rect 5840 35334 5892 35386
rect 5904 35334 5956 35386
rect 5968 35334 6020 35386
rect 6032 35334 6084 35386
rect 5264 35164 5316 35216
rect 5540 35164 5592 35216
rect 5264 35071 5316 35080
rect 5264 35037 5273 35071
rect 5273 35037 5307 35071
rect 5307 35037 5316 35071
rect 5264 35028 5316 35037
rect 2880 34790 2932 34842
rect 2944 34790 2996 34842
rect 3008 34790 3060 34842
rect 3072 34790 3124 34842
rect 3136 34790 3188 34842
rect 4811 34790 4863 34842
rect 4875 34790 4927 34842
rect 4939 34790 4991 34842
rect 5003 34790 5055 34842
rect 5067 34790 5119 34842
rect 2596 34688 2648 34740
rect 4344 34620 4396 34672
rect 1860 34595 1912 34604
rect 1860 34561 1869 34595
rect 1869 34561 1903 34595
rect 1903 34561 1912 34595
rect 1860 34552 1912 34561
rect 1216 34484 1268 34536
rect 2596 34484 2648 34536
rect 3424 34552 3476 34604
rect 4988 34527 5040 34536
rect 4988 34493 4997 34527
rect 4997 34493 5031 34527
rect 5031 34493 5040 34527
rect 4988 34484 5040 34493
rect 1915 34246 1967 34298
rect 1979 34246 2031 34298
rect 2043 34246 2095 34298
rect 2107 34246 2159 34298
rect 2171 34246 2223 34298
rect 3846 34246 3898 34298
rect 3910 34246 3962 34298
rect 3974 34246 4026 34298
rect 4038 34246 4090 34298
rect 4102 34246 4154 34298
rect 5776 34246 5828 34298
rect 5840 34246 5892 34298
rect 5904 34246 5956 34298
rect 5968 34246 6020 34298
rect 6032 34246 6084 34298
rect 2688 34144 2740 34196
rect 1400 34076 1452 34128
rect 2780 34008 2832 34060
rect 5264 33983 5316 33992
rect 1860 33915 1912 33924
rect 1860 33881 1869 33915
rect 1869 33881 1903 33915
rect 1903 33881 1912 33915
rect 1860 33872 1912 33881
rect 5264 33949 5273 33983
rect 5273 33949 5307 33983
rect 5307 33949 5316 33983
rect 5264 33940 5316 33949
rect 2880 33702 2932 33754
rect 2944 33702 2996 33754
rect 3008 33702 3060 33754
rect 3072 33702 3124 33754
rect 3136 33702 3188 33754
rect 4811 33702 4863 33754
rect 4875 33702 4927 33754
rect 4939 33702 4991 33754
rect 5003 33702 5055 33754
rect 5067 33702 5119 33754
rect 2688 33600 2740 33652
rect 5356 33600 5408 33652
rect 2412 33532 2464 33584
rect 1400 33464 1452 33516
rect 3516 33464 3568 33516
rect 1124 33396 1176 33448
rect 2412 33396 2464 33448
rect 4988 33439 5040 33448
rect 4988 33405 4997 33439
rect 4997 33405 5031 33439
rect 5031 33405 5040 33439
rect 4988 33396 5040 33405
rect 1915 33158 1967 33210
rect 1979 33158 2031 33210
rect 2043 33158 2095 33210
rect 2107 33158 2159 33210
rect 2171 33158 2223 33210
rect 3846 33158 3898 33210
rect 3910 33158 3962 33210
rect 3974 33158 4026 33210
rect 4038 33158 4090 33210
rect 4102 33158 4154 33210
rect 5776 33158 5828 33210
rect 5840 33158 5892 33210
rect 5904 33158 5956 33210
rect 5968 33158 6020 33210
rect 6032 33158 6084 33210
rect 5264 32895 5316 32904
rect 5264 32861 5273 32895
rect 5273 32861 5307 32895
rect 5307 32861 5316 32895
rect 5264 32852 5316 32861
rect 2880 32614 2932 32666
rect 2944 32614 2996 32666
rect 3008 32614 3060 32666
rect 3072 32614 3124 32666
rect 3136 32614 3188 32666
rect 4811 32614 4863 32666
rect 4875 32614 4927 32666
rect 4939 32614 4991 32666
rect 5003 32614 5055 32666
rect 5067 32614 5119 32666
rect 2044 32487 2096 32496
rect 2044 32453 2053 32487
rect 2053 32453 2087 32487
rect 2087 32453 2096 32487
rect 2044 32444 2096 32453
rect 1400 32376 1452 32428
rect 5632 32376 5684 32428
rect 4988 32351 5040 32360
rect 4988 32317 4997 32351
rect 4997 32317 5031 32351
rect 5031 32317 5040 32351
rect 4988 32308 5040 32317
rect 5172 32308 5224 32360
rect 5448 32308 5500 32360
rect 1915 32070 1967 32122
rect 1979 32070 2031 32122
rect 2043 32070 2095 32122
rect 2107 32070 2159 32122
rect 2171 32070 2223 32122
rect 3846 32070 3898 32122
rect 3910 32070 3962 32122
rect 3974 32070 4026 32122
rect 4038 32070 4090 32122
rect 4102 32070 4154 32122
rect 5776 32070 5828 32122
rect 5840 32070 5892 32122
rect 5904 32070 5956 32122
rect 5968 32070 6020 32122
rect 6032 32070 6084 32122
rect 1400 31968 1452 32020
rect 1768 31968 1820 32020
rect 2596 31968 2648 32020
rect 4344 31832 4396 31884
rect 1860 31807 1912 31816
rect 1860 31773 1869 31807
rect 1869 31773 1903 31807
rect 1903 31773 1912 31807
rect 1860 31764 1912 31773
rect 3424 31764 3476 31816
rect 6828 31832 6880 31884
rect 4344 31740 4396 31792
rect 6828 31696 6880 31748
rect 2880 31526 2932 31578
rect 2944 31526 2996 31578
rect 3008 31526 3060 31578
rect 3072 31526 3124 31578
rect 3136 31526 3188 31578
rect 4811 31526 4863 31578
rect 4875 31526 4927 31578
rect 4939 31526 4991 31578
rect 5003 31526 5055 31578
rect 5067 31526 5119 31578
rect 1400 31288 1452 31340
rect 6184 31288 6236 31340
rect 1915 30982 1967 31034
rect 1979 30982 2031 31034
rect 2043 30982 2095 31034
rect 2107 30982 2159 31034
rect 2171 30982 2223 31034
rect 3846 30982 3898 31034
rect 3910 30982 3962 31034
rect 3974 30982 4026 31034
rect 4038 30982 4090 31034
rect 4102 30982 4154 31034
rect 5776 30982 5828 31034
rect 5840 30982 5892 31034
rect 5904 30982 5956 31034
rect 5968 30982 6020 31034
rect 6032 30982 6084 31034
rect 5264 30923 5316 30932
rect 5264 30889 5273 30923
rect 5273 30889 5307 30923
rect 5307 30889 5316 30923
rect 5264 30880 5316 30889
rect 5172 30812 5224 30864
rect 5448 30812 5500 30864
rect 2412 30744 2464 30796
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 5448 30719 5500 30728
rect 5448 30685 5457 30719
rect 5457 30685 5491 30719
rect 5491 30685 5500 30719
rect 5448 30676 5500 30685
rect 6184 30676 6236 30728
rect 5080 30608 5132 30660
rect 5540 30608 5592 30660
rect 2880 30438 2932 30490
rect 2944 30438 2996 30490
rect 3008 30438 3060 30490
rect 3072 30438 3124 30490
rect 3136 30438 3188 30490
rect 4811 30438 4863 30490
rect 4875 30438 4927 30490
rect 4939 30438 4991 30490
rect 5003 30438 5055 30490
rect 5067 30438 5119 30490
rect 3700 30268 3752 30320
rect 1400 30200 1452 30252
rect 5356 30243 5408 30252
rect 5356 30209 5365 30243
rect 5365 30209 5399 30243
rect 5399 30209 5408 30243
rect 5356 30200 5408 30209
rect 1768 30064 1820 30116
rect 1915 29894 1967 29946
rect 1979 29894 2031 29946
rect 2043 29894 2095 29946
rect 2107 29894 2159 29946
rect 2171 29894 2223 29946
rect 3846 29894 3898 29946
rect 3910 29894 3962 29946
rect 3974 29894 4026 29946
rect 4038 29894 4090 29946
rect 4102 29894 4154 29946
rect 5776 29894 5828 29946
rect 5840 29894 5892 29946
rect 5904 29894 5956 29946
rect 5968 29894 6020 29946
rect 6032 29894 6084 29946
rect 1584 29724 1636 29776
rect 1768 29724 1820 29776
rect 2872 29767 2924 29776
rect 2872 29733 2881 29767
rect 2881 29733 2915 29767
rect 2915 29733 2924 29767
rect 2872 29724 2924 29733
rect 4160 29724 4212 29776
rect 5264 29724 5316 29776
rect 1584 29631 1636 29640
rect 1584 29597 1593 29631
rect 1593 29597 1627 29631
rect 1627 29597 1636 29631
rect 1584 29588 1636 29597
rect 5264 29631 5316 29640
rect 5264 29597 5273 29631
rect 5273 29597 5307 29631
rect 5307 29597 5316 29631
rect 5264 29588 5316 29597
rect 2320 29520 2372 29572
rect 2596 29452 2648 29504
rect 2880 29350 2932 29402
rect 2944 29350 2996 29402
rect 3008 29350 3060 29402
rect 3072 29350 3124 29402
rect 3136 29350 3188 29402
rect 4811 29350 4863 29402
rect 4875 29350 4927 29402
rect 4939 29350 4991 29402
rect 5003 29350 5055 29402
rect 5067 29350 5119 29402
rect 5356 29248 5408 29300
rect 2596 29180 2648 29232
rect 4160 29180 4212 29232
rect 1400 29112 1452 29164
rect 2412 29112 2464 29164
rect 3332 29112 3384 29164
rect 2688 29044 2740 29096
rect 4988 29087 5040 29096
rect 4988 29053 4997 29087
rect 4997 29053 5031 29087
rect 5031 29053 5040 29087
rect 4988 29044 5040 29053
rect 3424 28976 3476 29028
rect 5264 28976 5316 29028
rect 1915 28806 1967 28858
rect 1979 28806 2031 28858
rect 2043 28806 2095 28858
rect 2107 28806 2159 28858
rect 2171 28806 2223 28858
rect 3846 28806 3898 28858
rect 3910 28806 3962 28858
rect 3974 28806 4026 28858
rect 4038 28806 4090 28858
rect 4102 28806 4154 28858
rect 5776 28806 5828 28858
rect 5840 28806 5892 28858
rect 5904 28806 5956 28858
rect 5968 28806 6020 28858
rect 6032 28806 6084 28858
rect 1768 28747 1820 28756
rect 1768 28713 1777 28747
rect 1777 28713 1811 28747
rect 1811 28713 1820 28747
rect 1768 28704 1820 28713
rect 5172 28747 5224 28756
rect 5172 28713 5181 28747
rect 5181 28713 5215 28747
rect 5215 28713 5224 28747
rect 5172 28704 5224 28713
rect 6092 28543 6144 28552
rect 6092 28509 6101 28543
rect 6101 28509 6135 28543
rect 6135 28509 6144 28543
rect 6092 28500 6144 28509
rect 2228 28432 2280 28484
rect 2880 28262 2932 28314
rect 2944 28262 2996 28314
rect 3008 28262 3060 28314
rect 3072 28262 3124 28314
rect 3136 28262 3188 28314
rect 4811 28262 4863 28314
rect 4875 28262 4927 28314
rect 4939 28262 4991 28314
rect 5003 28262 5055 28314
rect 5067 28262 5119 28314
rect 1676 28160 1728 28212
rect 2228 28203 2280 28212
rect 2228 28169 2237 28203
rect 2237 28169 2271 28203
rect 2271 28169 2280 28203
rect 2228 28160 2280 28169
rect 2780 28024 2832 28076
rect 6184 28024 6236 28076
rect 5172 27956 5224 28008
rect 5540 27820 5592 27872
rect 1915 27718 1967 27770
rect 1979 27718 2031 27770
rect 2043 27718 2095 27770
rect 2107 27718 2159 27770
rect 2171 27718 2223 27770
rect 3846 27718 3898 27770
rect 3910 27718 3962 27770
rect 3974 27718 4026 27770
rect 4038 27718 4090 27770
rect 4102 27718 4154 27770
rect 5776 27718 5828 27770
rect 5840 27718 5892 27770
rect 5904 27718 5956 27770
rect 5968 27718 6020 27770
rect 6032 27718 6084 27770
rect 6460 27480 6512 27532
rect 5632 27412 5684 27464
rect 5816 27455 5868 27464
rect 5816 27421 5825 27455
rect 5825 27421 5859 27455
rect 5859 27421 5868 27455
rect 5816 27412 5868 27421
rect 1676 27344 1728 27396
rect 2044 27344 2096 27396
rect 2880 27174 2932 27226
rect 2944 27174 2996 27226
rect 3008 27174 3060 27226
rect 3072 27174 3124 27226
rect 3136 27174 3188 27226
rect 4811 27174 4863 27226
rect 4875 27174 4927 27226
rect 4939 27174 4991 27226
rect 5003 27174 5055 27226
rect 5067 27174 5119 27226
rect 2044 27072 2096 27124
rect 2504 27072 2556 27124
rect 5172 27072 5224 27124
rect 5540 27004 5592 27056
rect 1584 26979 1636 26988
rect 1584 26945 1593 26979
rect 1593 26945 1627 26979
rect 1627 26945 1636 26979
rect 1584 26936 1636 26945
rect 5080 26979 5132 26988
rect 5080 26945 5089 26979
rect 5089 26945 5123 26979
rect 5123 26945 5132 26979
rect 5080 26936 5132 26945
rect 5540 26868 5592 26920
rect 5172 26800 5224 26852
rect 5816 26800 5868 26852
rect 1915 26630 1967 26682
rect 1979 26630 2031 26682
rect 2043 26630 2095 26682
rect 2107 26630 2159 26682
rect 2171 26630 2223 26682
rect 3846 26630 3898 26682
rect 3910 26630 3962 26682
rect 3974 26630 4026 26682
rect 4038 26630 4090 26682
rect 4102 26630 4154 26682
rect 5776 26630 5828 26682
rect 5840 26630 5892 26682
rect 5904 26630 5956 26682
rect 5968 26630 6020 26682
rect 6032 26630 6084 26682
rect 2412 26528 2464 26580
rect 5264 26571 5316 26580
rect 5264 26537 5273 26571
rect 5273 26537 5307 26571
rect 5307 26537 5316 26571
rect 5264 26528 5316 26537
rect 6184 26528 6236 26580
rect 6552 26528 6604 26580
rect 5448 26460 5500 26512
rect 5264 26392 5316 26444
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 5448 26367 5500 26376
rect 5448 26333 5457 26367
rect 5457 26333 5491 26367
rect 5491 26333 5500 26367
rect 5448 26324 5500 26333
rect 6828 26188 6880 26240
rect 2880 26086 2932 26138
rect 2944 26086 2996 26138
rect 3008 26086 3060 26138
rect 3072 26086 3124 26138
rect 3136 26086 3188 26138
rect 4811 26086 4863 26138
rect 4875 26086 4927 26138
rect 4939 26086 4991 26138
rect 5003 26086 5055 26138
rect 5067 26086 5119 26138
rect 1676 25984 1728 26036
rect 4712 26027 4764 26036
rect 4712 25993 4721 26027
rect 4721 25993 4755 26027
rect 4755 25993 4764 26027
rect 4712 25984 4764 25993
rect 3700 25916 3752 25968
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 3516 25848 3568 25900
rect 4436 25780 4488 25832
rect 4712 25780 4764 25832
rect 1915 25542 1967 25594
rect 1979 25542 2031 25594
rect 2043 25542 2095 25594
rect 2107 25542 2159 25594
rect 2171 25542 2223 25594
rect 3846 25542 3898 25594
rect 3910 25542 3962 25594
rect 3974 25542 4026 25594
rect 4038 25542 4090 25594
rect 4102 25542 4154 25594
rect 5776 25542 5828 25594
rect 5840 25542 5892 25594
rect 5904 25542 5956 25594
rect 5968 25542 6020 25594
rect 6032 25542 6084 25594
rect 5172 25304 5224 25356
rect 5448 25304 5500 25356
rect 6092 25279 6144 25288
rect 6092 25245 6101 25279
rect 6101 25245 6135 25279
rect 6135 25245 6144 25279
rect 6092 25236 6144 25245
rect 5172 25211 5224 25220
rect 5172 25177 5181 25211
rect 5181 25177 5215 25211
rect 5215 25177 5224 25211
rect 5172 25168 5224 25177
rect 2880 24998 2932 25050
rect 2944 24998 2996 25050
rect 3008 24998 3060 25050
rect 3072 24998 3124 25050
rect 3136 24998 3188 25050
rect 4811 24998 4863 25050
rect 4875 24998 4927 25050
rect 4939 24998 4991 25050
rect 5003 24998 5055 25050
rect 5067 24998 5119 25050
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 6184 24760 6236 24812
rect 5540 24624 5592 24676
rect 1915 24454 1967 24506
rect 1979 24454 2031 24506
rect 2043 24454 2095 24506
rect 2107 24454 2159 24506
rect 2171 24454 2223 24506
rect 3846 24454 3898 24506
rect 3910 24454 3962 24506
rect 3974 24454 4026 24506
rect 4038 24454 4090 24506
rect 4102 24454 4154 24506
rect 5776 24454 5828 24506
rect 5840 24454 5892 24506
rect 5904 24454 5956 24506
rect 5968 24454 6020 24506
rect 6032 24454 6084 24506
rect 1492 24395 1544 24404
rect 1492 24361 1501 24395
rect 1501 24361 1535 24395
rect 1535 24361 1544 24395
rect 1492 24352 1544 24361
rect 4528 24352 4580 24404
rect 5448 24191 5500 24200
rect 5448 24157 5457 24191
rect 5457 24157 5491 24191
rect 5491 24157 5500 24191
rect 5448 24148 5500 24157
rect 6184 24148 6236 24200
rect 2780 24080 2832 24132
rect 2880 23910 2932 23962
rect 2944 23910 2996 23962
rect 3008 23910 3060 23962
rect 3072 23910 3124 23962
rect 3136 23910 3188 23962
rect 4811 23910 4863 23962
rect 4875 23910 4927 23962
rect 4939 23910 4991 23962
rect 5003 23910 5055 23962
rect 5067 23910 5119 23962
rect 5172 23808 5224 23860
rect 1584 23715 1636 23724
rect 1584 23681 1593 23715
rect 1593 23681 1627 23715
rect 1627 23681 1636 23715
rect 1584 23672 1636 23681
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 5448 23511 5500 23520
rect 5448 23477 5457 23511
rect 5457 23477 5491 23511
rect 5491 23477 5500 23511
rect 5448 23468 5500 23477
rect 6828 23468 6880 23520
rect 1915 23366 1967 23418
rect 1979 23366 2031 23418
rect 2043 23366 2095 23418
rect 2107 23366 2159 23418
rect 2171 23366 2223 23418
rect 3846 23366 3898 23418
rect 3910 23366 3962 23418
rect 3974 23366 4026 23418
rect 4038 23366 4090 23418
rect 4102 23366 4154 23418
rect 5776 23366 5828 23418
rect 5840 23366 5892 23418
rect 5904 23366 5956 23418
rect 5968 23366 6020 23418
rect 6032 23366 6084 23418
rect 3700 23264 3752 23316
rect 5540 23264 5592 23316
rect 6460 23264 6512 23316
rect 5264 23196 5316 23248
rect 1584 23103 1636 23112
rect 1584 23069 1593 23103
rect 1593 23069 1627 23103
rect 1627 23069 1636 23103
rect 1584 23060 1636 23069
rect 5264 23060 5316 23112
rect 3240 22992 3292 23044
rect 3424 22992 3476 23044
rect 6828 23060 6880 23112
rect 2880 22822 2932 22874
rect 2944 22822 2996 22874
rect 3008 22822 3060 22874
rect 3072 22822 3124 22874
rect 3136 22822 3188 22874
rect 4811 22822 4863 22874
rect 4875 22822 4927 22874
rect 4939 22822 4991 22874
rect 5003 22822 5055 22874
rect 5067 22822 5119 22874
rect 3516 22720 3568 22772
rect 5172 22720 5224 22772
rect 5632 22763 5684 22772
rect 5632 22729 5641 22763
rect 5641 22729 5675 22763
rect 5675 22729 5684 22763
rect 5632 22720 5684 22729
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 5172 22627 5224 22636
rect 5172 22593 5181 22627
rect 5181 22593 5215 22627
rect 5215 22593 5224 22627
rect 5172 22584 5224 22593
rect 6184 22584 6236 22636
rect 1915 22278 1967 22330
rect 1979 22278 2031 22330
rect 2043 22278 2095 22330
rect 2107 22278 2159 22330
rect 2171 22278 2223 22330
rect 3846 22278 3898 22330
rect 3910 22278 3962 22330
rect 3974 22278 4026 22330
rect 4038 22278 4090 22330
rect 4102 22278 4154 22330
rect 5776 22278 5828 22330
rect 5840 22278 5892 22330
rect 5904 22278 5956 22330
rect 5968 22278 6020 22330
rect 6032 22278 6084 22330
rect 5540 22176 5592 22228
rect 6460 22176 6512 22228
rect 4436 22040 4488 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 4528 21947 4580 21956
rect 4528 21913 4537 21947
rect 4537 21913 4571 21947
rect 4571 21913 4580 21947
rect 4528 21904 4580 21913
rect 5632 21947 5684 21956
rect 5632 21913 5641 21947
rect 5641 21913 5675 21947
rect 5675 21913 5684 21947
rect 5632 21904 5684 21913
rect 2780 21836 2832 21888
rect 2880 21734 2932 21786
rect 2944 21734 2996 21786
rect 3008 21734 3060 21786
rect 3072 21734 3124 21786
rect 3136 21734 3188 21786
rect 4811 21734 4863 21786
rect 4875 21734 4927 21786
rect 4939 21734 4991 21786
rect 5003 21734 5055 21786
rect 5067 21734 5119 21786
rect 5448 21632 5500 21684
rect 6184 21496 6236 21548
rect 1915 21190 1967 21242
rect 1979 21190 2031 21242
rect 2043 21190 2095 21242
rect 2107 21190 2159 21242
rect 2171 21190 2223 21242
rect 3846 21190 3898 21242
rect 3910 21190 3962 21242
rect 3974 21190 4026 21242
rect 4038 21190 4090 21242
rect 4102 21190 4154 21242
rect 5776 21190 5828 21242
rect 5840 21190 5892 21242
rect 5904 21190 5956 21242
rect 5968 21190 6020 21242
rect 6032 21190 6084 21242
rect 4528 21088 4580 21140
rect 1584 20927 1636 20936
rect 1584 20893 1593 20927
rect 1593 20893 1627 20927
rect 1627 20893 1636 20927
rect 1584 20884 1636 20893
rect 6092 20927 6144 20936
rect 6092 20893 6101 20927
rect 6101 20893 6135 20927
rect 6135 20893 6144 20927
rect 6092 20884 6144 20893
rect 2880 20646 2932 20698
rect 2944 20646 2996 20698
rect 3008 20646 3060 20698
rect 3072 20646 3124 20698
rect 3136 20646 3188 20698
rect 4811 20646 4863 20698
rect 4875 20646 4927 20698
rect 4939 20646 4991 20698
rect 5003 20646 5055 20698
rect 5067 20646 5119 20698
rect 1768 20544 1820 20596
rect 5632 20587 5684 20596
rect 5632 20553 5641 20587
rect 5641 20553 5675 20587
rect 5675 20553 5684 20587
rect 5632 20544 5684 20553
rect 1584 20451 1636 20460
rect 1584 20417 1593 20451
rect 1593 20417 1627 20451
rect 1627 20417 1636 20451
rect 1584 20408 1636 20417
rect 6184 20408 6236 20460
rect 1915 20102 1967 20154
rect 1979 20102 2031 20154
rect 2043 20102 2095 20154
rect 2107 20102 2159 20154
rect 2171 20102 2223 20154
rect 3846 20102 3898 20154
rect 3910 20102 3962 20154
rect 3974 20102 4026 20154
rect 4038 20102 4090 20154
rect 4102 20102 4154 20154
rect 5776 20102 5828 20154
rect 5840 20102 5892 20154
rect 5904 20102 5956 20154
rect 5968 20102 6020 20154
rect 6032 20102 6084 20154
rect 6736 19932 6788 19984
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 1400 19728 1452 19780
rect 2880 19558 2932 19610
rect 2944 19558 2996 19610
rect 3008 19558 3060 19610
rect 3072 19558 3124 19610
rect 3136 19558 3188 19610
rect 4811 19558 4863 19610
rect 4875 19558 4927 19610
rect 4939 19558 4991 19610
rect 5003 19558 5055 19610
rect 5067 19558 5119 19610
rect 5540 19456 5592 19508
rect 1584 19363 1636 19372
rect 1584 19329 1593 19363
rect 1593 19329 1627 19363
rect 1627 19329 1636 19363
rect 1584 19320 1636 19329
rect 6460 19252 6512 19304
rect 6368 19184 6420 19236
rect 1915 19014 1967 19066
rect 1979 19014 2031 19066
rect 2043 19014 2095 19066
rect 2107 19014 2159 19066
rect 2171 19014 2223 19066
rect 3846 19014 3898 19066
rect 3910 19014 3962 19066
rect 3974 19014 4026 19066
rect 4038 19014 4090 19066
rect 4102 19014 4154 19066
rect 5776 19014 5828 19066
rect 5840 19014 5892 19066
rect 5904 19014 5956 19066
rect 5968 19014 6020 19066
rect 6032 19014 6084 19066
rect 3240 18912 3292 18964
rect 1584 18751 1636 18760
rect 1584 18717 1593 18751
rect 1593 18717 1627 18751
rect 1627 18717 1636 18751
rect 1584 18708 1636 18717
rect 6092 18751 6144 18760
rect 6092 18717 6101 18751
rect 6101 18717 6135 18751
rect 6135 18717 6144 18751
rect 6092 18708 6144 18717
rect 2880 18470 2932 18522
rect 2944 18470 2996 18522
rect 3008 18470 3060 18522
rect 3072 18470 3124 18522
rect 3136 18470 3188 18522
rect 4811 18470 4863 18522
rect 4875 18470 4927 18522
rect 4939 18470 4991 18522
rect 5003 18470 5055 18522
rect 5067 18470 5119 18522
rect 3424 18368 3476 18420
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 6184 18232 6236 18284
rect 5540 18028 5592 18080
rect 1915 17926 1967 17978
rect 1979 17926 2031 17978
rect 2043 17926 2095 17978
rect 2107 17926 2159 17978
rect 2171 17926 2223 17978
rect 3846 17926 3898 17978
rect 3910 17926 3962 17978
rect 3974 17926 4026 17978
rect 4038 17926 4090 17978
rect 4102 17926 4154 17978
rect 5776 17926 5828 17978
rect 5840 17926 5892 17978
rect 5904 17926 5956 17978
rect 5968 17926 6020 17978
rect 6032 17926 6084 17978
rect 4620 17867 4672 17876
rect 4620 17833 4629 17867
rect 4629 17833 4663 17867
rect 4663 17833 4672 17867
rect 4620 17824 4672 17833
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 6184 17620 6236 17672
rect 4528 17595 4580 17604
rect 4528 17561 4537 17595
rect 4537 17561 4571 17595
rect 4571 17561 4580 17595
rect 4528 17552 4580 17561
rect 2880 17382 2932 17434
rect 2944 17382 2996 17434
rect 3008 17382 3060 17434
rect 3072 17382 3124 17434
rect 3136 17382 3188 17434
rect 4811 17382 4863 17434
rect 4875 17382 4927 17434
rect 4939 17382 4991 17434
rect 5003 17382 5055 17434
rect 5067 17382 5119 17434
rect 1400 17323 1452 17332
rect 1400 17289 1409 17323
rect 1409 17289 1443 17323
rect 1443 17289 1452 17323
rect 1400 17280 1452 17289
rect 4252 17280 4304 17332
rect 1584 17187 1636 17196
rect 1584 17153 1593 17187
rect 1593 17153 1627 17187
rect 1627 17153 1636 17187
rect 1584 17144 1636 17153
rect 4436 17144 4488 17196
rect 6368 17144 6420 17196
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 5632 16940 5684 16949
rect 1915 16838 1967 16890
rect 1979 16838 2031 16890
rect 2043 16838 2095 16890
rect 2107 16838 2159 16890
rect 2171 16838 2223 16890
rect 3846 16838 3898 16890
rect 3910 16838 3962 16890
rect 3974 16838 4026 16890
rect 4038 16838 4090 16890
rect 4102 16838 4154 16890
rect 5776 16838 5828 16890
rect 5840 16838 5892 16890
rect 5904 16838 5956 16890
rect 5968 16838 6020 16890
rect 6032 16838 6084 16890
rect 4344 16779 4396 16788
rect 4344 16745 4353 16779
rect 4353 16745 4387 16779
rect 4387 16745 4396 16779
rect 4344 16736 4396 16745
rect 5816 16668 5868 16720
rect 6644 16668 6696 16720
rect 5632 16600 5684 16652
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 5264 16532 5316 16584
rect 4252 16507 4304 16516
rect 4252 16473 4261 16507
rect 4261 16473 4295 16507
rect 4295 16473 4304 16507
rect 4252 16464 4304 16473
rect 5540 16464 5592 16516
rect 4436 16396 4488 16448
rect 6276 16396 6328 16448
rect 2880 16294 2932 16346
rect 2944 16294 2996 16346
rect 3008 16294 3060 16346
rect 3072 16294 3124 16346
rect 3136 16294 3188 16346
rect 4811 16294 4863 16346
rect 4875 16294 4927 16346
rect 4939 16294 4991 16346
rect 5003 16294 5055 16346
rect 5067 16294 5119 16346
rect 5816 16192 5868 16244
rect 4344 16056 4396 16108
rect 6184 16056 6236 16108
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 1915 15750 1967 15802
rect 1979 15750 2031 15802
rect 2043 15750 2095 15802
rect 2107 15750 2159 15802
rect 2171 15750 2223 15802
rect 3846 15750 3898 15802
rect 3910 15750 3962 15802
rect 3974 15750 4026 15802
rect 4038 15750 4090 15802
rect 4102 15750 4154 15802
rect 5776 15750 5828 15802
rect 5840 15750 5892 15802
rect 5904 15750 5956 15802
rect 5968 15750 6020 15802
rect 6032 15750 6084 15802
rect 4528 15648 4580 15700
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 5448 15487 5500 15496
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 6184 15444 6236 15496
rect 5540 15308 5592 15360
rect 2880 15206 2932 15258
rect 2944 15206 2996 15258
rect 3008 15206 3060 15258
rect 3072 15206 3124 15258
rect 3136 15206 3188 15258
rect 4811 15206 4863 15258
rect 4875 15206 4927 15258
rect 4939 15206 4991 15258
rect 5003 15206 5055 15258
rect 5067 15206 5119 15258
rect 4252 15104 4304 15156
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 5356 15011 5408 15020
rect 5356 14977 5365 15011
rect 5365 14977 5399 15011
rect 5399 14977 5408 15011
rect 5356 14968 5408 14977
rect 6276 14900 6328 14952
rect 1915 14662 1967 14714
rect 1979 14662 2031 14714
rect 2043 14662 2095 14714
rect 2107 14662 2159 14714
rect 2171 14662 2223 14714
rect 3846 14662 3898 14714
rect 3910 14662 3962 14714
rect 3974 14662 4026 14714
rect 4038 14662 4090 14714
rect 4102 14662 4154 14714
rect 5776 14662 5828 14714
rect 5840 14662 5892 14714
rect 5904 14662 5956 14714
rect 5968 14662 6020 14714
rect 6032 14662 6084 14714
rect 4344 14560 4396 14612
rect 5540 14560 5592 14612
rect 5356 14492 5408 14544
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 5632 14220 5684 14272
rect 2880 14118 2932 14170
rect 2944 14118 2996 14170
rect 3008 14118 3060 14170
rect 3072 14118 3124 14170
rect 3136 14118 3188 14170
rect 4811 14118 4863 14170
rect 4875 14118 4927 14170
rect 4939 14118 4991 14170
rect 5003 14118 5055 14170
rect 5067 14118 5119 14170
rect 5816 14016 5868 14068
rect 6552 13948 6604 14000
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 1915 13574 1967 13626
rect 1979 13574 2031 13626
rect 2043 13574 2095 13626
rect 2107 13574 2159 13626
rect 2171 13574 2223 13626
rect 3846 13574 3898 13626
rect 3910 13574 3962 13626
rect 3974 13574 4026 13626
rect 4038 13574 4090 13626
rect 4102 13574 4154 13626
rect 5776 13574 5828 13626
rect 5840 13574 5892 13626
rect 5904 13574 5956 13626
rect 5968 13574 6020 13626
rect 6032 13574 6084 13626
rect 3148 13472 3200 13524
rect 6460 13404 6512 13456
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 6092 13311 6144 13320
rect 6092 13277 6101 13311
rect 6101 13277 6135 13311
rect 6135 13277 6144 13311
rect 6092 13268 6144 13277
rect 1400 13200 1452 13252
rect 5540 13132 5592 13184
rect 2880 13030 2932 13082
rect 2944 13030 2996 13082
rect 3008 13030 3060 13082
rect 3072 13030 3124 13082
rect 3136 13030 3188 13082
rect 4811 13030 4863 13082
rect 4875 13030 4927 13082
rect 4939 13030 4991 13082
rect 5003 13030 5055 13082
rect 5067 13030 5119 13082
rect 1400 12971 1452 12980
rect 1400 12937 1409 12971
rect 1409 12937 1443 12971
rect 1443 12937 1452 12971
rect 1400 12928 1452 12937
rect 5632 12971 5684 12980
rect 5632 12937 5641 12971
rect 5641 12937 5675 12971
rect 5675 12937 5684 12971
rect 5632 12928 5684 12937
rect 5172 12903 5224 12912
rect 5172 12869 5181 12903
rect 5181 12869 5215 12903
rect 5215 12869 5224 12903
rect 5172 12860 5224 12869
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 4252 12792 4304 12844
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 1915 12486 1967 12538
rect 1979 12486 2031 12538
rect 2043 12486 2095 12538
rect 2107 12486 2159 12538
rect 2171 12486 2223 12538
rect 3846 12486 3898 12538
rect 3910 12486 3962 12538
rect 3974 12486 4026 12538
rect 4038 12486 4090 12538
rect 4102 12486 4154 12538
rect 5776 12486 5828 12538
rect 5840 12486 5892 12538
rect 5904 12486 5956 12538
rect 5968 12486 6020 12538
rect 6032 12486 6084 12538
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 5632 12044 5684 12096
rect 2880 11942 2932 11994
rect 2944 11942 2996 11994
rect 3008 11942 3060 11994
rect 3072 11942 3124 11994
rect 3136 11942 3188 11994
rect 4811 11942 4863 11994
rect 4875 11942 4927 11994
rect 4939 11942 4991 11994
rect 5003 11942 5055 11994
rect 5067 11942 5119 11994
rect 4252 11840 4304 11892
rect 5540 11772 5592 11824
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 5448 11704 5500 11756
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 1915 11398 1967 11450
rect 1979 11398 2031 11450
rect 2043 11398 2095 11450
rect 2107 11398 2159 11450
rect 2171 11398 2223 11450
rect 3846 11398 3898 11450
rect 3910 11398 3962 11450
rect 3974 11398 4026 11450
rect 4038 11398 4090 11450
rect 4102 11398 4154 11450
rect 5776 11398 5828 11450
rect 5840 11398 5892 11450
rect 5904 11398 5956 11450
rect 5968 11398 6020 11450
rect 6032 11398 6084 11450
rect 5448 11296 5500 11348
rect 5540 11296 5592 11348
rect 4252 11092 4304 11144
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 5356 11092 5408 11144
rect 6184 11092 6236 11144
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 2880 10854 2932 10906
rect 2944 10854 2996 10906
rect 3008 10854 3060 10906
rect 3072 10854 3124 10906
rect 3136 10854 3188 10906
rect 4811 10854 4863 10906
rect 4875 10854 4927 10906
rect 4939 10854 4991 10906
rect 5003 10854 5055 10906
rect 5067 10854 5119 10906
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 1915 10310 1967 10362
rect 1979 10310 2031 10362
rect 2043 10310 2095 10362
rect 2107 10310 2159 10362
rect 2171 10310 2223 10362
rect 3846 10310 3898 10362
rect 3910 10310 3962 10362
rect 3974 10310 4026 10362
rect 4038 10310 4090 10362
rect 4102 10310 4154 10362
rect 5776 10310 5828 10362
rect 5840 10310 5892 10362
rect 5904 10310 5956 10362
rect 5968 10310 6020 10362
rect 6032 10310 6084 10362
rect 1400 10208 1452 10260
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 2880 9766 2932 9818
rect 2944 9766 2996 9818
rect 3008 9766 3060 9818
rect 3072 9766 3124 9818
rect 3136 9766 3188 9818
rect 4811 9766 4863 9818
rect 4875 9766 4927 9818
rect 4939 9766 4991 9818
rect 5003 9766 5055 9818
rect 5067 9766 5119 9818
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 4252 9324 4304 9376
rect 1915 9222 1967 9274
rect 1979 9222 2031 9274
rect 2043 9222 2095 9274
rect 2107 9222 2159 9274
rect 2171 9222 2223 9274
rect 3846 9222 3898 9274
rect 3910 9222 3962 9274
rect 3974 9222 4026 9274
rect 4038 9222 4090 9274
rect 4102 9222 4154 9274
rect 5776 9222 5828 9274
rect 5840 9222 5892 9274
rect 5904 9222 5956 9274
rect 5968 9222 6020 9274
rect 6032 9222 6084 9274
rect 1400 9120 1452 9172
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 5632 8984 5684 9036
rect 5356 8916 5408 8968
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 4528 8780 4580 8832
rect 6184 8780 6236 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 2880 8678 2932 8730
rect 2944 8678 2996 8730
rect 3008 8678 3060 8730
rect 3072 8678 3124 8730
rect 3136 8678 3188 8730
rect 4811 8678 4863 8730
rect 4875 8678 4927 8730
rect 4939 8678 4991 8730
rect 5003 8678 5055 8730
rect 5067 8678 5119 8730
rect 1400 8576 1452 8628
rect 4252 8440 4304 8492
rect 5264 8440 5316 8492
rect 4436 8415 4488 8424
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 5448 8236 5500 8288
rect 1915 8134 1967 8186
rect 1979 8134 2031 8186
rect 2043 8134 2095 8186
rect 2107 8134 2159 8186
rect 2171 8134 2223 8186
rect 3846 8134 3898 8186
rect 3910 8134 3962 8186
rect 3974 8134 4026 8186
rect 4038 8134 4090 8186
rect 4102 8134 4154 8186
rect 5776 8134 5828 8186
rect 5840 8134 5892 8186
rect 5904 8134 5956 8186
rect 5968 8134 6020 8186
rect 6032 8134 6084 8186
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 5172 7828 5224 7880
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 4344 7692 4396 7744
rect 6276 7692 6328 7744
rect 2880 7590 2932 7642
rect 2944 7590 2996 7642
rect 3008 7590 3060 7642
rect 3072 7590 3124 7642
rect 3136 7590 3188 7642
rect 4811 7590 4863 7642
rect 4875 7590 4927 7642
rect 4939 7590 4991 7642
rect 5003 7590 5055 7642
rect 5067 7590 5119 7642
rect 1400 7488 1452 7540
rect 4436 7488 4488 7540
rect 3240 7352 3292 7404
rect 4528 7420 4580 7472
rect 4252 7352 4304 7404
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 5448 7352 5500 7404
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3700 7148 3752 7200
rect 5356 7148 5408 7200
rect 1915 7046 1967 7098
rect 1979 7046 2031 7098
rect 2043 7046 2095 7098
rect 2107 7046 2159 7098
rect 2171 7046 2223 7098
rect 3846 7046 3898 7098
rect 3910 7046 3962 7098
rect 3974 7046 4026 7098
rect 4038 7046 4090 7098
rect 4102 7046 4154 7098
rect 5776 7046 5828 7098
rect 5840 7046 5892 7098
rect 5904 7046 5956 7098
rect 5968 7046 6020 7098
rect 6032 7046 6084 7098
rect 7012 7012 7064 7064
rect 3240 6944 3292 6996
rect 4252 6944 4304 6996
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 4712 6672 4764 6724
rect 5632 6876 5684 6928
rect 6184 6672 6236 6724
rect 2880 6502 2932 6554
rect 2944 6502 2996 6554
rect 3008 6502 3060 6554
rect 3072 6502 3124 6554
rect 3136 6502 3188 6554
rect 4811 6502 4863 6554
rect 4875 6502 4927 6554
rect 4939 6502 4991 6554
rect 5003 6502 5055 6554
rect 5067 6502 5119 6554
rect 1400 6400 1452 6452
rect 4436 6400 4488 6452
rect 4344 6332 4396 6384
rect 3700 6264 3752 6316
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 4528 6128 4580 6180
rect 4436 6060 4488 6112
rect 1915 5958 1967 6010
rect 1979 5958 2031 6010
rect 2043 5958 2095 6010
rect 2107 5958 2159 6010
rect 2171 5958 2223 6010
rect 3846 5958 3898 6010
rect 3910 5958 3962 6010
rect 3974 5958 4026 6010
rect 4038 5958 4090 6010
rect 4102 5958 4154 6010
rect 5776 5958 5828 6010
rect 5840 5958 5892 6010
rect 5904 5958 5956 6010
rect 5968 5958 6020 6010
rect 6032 5958 6084 6010
rect 7012 5967 7064 5976
rect 7012 5933 7021 5967
rect 7021 5933 7055 5967
rect 7055 5933 7064 5967
rect 7012 5924 7064 5933
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 6276 5652 6328 5704
rect 4252 5584 4304 5636
rect 4712 5516 4764 5568
rect 2880 5414 2932 5466
rect 2944 5414 2996 5466
rect 3008 5414 3060 5466
rect 3072 5414 3124 5466
rect 3136 5414 3188 5466
rect 4811 5414 4863 5466
rect 4875 5414 4927 5466
rect 4939 5414 4991 5466
rect 5003 5414 5055 5466
rect 5067 5414 5119 5466
rect 5632 5312 5684 5364
rect 4804 5244 4856 5296
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 1915 4870 1967 4922
rect 1979 4870 2031 4922
rect 2043 4870 2095 4922
rect 2107 4870 2159 4922
rect 2171 4870 2223 4922
rect 3846 4870 3898 4922
rect 3910 4870 3962 4922
rect 3974 4870 4026 4922
rect 4038 4870 4090 4922
rect 4102 4870 4154 4922
rect 5776 4870 5828 4922
rect 5840 4870 5892 4922
rect 5904 4870 5956 4922
rect 5968 4870 6020 4922
rect 6032 4870 6084 4922
rect 4804 4768 4856 4820
rect 4436 4632 4488 4684
rect 4344 4564 4396 4616
rect 5172 4632 5224 4684
rect 5356 4632 5408 4684
rect 5448 4607 5500 4616
rect 4620 4496 4672 4548
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 5356 4496 5408 4548
rect 2320 4428 2372 4480
rect 2596 4471 2648 4480
rect 2596 4437 2605 4471
rect 2605 4437 2639 4471
rect 2639 4437 2648 4471
rect 2596 4428 2648 4437
rect 2780 4428 2832 4480
rect 2880 4326 2932 4378
rect 2944 4326 2996 4378
rect 3008 4326 3060 4378
rect 3072 4326 3124 4378
rect 3136 4326 3188 4378
rect 4811 4326 4863 4378
rect 4875 4326 4927 4378
rect 4939 4326 4991 4378
rect 5003 4326 5055 4378
rect 5067 4326 5119 4378
rect 1400 3952 1452 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 4528 4088 4580 4140
rect 4988 4088 5040 4140
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 5632 3884 5684 3893
rect 1915 3782 1967 3834
rect 1979 3782 2031 3834
rect 2043 3782 2095 3834
rect 2107 3782 2159 3834
rect 2171 3782 2223 3834
rect 3846 3782 3898 3834
rect 3910 3782 3962 3834
rect 3974 3782 4026 3834
rect 4038 3782 4090 3834
rect 4102 3782 4154 3834
rect 5776 3782 5828 3834
rect 5840 3782 5892 3834
rect 5904 3782 5956 3834
rect 5968 3782 6020 3834
rect 6032 3782 6084 3834
rect 4344 3723 4396 3732
rect 4344 3689 4353 3723
rect 4353 3689 4387 3723
rect 4387 3689 4396 3723
rect 4344 3680 4396 3689
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 2780 3476 2832 3528
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 5264 3476 5316 3528
rect 5632 3476 5684 3528
rect 1400 3340 1452 3392
rect 6000 3383 6052 3392
rect 6000 3349 6009 3383
rect 6009 3349 6043 3383
rect 6043 3349 6052 3383
rect 6000 3340 6052 3349
rect 2880 3238 2932 3290
rect 2944 3238 2996 3290
rect 3008 3238 3060 3290
rect 3072 3238 3124 3290
rect 3136 3238 3188 3290
rect 4811 3238 4863 3290
rect 4875 3238 4927 3290
rect 4939 3238 4991 3290
rect 5003 3238 5055 3290
rect 5067 3238 5119 3290
rect 4436 3136 4488 3188
rect 5540 3136 5592 3188
rect 4620 3068 4672 3120
rect 2596 3000 2648 3052
rect 4712 3000 4764 3052
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 6184 3000 6236 3052
rect 1492 2796 1544 2848
rect 1915 2694 1967 2746
rect 1979 2694 2031 2746
rect 2043 2694 2095 2746
rect 2107 2694 2159 2746
rect 2171 2694 2223 2746
rect 3846 2694 3898 2746
rect 3910 2694 3962 2746
rect 3974 2694 4026 2746
rect 4038 2694 4090 2746
rect 4102 2694 4154 2746
rect 5776 2694 5828 2746
rect 5840 2694 5892 2746
rect 5904 2694 5956 2746
rect 5968 2694 6020 2746
rect 6032 2694 6084 2746
rect 5448 2592 5500 2644
rect 5356 2524 5408 2576
rect 5264 2456 5316 2508
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2780 2252 2832 2304
rect 2880 2150 2932 2202
rect 2944 2150 2996 2202
rect 3008 2150 3060 2202
rect 3072 2150 3124 2202
rect 3136 2150 3188 2202
rect 4811 2150 4863 2202
rect 4875 2150 4927 2202
rect 4939 2150 4991 2202
rect 5003 2150 5055 2202
rect 5067 2150 5119 2202
<< metal2 >>
rect 4526 59664 4582 59673
rect 4526 59599 4582 59608
rect 3330 59528 3386 59537
rect 3330 59463 3386 59472
rect 3238 58712 3294 58721
rect 3238 58647 3294 58656
rect 2778 58032 2834 58041
rect 2778 57967 2834 57976
rect 2792 57594 2820 57967
rect 2880 57692 3188 57712
rect 2880 57690 2886 57692
rect 2942 57690 2966 57692
rect 3022 57690 3046 57692
rect 3102 57690 3126 57692
rect 3182 57690 3188 57692
rect 2942 57638 2944 57690
rect 3124 57638 3126 57690
rect 2880 57636 2886 57638
rect 2942 57636 2966 57638
rect 3022 57636 3046 57638
rect 3102 57636 3126 57638
rect 3182 57636 3188 57638
rect 2880 57616 3188 57636
rect 3252 57594 3280 58647
rect 2780 57588 2832 57594
rect 2780 57530 2832 57536
rect 3240 57588 3292 57594
rect 3240 57530 3292 57536
rect 2780 57452 2832 57458
rect 2780 57394 2832 57400
rect 1584 57248 1636 57254
rect 1582 57216 1584 57225
rect 1636 57216 1638 57225
rect 1582 57151 1638 57160
rect 1915 57148 2223 57168
rect 1915 57146 1921 57148
rect 1977 57146 2001 57148
rect 2057 57146 2081 57148
rect 2137 57146 2161 57148
rect 2217 57146 2223 57148
rect 1977 57094 1979 57146
rect 2159 57094 2161 57146
rect 1915 57092 1921 57094
rect 1977 57092 2001 57094
rect 2057 57092 2081 57094
rect 2137 57092 2161 57094
rect 2217 57092 2223 57094
rect 1915 57072 2223 57092
rect 1400 56840 1452 56846
rect 1400 56782 1452 56788
rect 1412 51490 1440 56782
rect 1584 56704 1636 56710
rect 1584 56646 1636 56652
rect 1596 56545 1624 56646
rect 1582 56536 1638 56545
rect 1582 56471 1638 56480
rect 1915 56060 2223 56080
rect 1915 56058 1921 56060
rect 1977 56058 2001 56060
rect 2057 56058 2081 56060
rect 2137 56058 2161 56060
rect 2217 56058 2223 56060
rect 1977 56006 1979 56058
rect 2159 56006 2161 56058
rect 1915 56004 1921 56006
rect 1977 56004 2001 56006
rect 2057 56004 2081 56006
rect 2137 56004 2161 56006
rect 2217 56004 2223 56006
rect 1915 55984 2223 56004
rect 1676 55752 1728 55758
rect 1582 55720 1638 55729
rect 1676 55694 1728 55700
rect 1582 55655 1638 55664
rect 1596 55622 1624 55655
rect 1584 55616 1636 55622
rect 1584 55558 1636 55564
rect 1492 55276 1544 55282
rect 1492 55218 1544 55224
rect 1320 51462 1440 51490
rect 1320 50402 1348 51462
rect 1400 51400 1452 51406
rect 1400 51342 1452 51348
rect 1412 51066 1440 51342
rect 1400 51060 1452 51066
rect 1400 51002 1452 51008
rect 1400 50924 1452 50930
rect 1400 50866 1452 50872
rect 1412 50522 1440 50866
rect 1400 50516 1452 50522
rect 1400 50458 1452 50464
rect 1320 50374 1440 50402
rect 1412 47138 1440 50374
rect 1320 47110 1440 47138
rect 1320 44962 1348 47110
rect 1400 47048 1452 47054
rect 1400 46990 1452 46996
rect 1412 45082 1440 46990
rect 1504 45642 1532 55218
rect 1688 55214 1716 55694
rect 2792 55418 2820 57394
rect 3240 57384 3292 57390
rect 3240 57326 3292 57332
rect 2880 56604 3188 56624
rect 2880 56602 2886 56604
rect 2942 56602 2966 56604
rect 3022 56602 3046 56604
rect 3102 56602 3126 56604
rect 3182 56602 3188 56604
rect 2942 56550 2944 56602
rect 3124 56550 3126 56602
rect 2880 56548 2886 56550
rect 2942 56548 2966 56550
rect 3022 56548 3046 56550
rect 3102 56548 3126 56550
rect 3182 56548 3188 56550
rect 2880 56528 3188 56548
rect 2880 55516 3188 55536
rect 2880 55514 2886 55516
rect 2942 55514 2966 55516
rect 3022 55514 3046 55516
rect 3102 55514 3126 55516
rect 3182 55514 3188 55516
rect 2942 55462 2944 55514
rect 3124 55462 3126 55514
rect 2880 55460 2886 55462
rect 2942 55460 2966 55462
rect 3022 55460 3046 55462
rect 3102 55460 3126 55462
rect 3182 55460 3188 55462
rect 2880 55440 3188 55460
rect 3252 55418 3280 57326
rect 3344 56506 3372 59463
rect 4250 59120 4306 59129
rect 4250 59055 4306 59064
rect 4264 57594 4292 59055
rect 4252 57588 4304 57594
rect 4252 57530 4304 57536
rect 4252 57452 4304 57458
rect 4252 57394 4304 57400
rect 3424 57384 3476 57390
rect 3424 57326 3476 57332
rect 3332 56500 3384 56506
rect 3332 56442 3384 56448
rect 3332 56364 3384 56370
rect 3332 56306 3384 56312
rect 2780 55412 2832 55418
rect 2780 55354 2832 55360
rect 3240 55412 3292 55418
rect 3240 55354 3292 55360
rect 2412 55276 2464 55282
rect 2412 55218 2464 55224
rect 1688 55186 2360 55214
rect 1584 55072 1636 55078
rect 1584 55014 1636 55020
rect 1596 54913 1624 55014
rect 1915 54972 2223 54992
rect 1915 54970 1921 54972
rect 1977 54970 2001 54972
rect 2057 54970 2081 54972
rect 2137 54970 2161 54972
rect 2217 54970 2223 54972
rect 1977 54918 1979 54970
rect 2159 54918 2161 54970
rect 1915 54916 1921 54918
rect 1977 54916 2001 54918
rect 2057 54916 2081 54918
rect 2137 54916 2161 54918
rect 2217 54916 2223 54918
rect 1582 54904 1638 54913
rect 1915 54896 2223 54916
rect 1582 54839 1638 54848
rect 1768 54664 1820 54670
rect 1768 54606 1820 54612
rect 1584 54528 1636 54534
rect 1584 54470 1636 54476
rect 1596 54233 1624 54470
rect 1582 54224 1638 54233
rect 1582 54159 1638 54168
rect 1584 53440 1636 53446
rect 1582 53408 1584 53417
rect 1636 53408 1638 53417
rect 1582 53343 1638 53352
rect 1584 52896 1636 52902
rect 1584 52838 1636 52844
rect 1596 52737 1624 52838
rect 1582 52728 1638 52737
rect 1582 52663 1638 52672
rect 1676 52012 1728 52018
rect 1676 51954 1728 51960
rect 1582 51912 1638 51921
rect 1582 51847 1584 51856
rect 1636 51847 1638 51856
rect 1584 51818 1636 51824
rect 1584 51264 1636 51270
rect 1582 51232 1584 51241
rect 1636 51232 1638 51241
rect 1582 51167 1638 51176
rect 1584 50720 1636 50726
rect 1584 50662 1636 50668
rect 1596 50425 1624 50662
rect 1582 50416 1638 50425
rect 1582 50351 1638 50360
rect 1688 49978 1716 51954
rect 1676 49972 1728 49978
rect 1676 49914 1728 49920
rect 1584 49632 1636 49638
rect 1582 49600 1584 49609
rect 1636 49600 1638 49609
rect 1582 49535 1638 49544
rect 1584 49088 1636 49094
rect 1584 49030 1636 49036
rect 1596 48929 1624 49030
rect 1582 48920 1638 48929
rect 1582 48855 1638 48864
rect 1582 48104 1638 48113
rect 1582 48039 1638 48048
rect 1596 48006 1624 48039
rect 1584 48000 1636 48006
rect 1584 47942 1636 47948
rect 1584 47456 1636 47462
rect 1582 47424 1584 47433
rect 1636 47424 1638 47433
rect 1582 47359 1638 47368
rect 1584 46912 1636 46918
rect 1584 46854 1636 46860
rect 1596 46617 1624 46854
rect 1582 46608 1638 46617
rect 1582 46543 1638 46552
rect 1584 45824 1636 45830
rect 1582 45792 1584 45801
rect 1636 45792 1638 45801
rect 1582 45727 1638 45736
rect 1504 45614 1716 45642
rect 1492 45484 1544 45490
rect 1492 45426 1544 45432
rect 1400 45076 1452 45082
rect 1400 45018 1452 45024
rect 1320 44934 1440 44962
rect 1216 43920 1268 43926
rect 1216 43862 1268 43868
rect 1124 41132 1176 41138
rect 1124 41074 1176 41080
rect 1136 33454 1164 41074
rect 1228 39914 1256 43862
rect 1412 43466 1440 44934
rect 1320 43438 1440 43466
rect 1320 41546 1348 43438
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42362 1440 43250
rect 1400 42356 1452 42362
rect 1400 42298 1452 42304
rect 1504 41857 1532 45426
rect 1584 45280 1636 45286
rect 1584 45222 1636 45228
rect 1596 45121 1624 45222
rect 1582 45112 1638 45121
rect 1582 45047 1638 45056
rect 1582 44296 1638 44305
rect 1582 44231 1584 44240
rect 1636 44231 1638 44240
rect 1584 44202 1636 44208
rect 1584 43648 1636 43654
rect 1582 43616 1584 43625
rect 1636 43616 1638 43625
rect 1582 43551 1638 43560
rect 1584 43104 1636 43110
rect 1584 43046 1636 43052
rect 1596 42809 1624 43046
rect 1582 42800 1638 42809
rect 1582 42735 1638 42744
rect 1582 42120 1638 42129
rect 1582 42055 1584 42064
rect 1636 42055 1638 42064
rect 1584 42026 1636 42032
rect 1490 41848 1546 41857
rect 1490 41783 1546 41792
rect 1688 41732 1716 45614
rect 1412 41704 1716 41732
rect 1308 41540 1360 41546
rect 1308 41482 1360 41488
rect 1412 40610 1440 41704
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1584 41472 1636 41478
rect 1490 41440 1546 41449
rect 1584 41414 1636 41420
rect 1490 41375 1546 41384
rect 1320 40582 1440 40610
rect 1216 39908 1268 39914
rect 1216 39850 1268 39856
rect 1216 39432 1268 39438
rect 1216 39374 1268 39380
rect 1228 34542 1256 39374
rect 1320 38418 1348 40582
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 38894 1440 40462
rect 1400 38888 1452 38894
rect 1400 38830 1452 38836
rect 1400 38752 1452 38758
rect 1400 38694 1452 38700
rect 1308 38412 1360 38418
rect 1308 38354 1360 38360
rect 1308 36032 1360 36038
rect 1306 36000 1308 36009
rect 1360 36000 1362 36009
rect 1306 35935 1362 35944
rect 1412 35850 1440 38694
rect 1504 36922 1532 41375
rect 1596 41313 1624 41414
rect 1582 41304 1638 41313
rect 1582 41239 1638 41248
rect 1584 40928 1636 40934
rect 1584 40870 1636 40876
rect 1596 40497 1624 40870
rect 1582 40488 1638 40497
rect 1582 40423 1638 40432
rect 1584 40384 1636 40390
rect 1584 40326 1636 40332
rect 1596 39817 1624 40326
rect 1688 40050 1716 41482
rect 1676 40044 1728 40050
rect 1676 39986 1728 39992
rect 1676 39908 1728 39914
rect 1676 39850 1728 39856
rect 1582 39808 1638 39817
rect 1582 39743 1638 39752
rect 1584 39296 1636 39302
rect 1584 39238 1636 39244
rect 1596 39001 1624 39238
rect 1688 39030 1716 39850
rect 1676 39024 1728 39030
rect 1582 38992 1638 39001
rect 1676 38966 1728 38972
rect 1582 38927 1638 38936
rect 1676 38888 1728 38894
rect 1676 38830 1728 38836
rect 1582 38312 1638 38321
rect 1582 38247 1638 38256
rect 1596 38214 1624 38247
rect 1584 38208 1636 38214
rect 1584 38150 1636 38156
rect 1584 37664 1636 37670
rect 1584 37606 1636 37612
rect 1596 37505 1624 37606
rect 1582 37496 1638 37505
rect 1582 37431 1638 37440
rect 1688 37074 1716 38830
rect 1780 37942 1808 54606
rect 1915 53884 2223 53904
rect 1915 53882 1921 53884
rect 1977 53882 2001 53884
rect 2057 53882 2081 53884
rect 2137 53882 2161 53884
rect 2217 53882 2223 53884
rect 1977 53830 1979 53882
rect 2159 53830 2161 53882
rect 1915 53828 1921 53830
rect 1977 53828 2001 53830
rect 2057 53828 2081 53830
rect 2137 53828 2161 53830
rect 2217 53828 2223 53830
rect 1915 53808 2223 53828
rect 1915 52796 2223 52816
rect 1915 52794 1921 52796
rect 1977 52794 2001 52796
rect 2057 52794 2081 52796
rect 2137 52794 2161 52796
rect 2217 52794 2223 52796
rect 1977 52742 1979 52794
rect 2159 52742 2161 52794
rect 1915 52740 1921 52742
rect 1977 52740 2001 52742
rect 2057 52740 2081 52742
rect 2137 52740 2161 52742
rect 2217 52740 2223 52742
rect 1915 52720 2223 52740
rect 1915 51708 2223 51728
rect 1915 51706 1921 51708
rect 1977 51706 2001 51708
rect 2057 51706 2081 51708
rect 2137 51706 2161 51708
rect 2217 51706 2223 51708
rect 1977 51654 1979 51706
rect 2159 51654 2161 51706
rect 1915 51652 1921 51654
rect 1977 51652 2001 51654
rect 2057 51652 2081 51654
rect 2137 51652 2161 51654
rect 2217 51652 2223 51654
rect 1915 51632 2223 51652
rect 2332 51082 2360 55186
rect 2424 51218 2452 55218
rect 2780 54596 2832 54602
rect 2780 54538 2832 54544
rect 2792 52698 2820 54538
rect 2880 54428 3188 54448
rect 2880 54426 2886 54428
rect 2942 54426 2966 54428
rect 3022 54426 3046 54428
rect 3102 54426 3126 54428
rect 3182 54426 3188 54428
rect 2942 54374 2944 54426
rect 3124 54374 3126 54426
rect 2880 54372 2886 54374
rect 2942 54372 2966 54374
rect 3022 54372 3046 54374
rect 3102 54372 3126 54374
rect 3182 54372 3188 54374
rect 2880 54352 3188 54372
rect 3344 54330 3372 56306
rect 3436 54874 3464 57326
rect 3846 57148 4154 57168
rect 3846 57146 3852 57148
rect 3908 57146 3932 57148
rect 3988 57146 4012 57148
rect 4068 57146 4092 57148
rect 4148 57146 4154 57148
rect 3908 57094 3910 57146
rect 4090 57094 4092 57146
rect 3846 57092 3852 57094
rect 3908 57092 3932 57094
rect 3988 57092 4012 57094
rect 4068 57092 4092 57094
rect 4148 57092 4154 57094
rect 3846 57072 4154 57092
rect 3846 56060 4154 56080
rect 3846 56058 3852 56060
rect 3908 56058 3932 56060
rect 3988 56058 4012 56060
rect 4068 56058 4092 56060
rect 4148 56058 4154 56060
rect 3908 56006 3910 56058
rect 4090 56006 4092 56058
rect 3846 56004 3852 56006
rect 3908 56004 3932 56006
rect 3988 56004 4012 56006
rect 4068 56004 4092 56006
rect 4148 56004 4154 56006
rect 3846 55984 4154 56004
rect 4264 55962 4292 57394
rect 4540 57050 4568 59599
rect 5262 58576 5318 58585
rect 5262 58511 5318 58520
rect 4811 57692 5119 57712
rect 4811 57690 4817 57692
rect 4873 57690 4897 57692
rect 4953 57690 4977 57692
rect 5033 57690 5057 57692
rect 5113 57690 5119 57692
rect 4873 57638 4875 57690
rect 5055 57638 5057 57690
rect 4811 57636 4817 57638
rect 4873 57636 4897 57638
rect 4953 57636 4977 57638
rect 5033 57636 5057 57638
rect 5113 57636 5119 57638
rect 4811 57616 5119 57636
rect 4712 57316 4764 57322
rect 4712 57258 4764 57264
rect 4528 57044 4580 57050
rect 4528 56986 4580 56992
rect 4344 56840 4396 56846
rect 4344 56782 4396 56788
rect 4528 56840 4580 56846
rect 4528 56782 4580 56788
rect 4252 55956 4304 55962
rect 4252 55898 4304 55904
rect 4068 55684 4120 55690
rect 4068 55626 4120 55632
rect 4080 55282 4108 55626
rect 4250 55312 4306 55321
rect 4068 55276 4120 55282
rect 4250 55247 4252 55256
rect 4068 55218 4120 55224
rect 4304 55247 4306 55256
rect 4252 55218 4304 55224
rect 4252 55140 4304 55146
rect 4252 55082 4304 55088
rect 3846 54972 4154 54992
rect 3846 54970 3852 54972
rect 3908 54970 3932 54972
rect 3988 54970 4012 54972
rect 4068 54970 4092 54972
rect 4148 54970 4154 54972
rect 3908 54918 3910 54970
rect 4090 54918 4092 54970
rect 3846 54916 3852 54918
rect 3908 54916 3932 54918
rect 3988 54916 4012 54918
rect 4068 54916 4092 54918
rect 4148 54916 4154 54918
rect 3846 54896 4154 54916
rect 3424 54868 3476 54874
rect 3424 54810 3476 54816
rect 3516 54664 3568 54670
rect 3516 54606 3568 54612
rect 3332 54324 3384 54330
rect 3332 54266 3384 54272
rect 3424 53576 3476 53582
rect 3424 53518 3476 53524
rect 2880 53340 3188 53360
rect 2880 53338 2886 53340
rect 2942 53338 2966 53340
rect 3022 53338 3046 53340
rect 3102 53338 3126 53340
rect 3182 53338 3188 53340
rect 2942 53286 2944 53338
rect 3124 53286 3126 53338
rect 2880 53284 2886 53286
rect 2942 53284 2966 53286
rect 3022 53284 3046 53286
rect 3102 53284 3126 53286
rect 3182 53284 3188 53286
rect 2880 53264 3188 53284
rect 3436 53242 3464 53518
rect 3424 53236 3476 53242
rect 3424 53178 3476 53184
rect 2872 53100 2924 53106
rect 2872 53042 2924 53048
rect 2780 52692 2832 52698
rect 2780 52634 2832 52640
rect 2884 52442 2912 53042
rect 2792 52414 2912 52442
rect 3240 52488 3292 52494
rect 3240 52430 3292 52436
rect 2424 51190 2544 51218
rect 2332 51054 2452 51082
rect 2320 50924 2372 50930
rect 2320 50866 2372 50872
rect 1915 50620 2223 50640
rect 1915 50618 1921 50620
rect 1977 50618 2001 50620
rect 2057 50618 2081 50620
rect 2137 50618 2161 50620
rect 2217 50618 2223 50620
rect 1977 50566 1979 50618
rect 2159 50566 2161 50618
rect 1915 50564 1921 50566
rect 1977 50564 2001 50566
rect 2057 50564 2081 50566
rect 2137 50564 2161 50566
rect 2217 50564 2223 50566
rect 1915 50544 2223 50564
rect 1915 49532 2223 49552
rect 1915 49530 1921 49532
rect 1977 49530 2001 49532
rect 2057 49530 2081 49532
rect 2137 49530 2161 49532
rect 2217 49530 2223 49532
rect 1977 49478 1979 49530
rect 2159 49478 2161 49530
rect 1915 49476 1921 49478
rect 1977 49476 2001 49478
rect 2057 49476 2081 49478
rect 2137 49476 2161 49478
rect 2217 49476 2223 49478
rect 1915 49456 2223 49476
rect 1915 48444 2223 48464
rect 1915 48442 1921 48444
rect 1977 48442 2001 48444
rect 2057 48442 2081 48444
rect 2137 48442 2161 48444
rect 2217 48442 2223 48444
rect 1977 48390 1979 48442
rect 2159 48390 2161 48442
rect 1915 48388 1921 48390
rect 1977 48388 2001 48390
rect 2057 48388 2081 48390
rect 2137 48388 2161 48390
rect 2217 48388 2223 48390
rect 1915 48368 2223 48388
rect 1915 47356 2223 47376
rect 1915 47354 1921 47356
rect 1977 47354 2001 47356
rect 2057 47354 2081 47356
rect 2137 47354 2161 47356
rect 2217 47354 2223 47356
rect 1977 47302 1979 47354
rect 2159 47302 2161 47354
rect 1915 47300 1921 47302
rect 1977 47300 2001 47302
rect 2057 47300 2081 47302
rect 2137 47300 2161 47302
rect 2217 47300 2223 47302
rect 1915 47280 2223 47300
rect 1915 46268 2223 46288
rect 1915 46266 1921 46268
rect 1977 46266 2001 46268
rect 2057 46266 2081 46268
rect 2137 46266 2161 46268
rect 2217 46266 2223 46268
rect 1977 46214 1979 46266
rect 2159 46214 2161 46266
rect 1915 46212 1921 46214
rect 1977 46212 2001 46214
rect 2057 46212 2081 46214
rect 2137 46212 2161 46214
rect 2217 46212 2223 46214
rect 1915 46192 2223 46212
rect 1915 45180 2223 45200
rect 1915 45178 1921 45180
rect 1977 45178 2001 45180
rect 2057 45178 2081 45180
rect 2137 45178 2161 45180
rect 2217 45178 2223 45180
rect 1977 45126 1979 45178
rect 2159 45126 2161 45178
rect 1915 45124 1921 45126
rect 1977 45124 2001 45126
rect 2057 45124 2081 45126
rect 2137 45124 2161 45126
rect 2217 45124 2223 45126
rect 1915 45104 2223 45124
rect 1915 44092 2223 44112
rect 1915 44090 1921 44092
rect 1977 44090 2001 44092
rect 2057 44090 2081 44092
rect 2137 44090 2161 44092
rect 2217 44090 2223 44092
rect 1977 44038 1979 44090
rect 2159 44038 2161 44090
rect 1915 44036 1921 44038
rect 1977 44036 2001 44038
rect 2057 44036 2081 44038
rect 2137 44036 2161 44038
rect 2217 44036 2223 44038
rect 1915 44016 2223 44036
rect 1915 43004 2223 43024
rect 1915 43002 1921 43004
rect 1977 43002 2001 43004
rect 2057 43002 2081 43004
rect 2137 43002 2161 43004
rect 2217 43002 2223 43004
rect 1977 42950 1979 43002
rect 2159 42950 2161 43002
rect 1915 42948 1921 42950
rect 1977 42948 2001 42950
rect 2057 42948 2081 42950
rect 2137 42948 2161 42950
rect 2217 42948 2223 42950
rect 1915 42928 2223 42948
rect 1915 41916 2223 41936
rect 1915 41914 1921 41916
rect 1977 41914 2001 41916
rect 2057 41914 2081 41916
rect 2137 41914 2161 41916
rect 2217 41914 2223 41916
rect 1977 41862 1979 41914
rect 2159 41862 2161 41914
rect 1915 41860 1921 41862
rect 1977 41860 2001 41862
rect 2057 41860 2081 41862
rect 2137 41860 2161 41862
rect 2217 41860 2223 41862
rect 1915 41840 2223 41860
rect 2228 41608 2280 41614
rect 2228 41550 2280 41556
rect 2240 41002 2268 41550
rect 2228 40996 2280 41002
rect 2228 40938 2280 40944
rect 1915 40828 2223 40848
rect 1915 40826 1921 40828
rect 1977 40826 2001 40828
rect 2057 40826 2081 40828
rect 2137 40826 2161 40828
rect 2217 40826 2223 40828
rect 1977 40774 1979 40826
rect 2159 40774 2161 40826
rect 1915 40772 1921 40774
rect 1977 40772 2001 40774
rect 2057 40772 2081 40774
rect 2137 40772 2161 40774
rect 2217 40772 2223 40774
rect 1915 40752 2223 40772
rect 1915 39740 2223 39760
rect 1915 39738 1921 39740
rect 1977 39738 2001 39740
rect 2057 39738 2081 39740
rect 2137 39738 2161 39740
rect 2217 39738 2223 39740
rect 1977 39686 1979 39738
rect 2159 39686 2161 39738
rect 1915 39684 1921 39686
rect 1977 39684 2001 39686
rect 2057 39684 2081 39686
rect 2137 39684 2161 39686
rect 2217 39684 2223 39686
rect 1915 39664 2223 39684
rect 1915 38652 2223 38672
rect 1915 38650 1921 38652
rect 1977 38650 2001 38652
rect 2057 38650 2081 38652
rect 2137 38650 2161 38652
rect 2217 38650 2223 38652
rect 1977 38598 1979 38650
rect 2159 38598 2161 38650
rect 1915 38596 1921 38598
rect 1977 38596 2001 38598
rect 2057 38596 2081 38598
rect 2137 38596 2161 38598
rect 2217 38596 2223 38598
rect 1915 38576 2223 38596
rect 2332 38026 2360 50866
rect 2424 44962 2452 51054
rect 2516 51074 2544 51190
rect 2516 51046 2636 51074
rect 2792 51066 2820 52414
rect 2880 52252 3188 52272
rect 2880 52250 2886 52252
rect 2942 52250 2966 52252
rect 3022 52250 3046 52252
rect 3102 52250 3126 52252
rect 3182 52250 3188 52252
rect 2942 52198 2944 52250
rect 3124 52198 3126 52250
rect 2880 52196 2886 52198
rect 2942 52196 2966 52198
rect 3022 52196 3046 52198
rect 3102 52196 3126 52198
rect 3182 52196 3188 52198
rect 2880 52176 3188 52196
rect 2880 51164 3188 51184
rect 2880 51162 2886 51164
rect 2942 51162 2966 51164
rect 3022 51162 3046 51164
rect 3102 51162 3126 51164
rect 3182 51162 3188 51164
rect 2942 51110 2944 51162
rect 3124 51110 3126 51162
rect 2880 51108 2886 51110
rect 2942 51108 2966 51110
rect 3022 51108 3046 51110
rect 3102 51108 3126 51110
rect 3182 51108 3188 51110
rect 2880 51088 3188 51108
rect 2424 44934 2544 44962
rect 2412 44872 2464 44878
rect 2412 44814 2464 44820
rect 2424 41138 2452 44814
rect 2516 43926 2544 44934
rect 2504 43920 2556 43926
rect 2504 43862 2556 43868
rect 2504 43784 2556 43790
rect 2504 43726 2556 43732
rect 2412 41132 2464 41138
rect 2412 41074 2464 41080
rect 2412 40996 2464 41002
rect 2412 40938 2464 40944
rect 2424 38729 2452 40938
rect 2516 38758 2544 43726
rect 2608 41138 2636 51046
rect 2780 51060 2832 51066
rect 2780 51002 2832 51008
rect 2780 50924 2832 50930
rect 2780 50866 2832 50872
rect 2688 45960 2740 45966
rect 2688 45902 2740 45908
rect 2596 41132 2648 41138
rect 2596 41074 2648 41080
rect 2596 40996 2648 41002
rect 2596 40938 2648 40944
rect 2504 38752 2556 38758
rect 2410 38720 2466 38729
rect 2504 38694 2556 38700
rect 2410 38655 2466 38664
rect 2608 38457 2636 40938
rect 2594 38448 2650 38457
rect 2594 38383 2650 38392
rect 2596 38344 2648 38350
rect 2596 38286 2648 38292
rect 2332 37998 2544 38026
rect 1768 37936 1820 37942
rect 1768 37878 1820 37884
rect 2412 37936 2464 37942
rect 2412 37878 2464 37884
rect 2320 37868 2372 37874
rect 2320 37810 2372 37816
rect 1915 37564 2223 37584
rect 1915 37562 1921 37564
rect 1977 37562 2001 37564
rect 2057 37562 2081 37564
rect 2137 37562 2161 37564
rect 2217 37562 2223 37564
rect 1977 37510 1979 37562
rect 2159 37510 2161 37562
rect 1915 37508 1921 37510
rect 1977 37508 2001 37510
rect 2057 37508 2081 37510
rect 2137 37508 2161 37510
rect 2217 37508 2223 37510
rect 1915 37488 2223 37508
rect 1596 37046 1716 37074
rect 1492 36916 1544 36922
rect 1492 36858 1544 36864
rect 1596 36802 1624 37046
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1504 36774 1624 36802
rect 1676 36780 1728 36786
rect 1504 36258 1532 36774
rect 1676 36722 1728 36728
rect 1582 36680 1638 36689
rect 1582 36615 1584 36624
rect 1636 36615 1638 36624
rect 1584 36586 1636 36592
rect 1504 36230 1624 36258
rect 1492 36168 1544 36174
rect 1492 36110 1544 36116
rect 1320 35822 1440 35850
rect 1320 35034 1348 35822
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1412 35193 1440 35634
rect 1398 35184 1454 35193
rect 1398 35119 1454 35128
rect 1320 35006 1440 35034
rect 1216 34536 1268 34542
rect 1216 34478 1268 34484
rect 1412 34134 1440 35006
rect 1400 34128 1452 34134
rect 1400 34070 1452 34076
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1124 33448 1176 33454
rect 1124 33390 1176 33396
rect 1412 33017 1440 33458
rect 1398 33008 1454 33017
rect 1398 32943 1454 32952
rect 1400 32428 1452 32434
rect 1400 32370 1452 32376
rect 1412 32201 1440 32370
rect 1398 32192 1454 32201
rect 1398 32127 1454 32136
rect 1400 32020 1452 32026
rect 1400 31962 1452 31968
rect 1412 31346 1440 31962
rect 1400 31340 1452 31346
rect 1400 31282 1452 31288
rect 1400 30728 1452 30734
rect 1398 30696 1400 30705
rect 1452 30696 1454 30705
rect 1398 30631 1454 30640
rect 1400 30252 1452 30258
rect 1400 30194 1452 30200
rect 1412 29889 1440 30194
rect 1398 29880 1454 29889
rect 1398 29815 1454 29824
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 28393 1440 29106
rect 1398 28384 1454 28393
rect 1398 28319 1454 28328
rect 1504 24410 1532 36110
rect 1596 34218 1624 36230
rect 1688 34377 1716 36722
rect 1674 34368 1730 34377
rect 1674 34303 1730 34312
rect 1596 34190 1716 34218
rect 1582 34096 1638 34105
rect 1582 34031 1638 34040
rect 1596 29782 1624 34031
rect 1584 29776 1636 29782
rect 1584 29718 1636 29724
rect 1584 29640 1636 29646
rect 1584 29582 1636 29588
rect 1596 29209 1624 29582
rect 1582 29200 1638 29209
rect 1582 29135 1638 29144
rect 1688 28218 1716 34190
rect 1780 32026 1808 36858
rect 1915 36476 2223 36496
rect 1915 36474 1921 36476
rect 1977 36474 2001 36476
rect 2057 36474 2081 36476
rect 2137 36474 2161 36476
rect 2217 36474 2223 36476
rect 1977 36422 1979 36474
rect 2159 36422 2161 36474
rect 1915 36420 1921 36422
rect 1977 36420 2001 36422
rect 2057 36420 2081 36422
rect 2137 36420 2161 36422
rect 2217 36420 2223 36422
rect 1915 36400 2223 36420
rect 2044 36100 2096 36106
rect 2044 36042 2096 36048
rect 2056 35766 2084 36042
rect 2044 35760 2096 35766
rect 2044 35702 2096 35708
rect 1915 35388 2223 35408
rect 1915 35386 1921 35388
rect 1977 35386 2001 35388
rect 2057 35386 2081 35388
rect 2137 35386 2161 35388
rect 2217 35386 2223 35388
rect 1977 35334 1979 35386
rect 2159 35334 2161 35386
rect 1915 35332 1921 35334
rect 1977 35332 2001 35334
rect 2057 35332 2081 35334
rect 2137 35332 2161 35334
rect 2217 35332 2223 35334
rect 1915 35312 2223 35332
rect 1860 34604 1912 34610
rect 1860 34546 1912 34552
rect 1872 34513 1900 34546
rect 1858 34504 1914 34513
rect 1858 34439 1914 34448
rect 1915 34300 2223 34320
rect 1915 34298 1921 34300
rect 1977 34298 2001 34300
rect 2057 34298 2081 34300
rect 2137 34298 2161 34300
rect 2217 34298 2223 34300
rect 1977 34246 1979 34298
rect 2159 34246 2161 34298
rect 1915 34244 1921 34246
rect 1977 34244 2001 34246
rect 2057 34244 2081 34246
rect 2137 34244 2161 34246
rect 2217 34244 2223 34246
rect 1915 34224 2223 34244
rect 1860 33924 1912 33930
rect 1860 33866 1912 33872
rect 1872 33697 1900 33866
rect 1858 33688 1914 33697
rect 1858 33623 1914 33632
rect 1915 33212 2223 33232
rect 1915 33210 1921 33212
rect 1977 33210 2001 33212
rect 2057 33210 2081 33212
rect 2137 33210 2161 33212
rect 2217 33210 2223 33212
rect 1977 33158 1979 33210
rect 2159 33158 2161 33210
rect 1915 33156 1921 33158
rect 1977 33156 2001 33158
rect 2057 33156 2081 33158
rect 2137 33156 2161 33158
rect 2217 33156 2223 33158
rect 1915 33136 2223 33156
rect 2042 32872 2098 32881
rect 2042 32807 2098 32816
rect 2056 32502 2084 32807
rect 2044 32496 2096 32502
rect 2044 32438 2096 32444
rect 1915 32124 2223 32144
rect 1915 32122 1921 32124
rect 1977 32122 2001 32124
rect 2057 32122 2081 32124
rect 2137 32122 2161 32124
rect 2217 32122 2223 32124
rect 1977 32070 1979 32122
rect 2159 32070 2161 32122
rect 1915 32068 1921 32070
rect 1977 32068 2001 32070
rect 2057 32068 2081 32070
rect 2137 32068 2161 32070
rect 2217 32068 2223 32070
rect 1915 32048 2223 32068
rect 1768 32020 1820 32026
rect 1768 31962 1820 31968
rect 2332 31906 2360 37810
rect 2424 33590 2452 37878
rect 2516 35630 2544 37998
rect 2504 35624 2556 35630
rect 2504 35566 2556 35572
rect 2608 34746 2636 38286
rect 2700 37126 2728 45902
rect 2688 37120 2740 37126
rect 2688 37062 2740 37068
rect 2686 36952 2742 36961
rect 2686 36887 2742 36896
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 2596 34536 2648 34542
rect 2596 34478 2648 34484
rect 2412 33584 2464 33590
rect 2412 33526 2464 33532
rect 2412 33448 2464 33454
rect 2412 33390 2464 33396
rect 1780 31878 2360 31906
rect 1780 30122 1808 31878
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 1872 31385 1900 31758
rect 2424 31754 2452 33390
rect 2608 32026 2636 34478
rect 2700 34202 2728 36887
rect 2792 36786 2820 50866
rect 2880 50076 3188 50096
rect 2880 50074 2886 50076
rect 2942 50074 2966 50076
rect 3022 50074 3046 50076
rect 3102 50074 3126 50076
rect 3182 50074 3188 50076
rect 2942 50022 2944 50074
rect 3124 50022 3126 50074
rect 2880 50020 2886 50022
rect 2942 50020 2966 50022
rect 3022 50020 3046 50022
rect 3102 50020 3126 50022
rect 3182 50020 3188 50022
rect 2880 50000 3188 50020
rect 2880 48988 3188 49008
rect 2880 48986 2886 48988
rect 2942 48986 2966 48988
rect 3022 48986 3046 48988
rect 3102 48986 3126 48988
rect 3182 48986 3188 48988
rect 2942 48934 2944 48986
rect 3124 48934 3126 48986
rect 2880 48932 2886 48934
rect 2942 48932 2966 48934
rect 3022 48932 3046 48934
rect 3102 48932 3126 48934
rect 3182 48932 3188 48934
rect 2880 48912 3188 48932
rect 2872 48136 2924 48142
rect 2870 48104 2872 48113
rect 2924 48104 2926 48113
rect 2870 48039 2926 48048
rect 2880 47900 3188 47920
rect 2880 47898 2886 47900
rect 2942 47898 2966 47900
rect 3022 47898 3046 47900
rect 3102 47898 3126 47900
rect 3182 47898 3188 47900
rect 2942 47846 2944 47898
rect 3124 47846 3126 47898
rect 2880 47844 2886 47846
rect 2942 47844 2966 47846
rect 3022 47844 3046 47846
rect 3102 47844 3126 47846
rect 3182 47844 3188 47846
rect 2880 47824 3188 47844
rect 2880 46812 3188 46832
rect 2880 46810 2886 46812
rect 2942 46810 2966 46812
rect 3022 46810 3046 46812
rect 3102 46810 3126 46812
rect 3182 46810 3188 46812
rect 2942 46758 2944 46810
rect 3124 46758 3126 46810
rect 2880 46756 2886 46758
rect 2942 46756 2966 46758
rect 3022 46756 3046 46758
rect 3102 46756 3126 46758
rect 3182 46756 3188 46758
rect 2880 46736 3188 46756
rect 3252 46034 3280 52430
rect 3528 51074 3556 54606
rect 3846 53884 4154 53904
rect 3846 53882 3852 53884
rect 3908 53882 3932 53884
rect 3988 53882 4012 53884
rect 4068 53882 4092 53884
rect 4148 53882 4154 53884
rect 3908 53830 3910 53882
rect 4090 53830 4092 53882
rect 3846 53828 3852 53830
rect 3908 53828 3932 53830
rect 3988 53828 4012 53830
rect 4068 53828 4092 53830
rect 4148 53828 4154 53830
rect 3846 53808 4154 53828
rect 3846 52796 4154 52816
rect 3846 52794 3852 52796
rect 3908 52794 3932 52796
rect 3988 52794 4012 52796
rect 4068 52794 4092 52796
rect 4148 52794 4154 52796
rect 3908 52742 3910 52794
rect 4090 52742 4092 52794
rect 3846 52740 3852 52742
rect 3908 52740 3932 52742
rect 3988 52740 4012 52742
rect 4068 52740 4092 52742
rect 4148 52740 4154 52742
rect 3846 52720 4154 52740
rect 3700 52012 3752 52018
rect 3700 51954 3752 51960
rect 3528 51046 3648 51074
rect 3424 49768 3476 49774
rect 3424 49710 3476 49716
rect 3332 49224 3384 49230
rect 3332 49166 3384 49172
rect 3344 46714 3372 49166
rect 3436 48006 3464 49710
rect 3516 48136 3568 48142
rect 3516 48078 3568 48084
rect 3424 48000 3476 48006
rect 3424 47942 3476 47948
rect 3424 47048 3476 47054
rect 3424 46990 3476 46996
rect 3332 46708 3384 46714
rect 3332 46650 3384 46656
rect 3240 46028 3292 46034
rect 3240 45970 3292 45976
rect 3240 45824 3292 45830
rect 3240 45766 3292 45772
rect 2880 45724 3188 45744
rect 2880 45722 2886 45724
rect 2942 45722 2966 45724
rect 3022 45722 3046 45724
rect 3102 45722 3126 45724
rect 3182 45722 3188 45724
rect 2942 45670 2944 45722
rect 3124 45670 3126 45722
rect 2880 45668 2886 45670
rect 2942 45668 2966 45670
rect 3022 45668 3046 45670
rect 3102 45668 3126 45670
rect 3182 45668 3188 45670
rect 2880 45648 3188 45668
rect 2880 44636 3188 44656
rect 2880 44634 2886 44636
rect 2942 44634 2966 44636
rect 3022 44634 3046 44636
rect 3102 44634 3126 44636
rect 3182 44634 3188 44636
rect 2942 44582 2944 44634
rect 3124 44582 3126 44634
rect 2880 44580 2886 44582
rect 2942 44580 2966 44582
rect 3022 44580 3046 44582
rect 3102 44580 3126 44582
rect 3182 44580 3188 44582
rect 2880 44560 3188 44580
rect 3148 44396 3200 44402
rect 3148 44338 3200 44344
rect 3160 43761 3188 44338
rect 3146 43752 3202 43761
rect 3146 43687 3202 43696
rect 2880 43548 3188 43568
rect 2880 43546 2886 43548
rect 2942 43546 2966 43548
rect 3022 43546 3046 43548
rect 3102 43546 3126 43548
rect 3182 43546 3188 43548
rect 2942 43494 2944 43546
rect 3124 43494 3126 43546
rect 2880 43492 2886 43494
rect 2942 43492 2966 43494
rect 3022 43492 3046 43494
rect 3102 43492 3126 43494
rect 3182 43492 3188 43494
rect 2880 43472 3188 43492
rect 2880 42460 3188 42480
rect 2880 42458 2886 42460
rect 2942 42458 2966 42460
rect 3022 42458 3046 42460
rect 3102 42458 3126 42460
rect 3182 42458 3188 42460
rect 2942 42406 2944 42458
rect 3124 42406 3126 42458
rect 2880 42404 2886 42406
rect 2942 42404 2966 42406
rect 3022 42404 3046 42406
rect 3102 42404 3126 42406
rect 3182 42404 3188 42406
rect 2880 42384 3188 42404
rect 2880 41372 3188 41392
rect 2880 41370 2886 41372
rect 2942 41370 2966 41372
rect 3022 41370 3046 41372
rect 3102 41370 3126 41372
rect 3182 41370 3188 41372
rect 2942 41318 2944 41370
rect 3124 41318 3126 41370
rect 2880 41316 2886 41318
rect 2942 41316 2966 41318
rect 3022 41316 3046 41318
rect 3102 41316 3126 41318
rect 3182 41316 3188 41318
rect 2880 41296 3188 41316
rect 3252 41274 3280 45766
rect 3332 41608 3384 41614
rect 3332 41550 3384 41556
rect 3240 41268 3292 41274
rect 3240 41210 3292 41216
rect 3238 41168 3294 41177
rect 3238 41103 3294 41112
rect 2880 40284 3188 40304
rect 2880 40282 2886 40284
rect 2942 40282 2966 40284
rect 3022 40282 3046 40284
rect 3102 40282 3126 40284
rect 3182 40282 3188 40284
rect 2942 40230 2944 40282
rect 3124 40230 3126 40282
rect 2880 40228 2886 40230
rect 2942 40228 2966 40230
rect 3022 40228 3046 40230
rect 3102 40228 3126 40230
rect 3182 40228 3188 40230
rect 2880 40208 3188 40228
rect 2880 39196 3188 39216
rect 2880 39194 2886 39196
rect 2942 39194 2966 39196
rect 3022 39194 3046 39196
rect 3102 39194 3126 39196
rect 3182 39194 3188 39196
rect 2942 39142 2944 39194
rect 3124 39142 3126 39194
rect 2880 39140 2886 39142
rect 2942 39140 2966 39142
rect 3022 39140 3046 39142
rect 3102 39140 3126 39142
rect 3182 39140 3188 39142
rect 2880 39120 3188 39140
rect 3146 38992 3202 39001
rect 3146 38927 3202 38936
rect 3160 38654 3188 38927
rect 2976 38626 3188 38654
rect 2976 38350 3004 38626
rect 3056 38548 3108 38554
rect 3056 38490 3108 38496
rect 2964 38344 3016 38350
rect 2964 38286 3016 38292
rect 3068 38282 3096 38490
rect 3148 38412 3200 38418
rect 3148 38354 3200 38360
rect 3160 38282 3188 38354
rect 3056 38276 3108 38282
rect 3056 38218 3108 38224
rect 3148 38276 3200 38282
rect 3148 38218 3200 38224
rect 2880 38108 3188 38128
rect 2880 38106 2886 38108
rect 2942 38106 2966 38108
rect 3022 38106 3046 38108
rect 3102 38106 3126 38108
rect 3182 38106 3188 38108
rect 2942 38054 2944 38106
rect 3124 38054 3126 38106
rect 2880 38052 2886 38054
rect 2942 38052 2966 38054
rect 3022 38052 3046 38054
rect 3102 38052 3126 38054
rect 3182 38052 3188 38054
rect 2880 38032 3188 38052
rect 2880 37020 3188 37040
rect 2880 37018 2886 37020
rect 2942 37018 2966 37020
rect 3022 37018 3046 37020
rect 3102 37018 3126 37020
rect 3182 37018 3188 37020
rect 2942 36966 2944 37018
rect 3124 36966 3126 37018
rect 2880 36964 2886 36966
rect 2942 36964 2966 36966
rect 3022 36964 3046 36966
rect 3102 36964 3126 36966
rect 3182 36964 3188 36966
rect 2880 36944 3188 36964
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2872 36712 2924 36718
rect 2872 36654 2924 36660
rect 2780 36644 2832 36650
rect 2780 36586 2832 36592
rect 2688 34196 2740 34202
rect 2688 34138 2740 34144
rect 2792 34066 2820 36586
rect 2884 36106 2912 36654
rect 2872 36100 2924 36106
rect 2872 36042 2924 36048
rect 2880 35932 3188 35952
rect 2880 35930 2886 35932
rect 2942 35930 2966 35932
rect 3022 35930 3046 35932
rect 3102 35930 3126 35932
rect 3182 35930 3188 35932
rect 2942 35878 2944 35930
rect 3124 35878 3126 35930
rect 2880 35876 2886 35878
rect 2942 35876 2966 35878
rect 3022 35876 3046 35878
rect 3102 35876 3126 35878
rect 3182 35876 3188 35878
rect 2880 35856 3188 35876
rect 3252 35834 3280 41103
rect 3344 38554 3372 41550
rect 3436 41414 3464 46990
rect 3528 41585 3556 48078
rect 3514 41576 3570 41585
rect 3514 41511 3570 41520
rect 3436 41386 3556 41414
rect 3424 41268 3476 41274
rect 3424 41210 3476 41216
rect 3436 38554 3464 41210
rect 3528 38677 3556 41386
rect 3514 38668 3570 38677
rect 3514 38603 3570 38612
rect 3332 38548 3384 38554
rect 3332 38490 3384 38496
rect 3424 38548 3476 38554
rect 3424 38490 3476 38496
rect 3516 38344 3568 38350
rect 3516 38286 3568 38292
rect 3332 38208 3384 38214
rect 3332 38150 3384 38156
rect 3240 35828 3292 35834
rect 3240 35770 3292 35776
rect 2880 34844 3188 34864
rect 2880 34842 2886 34844
rect 2942 34842 2966 34844
rect 3022 34842 3046 34844
rect 3102 34842 3126 34844
rect 3182 34842 3188 34844
rect 2942 34790 2944 34842
rect 3124 34790 3126 34842
rect 2880 34788 2886 34790
rect 2942 34788 2966 34790
rect 3022 34788 3046 34790
rect 3102 34788 3126 34790
rect 3182 34788 3188 34790
rect 2880 34768 3188 34788
rect 2780 34060 2832 34066
rect 2780 34002 2832 34008
rect 2880 33756 3188 33776
rect 2880 33754 2886 33756
rect 2942 33754 2966 33756
rect 3022 33754 3046 33756
rect 3102 33754 3126 33756
rect 3182 33754 3188 33756
rect 2942 33702 2944 33754
rect 3124 33702 3126 33754
rect 2880 33700 2886 33702
rect 2942 33700 2966 33702
rect 3022 33700 3046 33702
rect 3102 33700 3126 33702
rect 3182 33700 3188 33702
rect 2880 33680 3188 33700
rect 2688 33652 2740 33658
rect 2688 33594 2740 33600
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2332 31726 2452 31754
rect 1858 31376 1914 31385
rect 2332 31362 2360 31726
rect 2332 31334 2544 31362
rect 1858 31311 1914 31320
rect 2410 31240 2466 31249
rect 2410 31175 2466 31184
rect 1915 31036 2223 31056
rect 1915 31034 1921 31036
rect 1977 31034 2001 31036
rect 2057 31034 2081 31036
rect 2137 31034 2161 31036
rect 2217 31034 2223 31036
rect 1977 30982 1979 31034
rect 2159 30982 2161 31034
rect 1915 30980 1921 30982
rect 1977 30980 2001 30982
rect 2057 30980 2081 30982
rect 2137 30980 2161 30982
rect 2217 30980 2223 30982
rect 1915 30960 2223 30980
rect 2424 30802 2452 31175
rect 2412 30796 2464 30802
rect 2412 30738 2464 30744
rect 1768 30116 1820 30122
rect 1768 30058 1820 30064
rect 1915 29948 2223 29968
rect 1915 29946 1921 29948
rect 1977 29946 2001 29948
rect 2057 29946 2081 29948
rect 2137 29946 2161 29948
rect 2217 29946 2223 29948
rect 1977 29894 1979 29946
rect 2159 29894 2161 29946
rect 1915 29892 1921 29894
rect 1977 29892 2001 29894
rect 2057 29892 2081 29894
rect 2137 29892 2161 29894
rect 2217 29892 2223 29894
rect 1915 29872 2223 29892
rect 1768 29776 1820 29782
rect 1768 29718 1820 29724
rect 1780 28762 1808 29718
rect 2320 29572 2372 29578
rect 2320 29514 2372 29520
rect 1915 28860 2223 28880
rect 1915 28858 1921 28860
rect 1977 28858 2001 28860
rect 2057 28858 2081 28860
rect 2137 28858 2161 28860
rect 2217 28858 2223 28860
rect 1977 28806 1979 28858
rect 2159 28806 2161 28858
rect 1915 28804 1921 28806
rect 1977 28804 2001 28806
rect 2057 28804 2081 28806
rect 2137 28804 2161 28806
rect 2217 28804 2223 28806
rect 1915 28784 2223 28804
rect 1768 28756 1820 28762
rect 1768 28698 1820 28704
rect 2228 28484 2280 28490
rect 2228 28426 2280 28432
rect 2240 28218 2268 28426
rect 1676 28212 1728 28218
rect 1676 28154 1728 28160
rect 2228 28212 2280 28218
rect 2228 28154 2280 28160
rect 1915 27772 2223 27792
rect 1915 27770 1921 27772
rect 1977 27770 2001 27772
rect 2057 27770 2081 27772
rect 2137 27770 2161 27772
rect 2217 27770 2223 27772
rect 1977 27718 1979 27770
rect 2159 27718 2161 27770
rect 1915 27716 1921 27718
rect 1977 27716 2001 27718
rect 2057 27716 2081 27718
rect 2137 27716 2161 27718
rect 2217 27716 2223 27718
rect 1915 27696 2223 27716
rect 1676 27396 1728 27402
rect 1676 27338 1728 27344
rect 2044 27396 2096 27402
rect 2044 27338 2096 27344
rect 1584 26988 1636 26994
rect 1584 26930 1636 26936
rect 1596 26897 1624 26930
rect 1582 26888 1638 26897
rect 1582 26823 1638 26832
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 26081 1624 26318
rect 1582 26072 1638 26081
rect 1688 26042 1716 27338
rect 2056 27130 2084 27338
rect 2044 27124 2096 27130
rect 2044 27066 2096 27072
rect 1915 26684 2223 26704
rect 1915 26682 1921 26684
rect 1977 26682 2001 26684
rect 2057 26682 2081 26684
rect 2137 26682 2161 26684
rect 2217 26682 2223 26684
rect 1977 26630 1979 26682
rect 2159 26630 2161 26682
rect 1915 26628 1921 26630
rect 1977 26628 2001 26630
rect 2057 26628 2081 26630
rect 2137 26628 2161 26630
rect 2217 26628 2223 26630
rect 1915 26608 2223 26628
rect 2332 26234 2360 29514
rect 2412 29164 2464 29170
rect 2412 29106 2464 29112
rect 2424 26586 2452 29106
rect 2516 27130 2544 31334
rect 2596 29504 2648 29510
rect 2596 29446 2648 29452
rect 2608 29238 2636 29446
rect 2596 29232 2648 29238
rect 2596 29174 2648 29180
rect 2700 29102 2728 33594
rect 2880 32668 3188 32688
rect 2880 32666 2886 32668
rect 2942 32666 2966 32668
rect 3022 32666 3046 32668
rect 3102 32666 3126 32668
rect 3182 32666 3188 32668
rect 2942 32614 2944 32666
rect 3124 32614 3126 32666
rect 2880 32612 2886 32614
rect 2942 32612 2966 32614
rect 3022 32612 3046 32614
rect 3102 32612 3126 32614
rect 3182 32612 3188 32614
rect 2880 32592 3188 32612
rect 2880 31580 3188 31600
rect 2880 31578 2886 31580
rect 2942 31578 2966 31580
rect 3022 31578 3046 31580
rect 3102 31578 3126 31580
rect 3182 31578 3188 31580
rect 2942 31526 2944 31578
rect 3124 31526 3126 31578
rect 2880 31524 2886 31526
rect 2942 31524 2966 31526
rect 3022 31524 3046 31526
rect 3102 31524 3126 31526
rect 3182 31524 3188 31526
rect 2880 31504 3188 31524
rect 2880 30492 3188 30512
rect 2880 30490 2886 30492
rect 2942 30490 2966 30492
rect 3022 30490 3046 30492
rect 3102 30490 3126 30492
rect 3182 30490 3188 30492
rect 2942 30438 2944 30490
rect 3124 30438 3126 30490
rect 2880 30436 2886 30438
rect 2942 30436 2966 30438
rect 3022 30436 3046 30438
rect 3102 30436 3126 30438
rect 3182 30436 3188 30438
rect 2880 30416 3188 30436
rect 2870 29880 2926 29889
rect 2870 29815 2926 29824
rect 2884 29782 2912 29815
rect 2872 29776 2924 29782
rect 2872 29718 2924 29724
rect 2880 29404 3188 29424
rect 2880 29402 2886 29404
rect 2942 29402 2966 29404
rect 3022 29402 3046 29404
rect 3102 29402 3126 29404
rect 3182 29402 3188 29404
rect 2942 29350 2944 29402
rect 3124 29350 3126 29402
rect 2880 29348 2886 29350
rect 2942 29348 2966 29350
rect 3022 29348 3046 29350
rect 3102 29348 3126 29350
rect 3182 29348 3188 29350
rect 2880 29328 3188 29348
rect 3344 29170 3372 38150
rect 3528 38026 3556 38286
rect 3436 37998 3556 38026
rect 3436 34610 3464 37998
rect 3514 37904 3570 37913
rect 3514 37839 3570 37848
rect 3424 34604 3476 34610
rect 3424 34546 3476 34552
rect 3528 33522 3556 37839
rect 3620 36650 3648 51046
rect 3608 36644 3660 36650
rect 3608 36586 3660 36592
rect 3516 33516 3568 33522
rect 3516 33458 3568 33464
rect 3424 31816 3476 31822
rect 3424 31758 3476 31764
rect 3332 29164 3384 29170
rect 3332 29106 3384 29112
rect 2688 29096 2740 29102
rect 2688 29038 2740 29044
rect 3436 29034 3464 31758
rect 3712 30326 3740 51954
rect 3846 51708 4154 51728
rect 3846 51706 3852 51708
rect 3908 51706 3932 51708
rect 3988 51706 4012 51708
rect 4068 51706 4092 51708
rect 4148 51706 4154 51708
rect 3908 51654 3910 51706
rect 4090 51654 4092 51706
rect 3846 51652 3852 51654
rect 3908 51652 3932 51654
rect 3988 51652 4012 51654
rect 4068 51652 4092 51654
rect 4148 51652 4154 51654
rect 3846 51632 4154 51652
rect 3846 50620 4154 50640
rect 3846 50618 3852 50620
rect 3908 50618 3932 50620
rect 3988 50618 4012 50620
rect 4068 50618 4092 50620
rect 4148 50618 4154 50620
rect 3908 50566 3910 50618
rect 4090 50566 4092 50618
rect 3846 50564 3852 50566
rect 3908 50564 3932 50566
rect 3988 50564 4012 50566
rect 4068 50564 4092 50566
rect 4148 50564 4154 50566
rect 3846 50544 4154 50564
rect 3846 49532 4154 49552
rect 3846 49530 3852 49532
rect 3908 49530 3932 49532
rect 3988 49530 4012 49532
rect 4068 49530 4092 49532
rect 4148 49530 4154 49532
rect 3908 49478 3910 49530
rect 4090 49478 4092 49530
rect 3846 49476 3852 49478
rect 3908 49476 3932 49478
rect 3988 49476 4012 49478
rect 4068 49476 4092 49478
rect 4148 49476 4154 49478
rect 3846 49456 4154 49476
rect 3846 48444 4154 48464
rect 3846 48442 3852 48444
rect 3908 48442 3932 48444
rect 3988 48442 4012 48444
rect 4068 48442 4092 48444
rect 4148 48442 4154 48444
rect 3908 48390 3910 48442
rect 4090 48390 4092 48442
rect 3846 48388 3852 48390
rect 3908 48388 3932 48390
rect 3988 48388 4012 48390
rect 4068 48388 4092 48390
rect 4148 48388 4154 48390
rect 3846 48368 4154 48388
rect 3846 47356 4154 47376
rect 3846 47354 3852 47356
rect 3908 47354 3932 47356
rect 3988 47354 4012 47356
rect 4068 47354 4092 47356
rect 4148 47354 4154 47356
rect 3908 47302 3910 47354
rect 4090 47302 4092 47354
rect 3846 47300 3852 47302
rect 3908 47300 3932 47302
rect 3988 47300 4012 47302
rect 4068 47300 4092 47302
rect 4148 47300 4154 47302
rect 3846 47280 4154 47300
rect 3846 46268 4154 46288
rect 3846 46266 3852 46268
rect 3908 46266 3932 46268
rect 3988 46266 4012 46268
rect 4068 46266 4092 46268
rect 4148 46266 4154 46268
rect 3908 46214 3910 46266
rect 4090 46214 4092 46266
rect 3846 46212 3852 46214
rect 3908 46212 3932 46214
rect 3988 46212 4012 46214
rect 4068 46212 4092 46214
rect 4148 46212 4154 46214
rect 3846 46192 4154 46212
rect 4264 46186 4292 55082
rect 4356 54330 4384 56782
rect 4436 55752 4488 55758
rect 4436 55694 4488 55700
rect 4344 54324 4396 54330
rect 4344 54266 4396 54272
rect 4448 50266 4476 55694
rect 4540 54874 4568 56782
rect 4724 55214 4752 57258
rect 5276 57050 5304 58511
rect 5446 58032 5502 58041
rect 5446 57967 5502 57976
rect 5460 57594 5488 57967
rect 5448 57588 5500 57594
rect 5448 57530 5500 57536
rect 6274 57488 6330 57497
rect 5540 57452 5592 57458
rect 6274 57423 6330 57432
rect 5540 57394 5592 57400
rect 5264 57044 5316 57050
rect 5264 56986 5316 56992
rect 4811 56604 5119 56624
rect 4811 56602 4817 56604
rect 4873 56602 4897 56604
rect 4953 56602 4977 56604
rect 5033 56602 5057 56604
rect 5113 56602 5119 56604
rect 4873 56550 4875 56602
rect 5055 56550 5057 56602
rect 4811 56548 4817 56550
rect 4873 56548 4897 56550
rect 4953 56548 4977 56550
rect 5033 56548 5057 56550
rect 5113 56548 5119 56550
rect 4811 56528 5119 56548
rect 4811 55516 5119 55536
rect 4811 55514 4817 55516
rect 4873 55514 4897 55516
rect 4953 55514 4977 55516
rect 5033 55514 5057 55516
rect 5113 55514 5119 55516
rect 4873 55462 4875 55514
rect 5055 55462 5057 55514
rect 4811 55460 4817 55462
rect 4873 55460 4897 55462
rect 4953 55460 4977 55462
rect 5033 55460 5057 55462
rect 5113 55460 5119 55462
rect 4811 55440 5119 55460
rect 5552 55418 5580 57394
rect 6184 57248 6236 57254
rect 6184 57190 6236 57196
rect 5776 57148 6084 57168
rect 5776 57146 5782 57148
rect 5838 57146 5862 57148
rect 5918 57146 5942 57148
rect 5998 57146 6022 57148
rect 6078 57146 6084 57148
rect 5838 57094 5840 57146
rect 6020 57094 6022 57146
rect 5776 57092 5782 57094
rect 5838 57092 5862 57094
rect 5918 57092 5942 57094
rect 5998 57092 6022 57094
rect 6078 57092 6084 57094
rect 5776 57072 6084 57092
rect 6196 56953 6224 57190
rect 6288 57050 6316 57423
rect 6276 57044 6328 57050
rect 6276 56986 6328 56992
rect 6182 56944 6238 56953
rect 6182 56879 6238 56888
rect 5632 56840 5684 56846
rect 5632 56782 5684 56788
rect 5540 55412 5592 55418
rect 5540 55354 5592 55360
rect 5644 55350 5672 56782
rect 5722 56264 5778 56273
rect 5722 56199 5724 56208
rect 5776 56199 5778 56208
rect 5724 56170 5776 56176
rect 5776 56060 6084 56080
rect 5776 56058 5782 56060
rect 5838 56058 5862 56060
rect 5918 56058 5942 56060
rect 5998 56058 6022 56060
rect 6078 56058 6084 56060
rect 5838 56006 5840 56058
rect 6020 56006 6022 56058
rect 5776 56004 5782 56006
rect 5838 56004 5862 56006
rect 5918 56004 5942 56006
rect 5998 56004 6022 56006
rect 6078 56004 6084 56006
rect 5776 55984 6084 56004
rect 5998 55720 6054 55729
rect 5998 55655 6054 55664
rect 6012 55622 6040 55655
rect 6000 55616 6052 55622
rect 6000 55558 6052 55564
rect 5632 55344 5684 55350
rect 5632 55286 5684 55292
rect 5356 55276 5408 55282
rect 5356 55218 5408 55224
rect 4724 55186 5212 55214
rect 4528 54868 4580 54874
rect 4528 54810 4580 54816
rect 4620 54528 4672 54534
rect 4620 54470 4672 54476
rect 4528 54120 4580 54126
rect 4528 54062 4580 54068
rect 4356 50238 4476 50266
rect 4356 49314 4384 50238
rect 4356 49286 4476 49314
rect 4344 49224 4396 49230
rect 4344 49166 4396 49172
rect 4356 47841 4384 49166
rect 4342 47832 4398 47841
rect 4342 47767 4398 47776
rect 4344 47660 4396 47666
rect 4344 47602 4396 47608
rect 4356 46714 4384 47602
rect 4344 46708 4396 46714
rect 4344 46650 4396 46656
rect 4264 46158 4384 46186
rect 4252 46096 4304 46102
rect 4252 46038 4304 46044
rect 3846 45180 4154 45200
rect 3846 45178 3852 45180
rect 3908 45178 3932 45180
rect 3988 45178 4012 45180
rect 4068 45178 4092 45180
rect 4148 45178 4154 45180
rect 3908 45126 3910 45178
rect 4090 45126 4092 45178
rect 3846 45124 3852 45126
rect 3908 45124 3932 45126
rect 3988 45124 4012 45126
rect 4068 45124 4092 45126
rect 4148 45124 4154 45126
rect 3846 45104 4154 45124
rect 3846 44092 4154 44112
rect 3846 44090 3852 44092
rect 3908 44090 3932 44092
rect 3988 44090 4012 44092
rect 4068 44090 4092 44092
rect 4148 44090 4154 44092
rect 3908 44038 3910 44090
rect 4090 44038 4092 44090
rect 3846 44036 3852 44038
rect 3908 44036 3932 44038
rect 3988 44036 4012 44038
rect 4068 44036 4092 44038
rect 4148 44036 4154 44038
rect 3846 44016 4154 44036
rect 3846 43004 4154 43024
rect 3846 43002 3852 43004
rect 3908 43002 3932 43004
rect 3988 43002 4012 43004
rect 4068 43002 4092 43004
rect 4148 43002 4154 43004
rect 3908 42950 3910 43002
rect 4090 42950 4092 43002
rect 3846 42948 3852 42950
rect 3908 42948 3932 42950
rect 3988 42948 4012 42950
rect 4068 42948 4092 42950
rect 4148 42948 4154 42950
rect 3846 42928 4154 42948
rect 3846 41916 4154 41936
rect 3846 41914 3852 41916
rect 3908 41914 3932 41916
rect 3988 41914 4012 41916
rect 4068 41914 4092 41916
rect 4148 41914 4154 41916
rect 3908 41862 3910 41914
rect 4090 41862 4092 41914
rect 3846 41860 3852 41862
rect 3908 41860 3932 41862
rect 3988 41860 4012 41862
rect 4068 41860 4092 41862
rect 4148 41860 4154 41862
rect 3846 41840 4154 41860
rect 4264 41682 4292 46038
rect 4356 41721 4384 46158
rect 4342 41712 4398 41721
rect 4252 41676 4304 41682
rect 4342 41647 4398 41656
rect 4252 41618 4304 41624
rect 4448 41290 4476 49286
rect 4540 41857 4568 54062
rect 4632 48822 4660 54470
rect 4811 54428 5119 54448
rect 4811 54426 4817 54428
rect 4873 54426 4897 54428
rect 4953 54426 4977 54428
rect 5033 54426 5057 54428
rect 5113 54426 5119 54428
rect 4873 54374 4875 54426
rect 5055 54374 5057 54426
rect 4811 54372 4817 54374
rect 4873 54372 4897 54374
rect 4953 54372 4977 54374
rect 5033 54372 5057 54374
rect 5113 54372 5119 54374
rect 4811 54352 5119 54372
rect 4811 53340 5119 53360
rect 4811 53338 4817 53340
rect 4873 53338 4897 53340
rect 4953 53338 4977 53340
rect 5033 53338 5057 53340
rect 5113 53338 5119 53340
rect 4873 53286 4875 53338
rect 5055 53286 5057 53338
rect 4811 53284 4817 53286
rect 4873 53284 4897 53286
rect 4953 53284 4977 53286
rect 5033 53284 5057 53286
rect 5113 53284 5119 53286
rect 4811 53264 5119 53284
rect 4811 52252 5119 52272
rect 4811 52250 4817 52252
rect 4873 52250 4897 52252
rect 4953 52250 4977 52252
rect 5033 52250 5057 52252
rect 5113 52250 5119 52252
rect 4873 52198 4875 52250
rect 5055 52198 5057 52250
rect 4811 52196 4817 52198
rect 4873 52196 4897 52198
rect 4953 52196 4977 52198
rect 5033 52196 5057 52198
rect 5113 52196 5119 52198
rect 4811 52176 5119 52196
rect 4811 51164 5119 51184
rect 4811 51162 4817 51164
rect 4873 51162 4897 51164
rect 4953 51162 4977 51164
rect 5033 51162 5057 51164
rect 5113 51162 5119 51164
rect 4873 51110 4875 51162
rect 5055 51110 5057 51162
rect 4811 51108 4817 51110
rect 4873 51108 4897 51110
rect 4953 51108 4977 51110
rect 5033 51108 5057 51110
rect 5113 51108 5119 51110
rect 4811 51088 5119 51108
rect 4811 50076 5119 50096
rect 4811 50074 4817 50076
rect 4873 50074 4897 50076
rect 4953 50074 4977 50076
rect 5033 50074 5057 50076
rect 5113 50074 5119 50076
rect 4873 50022 4875 50074
rect 5055 50022 5057 50074
rect 4811 50020 4817 50022
rect 4873 50020 4897 50022
rect 4953 50020 4977 50022
rect 5033 50020 5057 50022
rect 5113 50020 5119 50022
rect 4811 50000 5119 50020
rect 4712 49768 4764 49774
rect 4712 49710 4764 49716
rect 4620 48816 4672 48822
rect 4620 48758 4672 48764
rect 4620 48544 4672 48550
rect 4620 48486 4672 48492
rect 4632 43353 4660 48486
rect 4724 46102 4752 49710
rect 4811 48988 5119 49008
rect 4811 48986 4817 48988
rect 4873 48986 4897 48988
rect 4953 48986 4977 48988
rect 5033 48986 5057 48988
rect 5113 48986 5119 48988
rect 4873 48934 4875 48986
rect 5055 48934 5057 48986
rect 4811 48932 4817 48934
rect 4873 48932 4897 48934
rect 4953 48932 4977 48934
rect 5033 48932 5057 48934
rect 5113 48932 5119 48934
rect 4811 48912 5119 48932
rect 4804 48340 4856 48346
rect 4804 48282 4856 48288
rect 4816 48113 4844 48282
rect 4802 48104 4858 48113
rect 4802 48039 4858 48048
rect 4811 47900 5119 47920
rect 4811 47898 4817 47900
rect 4873 47898 4897 47900
rect 4953 47898 4977 47900
rect 5033 47898 5057 47900
rect 5113 47898 5119 47900
rect 4873 47846 4875 47898
rect 5055 47846 5057 47898
rect 4811 47844 4817 47846
rect 4873 47844 4897 47846
rect 4953 47844 4977 47846
rect 5033 47844 5057 47846
rect 5113 47844 5119 47846
rect 4811 47824 5119 47844
rect 4811 46812 5119 46832
rect 4811 46810 4817 46812
rect 4873 46810 4897 46812
rect 4953 46810 4977 46812
rect 5033 46810 5057 46812
rect 5113 46810 5119 46812
rect 4873 46758 4875 46810
rect 5055 46758 5057 46810
rect 4811 46756 4817 46758
rect 4873 46756 4897 46758
rect 4953 46756 4977 46758
rect 5033 46756 5057 46758
rect 5113 46756 5119 46758
rect 4811 46736 5119 46756
rect 5080 46368 5132 46374
rect 5080 46310 5132 46316
rect 4712 46096 4764 46102
rect 4712 46038 4764 46044
rect 5092 45898 5120 46310
rect 5080 45892 5132 45898
rect 5080 45834 5132 45840
rect 4811 45724 5119 45744
rect 4811 45722 4817 45724
rect 4873 45722 4897 45724
rect 4953 45722 4977 45724
rect 5033 45722 5057 45724
rect 5113 45722 5119 45724
rect 4873 45670 4875 45722
rect 5055 45670 5057 45722
rect 4811 45668 4817 45670
rect 4873 45668 4897 45670
rect 4953 45668 4977 45670
rect 5033 45668 5057 45670
rect 5113 45668 5119 45670
rect 4811 45648 5119 45668
rect 4712 45280 4764 45286
rect 4712 45222 4764 45228
rect 4618 43344 4674 43353
rect 4618 43279 4674 43288
rect 4724 41993 4752 45222
rect 4811 44636 5119 44656
rect 4811 44634 4817 44636
rect 4873 44634 4897 44636
rect 4953 44634 4977 44636
rect 5033 44634 5057 44636
rect 5113 44634 5119 44636
rect 4873 44582 4875 44634
rect 5055 44582 5057 44634
rect 4811 44580 4817 44582
rect 4873 44580 4897 44582
rect 4953 44580 4977 44582
rect 5033 44580 5057 44582
rect 5113 44580 5119 44582
rect 4811 44560 5119 44580
rect 4811 43548 5119 43568
rect 4811 43546 4817 43548
rect 4873 43546 4897 43548
rect 4953 43546 4977 43548
rect 5033 43546 5057 43548
rect 5113 43546 5119 43548
rect 4873 43494 4875 43546
rect 5055 43494 5057 43546
rect 4811 43492 4817 43494
rect 4873 43492 4897 43494
rect 4953 43492 4977 43494
rect 5033 43492 5057 43494
rect 5113 43492 5119 43494
rect 4811 43472 5119 43492
rect 4811 42460 5119 42480
rect 4811 42458 4817 42460
rect 4873 42458 4897 42460
rect 4953 42458 4977 42460
rect 5033 42458 5057 42460
rect 5113 42458 5119 42460
rect 4873 42406 4875 42458
rect 5055 42406 5057 42458
rect 4811 42404 4817 42406
rect 4873 42404 4897 42406
rect 4953 42404 4977 42406
rect 5033 42404 5057 42406
rect 5113 42404 5119 42406
rect 4811 42384 5119 42404
rect 5080 42288 5132 42294
rect 4802 42256 4858 42265
rect 5080 42230 5132 42236
rect 4802 42191 4858 42200
rect 4710 41984 4766 41993
rect 4710 41919 4766 41928
rect 4526 41848 4582 41857
rect 4526 41783 4582 41792
rect 4618 41712 4674 41721
rect 4528 41676 4580 41682
rect 4816 41698 4844 42191
rect 4618 41647 4674 41656
rect 4724 41670 4844 41698
rect 5092 41698 5120 42230
rect 5184 41818 5212 55186
rect 5368 54534 5396 55218
rect 5722 55176 5778 55185
rect 5722 55111 5724 55120
rect 5776 55111 5778 55120
rect 5724 55082 5776 55088
rect 5776 54972 6084 54992
rect 5776 54970 5782 54972
rect 5838 54970 5862 54972
rect 5918 54970 5942 54972
rect 5998 54970 6022 54972
rect 6078 54970 6084 54972
rect 5838 54918 5840 54970
rect 6020 54918 6022 54970
rect 5776 54916 5782 54918
rect 5838 54916 5862 54918
rect 5918 54916 5942 54918
rect 5998 54916 6022 54918
rect 6078 54916 6084 54918
rect 5776 54896 6084 54916
rect 5998 54632 6054 54641
rect 5998 54567 6054 54576
rect 6012 54534 6040 54567
rect 5356 54528 5408 54534
rect 5356 54470 5408 54476
rect 6000 54528 6052 54534
rect 6000 54470 6052 54476
rect 5356 54188 5408 54194
rect 5356 54130 5408 54136
rect 5264 52896 5316 52902
rect 5264 52838 5316 52844
rect 5276 46374 5304 52838
rect 5368 51074 5396 54130
rect 5722 54088 5778 54097
rect 5722 54023 5724 54032
rect 5776 54023 5778 54032
rect 5724 53994 5776 54000
rect 5776 53884 6084 53904
rect 5776 53882 5782 53884
rect 5838 53882 5862 53884
rect 5918 53882 5942 53884
rect 5998 53882 6022 53884
rect 6078 53882 6084 53884
rect 5838 53830 5840 53882
rect 6020 53830 6022 53882
rect 5776 53828 5782 53830
rect 5838 53828 5862 53830
rect 5918 53828 5942 53830
rect 5998 53828 6022 53830
rect 6078 53828 6084 53830
rect 5776 53808 6084 53828
rect 5998 53544 6054 53553
rect 5998 53479 6054 53488
rect 6012 53446 6040 53479
rect 6000 53440 6052 53446
rect 6000 53382 6052 53388
rect 6184 52896 6236 52902
rect 6182 52864 6184 52873
rect 6236 52864 6238 52873
rect 5776 52796 6084 52816
rect 6182 52799 6238 52808
rect 5776 52794 5782 52796
rect 5838 52794 5862 52796
rect 5918 52794 5942 52796
rect 5998 52794 6022 52796
rect 6078 52794 6084 52796
rect 5838 52742 5840 52794
rect 6020 52742 6022 52794
rect 5776 52740 5782 52742
rect 5838 52740 5862 52742
rect 5918 52740 5942 52742
rect 5998 52740 6022 52742
rect 6078 52740 6084 52742
rect 5776 52720 6084 52740
rect 6460 52488 6512 52494
rect 6460 52430 6512 52436
rect 6000 52352 6052 52358
rect 5998 52320 6000 52329
rect 6052 52320 6054 52329
rect 5998 52255 6054 52264
rect 6184 51808 6236 51814
rect 6182 51776 6184 51785
rect 6236 51776 6238 51785
rect 5776 51708 6084 51728
rect 6182 51711 6238 51720
rect 5776 51706 5782 51708
rect 5838 51706 5862 51708
rect 5918 51706 5942 51708
rect 5998 51706 6022 51708
rect 6078 51706 6084 51708
rect 5838 51654 5840 51706
rect 6020 51654 6022 51706
rect 5776 51652 5782 51654
rect 5838 51652 5862 51654
rect 5918 51652 5942 51654
rect 5998 51652 6022 51654
rect 6078 51652 6084 51654
rect 5776 51632 6084 51652
rect 6000 51264 6052 51270
rect 5998 51232 6000 51241
rect 6052 51232 6054 51241
rect 5998 51167 6054 51176
rect 5368 51046 5488 51074
rect 5356 48816 5408 48822
rect 5356 48758 5408 48764
rect 5264 46368 5316 46374
rect 5264 46310 5316 46316
rect 5368 46170 5396 48758
rect 5356 46164 5408 46170
rect 5356 46106 5408 46112
rect 5264 46028 5316 46034
rect 5264 45970 5316 45976
rect 5276 42129 5304 45970
rect 5356 45824 5408 45830
rect 5356 45766 5408 45772
rect 5262 42120 5318 42129
rect 5262 42055 5318 42064
rect 5172 41812 5224 41818
rect 5172 41754 5224 41760
rect 5092 41670 5212 41698
rect 4528 41618 4580 41624
rect 4356 41262 4476 41290
rect 4250 40896 4306 40905
rect 3846 40828 4154 40848
rect 4250 40831 4306 40840
rect 3846 40826 3852 40828
rect 3908 40826 3932 40828
rect 3988 40826 4012 40828
rect 4068 40826 4092 40828
rect 4148 40826 4154 40828
rect 3908 40774 3910 40826
rect 4090 40774 4092 40826
rect 3846 40772 3852 40774
rect 3908 40772 3932 40774
rect 3988 40772 4012 40774
rect 4068 40772 4092 40774
rect 4148 40772 4154 40774
rect 3846 40752 4154 40772
rect 3846 39740 4154 39760
rect 3846 39738 3852 39740
rect 3908 39738 3932 39740
rect 3988 39738 4012 39740
rect 4068 39738 4092 39740
rect 4148 39738 4154 39740
rect 3908 39686 3910 39738
rect 4090 39686 4092 39738
rect 3846 39684 3852 39686
rect 3908 39684 3932 39686
rect 3988 39684 4012 39686
rect 4068 39684 4092 39686
rect 4148 39684 4154 39686
rect 3846 39664 4154 39684
rect 3846 38652 4154 38672
rect 3846 38650 3852 38652
rect 3908 38650 3932 38652
rect 3988 38650 4012 38652
rect 4068 38650 4092 38652
rect 4148 38650 4154 38652
rect 3908 38598 3910 38650
rect 4090 38598 4092 38650
rect 3846 38596 3852 38598
rect 3908 38596 3932 38598
rect 3988 38596 4012 38598
rect 4068 38596 4092 38598
rect 4148 38596 4154 38598
rect 3846 38576 4154 38596
rect 3884 38412 3936 38418
rect 3884 38354 3936 38360
rect 3896 37874 3924 38354
rect 3884 37868 3936 37874
rect 3884 37810 3936 37816
rect 3846 37564 4154 37584
rect 3846 37562 3852 37564
rect 3908 37562 3932 37564
rect 3988 37562 4012 37564
rect 4068 37562 4092 37564
rect 4148 37562 4154 37564
rect 3908 37510 3910 37562
rect 4090 37510 4092 37562
rect 3846 37508 3852 37510
rect 3908 37508 3932 37510
rect 3988 37508 4012 37510
rect 4068 37508 4092 37510
rect 4148 37508 4154 37510
rect 3846 37488 4154 37508
rect 3884 37392 3936 37398
rect 3884 37334 3936 37340
rect 3896 36718 3924 37334
rect 3884 36712 3936 36718
rect 3884 36654 3936 36660
rect 3846 36476 4154 36496
rect 3846 36474 3852 36476
rect 3908 36474 3932 36476
rect 3988 36474 4012 36476
rect 4068 36474 4092 36476
rect 4148 36474 4154 36476
rect 3908 36422 3910 36474
rect 4090 36422 4092 36474
rect 3846 36420 3852 36422
rect 3908 36420 3932 36422
rect 3988 36420 4012 36422
rect 4068 36420 4092 36422
rect 4148 36420 4154 36422
rect 3846 36400 4154 36420
rect 3846 35388 4154 35408
rect 3846 35386 3852 35388
rect 3908 35386 3932 35388
rect 3988 35386 4012 35388
rect 4068 35386 4092 35388
rect 4148 35386 4154 35388
rect 3908 35334 3910 35386
rect 4090 35334 4092 35386
rect 3846 35332 3852 35334
rect 3908 35332 3932 35334
rect 3988 35332 4012 35334
rect 4068 35332 4092 35334
rect 4148 35332 4154 35334
rect 3846 35312 4154 35332
rect 3846 34300 4154 34320
rect 3846 34298 3852 34300
rect 3908 34298 3932 34300
rect 3988 34298 4012 34300
rect 4068 34298 4092 34300
rect 4148 34298 4154 34300
rect 3908 34246 3910 34298
rect 4090 34246 4092 34298
rect 3846 34244 3852 34246
rect 3908 34244 3932 34246
rect 3988 34244 4012 34246
rect 4068 34244 4092 34246
rect 4148 34244 4154 34246
rect 3846 34224 4154 34244
rect 3846 33212 4154 33232
rect 3846 33210 3852 33212
rect 3908 33210 3932 33212
rect 3988 33210 4012 33212
rect 4068 33210 4092 33212
rect 4148 33210 4154 33212
rect 3908 33158 3910 33210
rect 4090 33158 4092 33210
rect 3846 33156 3852 33158
rect 3908 33156 3932 33158
rect 3988 33156 4012 33158
rect 4068 33156 4092 33158
rect 4148 33156 4154 33158
rect 3846 33136 4154 33156
rect 3846 32124 4154 32144
rect 3846 32122 3852 32124
rect 3908 32122 3932 32124
rect 3988 32122 4012 32124
rect 4068 32122 4092 32124
rect 4148 32122 4154 32124
rect 3908 32070 3910 32122
rect 4090 32070 4092 32122
rect 3846 32068 3852 32070
rect 3908 32068 3932 32070
rect 3988 32068 4012 32070
rect 4068 32068 4092 32070
rect 4148 32068 4154 32070
rect 3846 32048 4154 32068
rect 3846 31036 4154 31056
rect 3846 31034 3852 31036
rect 3908 31034 3932 31036
rect 3988 31034 4012 31036
rect 4068 31034 4092 31036
rect 4148 31034 4154 31036
rect 3908 30982 3910 31034
rect 4090 30982 4092 31034
rect 3846 30980 3852 30982
rect 3908 30980 3932 30982
rect 3988 30980 4012 30982
rect 4068 30980 4092 30982
rect 4148 30980 4154 30982
rect 3846 30960 4154 30980
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 3846 29948 4154 29968
rect 3846 29946 3852 29948
rect 3908 29946 3932 29948
rect 3988 29946 4012 29948
rect 4068 29946 4092 29948
rect 4148 29946 4154 29948
rect 3908 29894 3910 29946
rect 4090 29894 4092 29946
rect 3846 29892 3852 29894
rect 3908 29892 3932 29894
rect 3988 29892 4012 29894
rect 4068 29892 4092 29894
rect 4148 29892 4154 29894
rect 3846 29872 4154 29892
rect 4160 29776 4212 29782
rect 4160 29718 4212 29724
rect 4172 29238 4200 29718
rect 4160 29232 4212 29238
rect 4160 29174 4212 29180
rect 3424 29028 3476 29034
rect 3424 28970 3476 28976
rect 3846 28860 4154 28880
rect 3846 28858 3852 28860
rect 3908 28858 3932 28860
rect 3988 28858 4012 28860
rect 4068 28858 4092 28860
rect 4148 28858 4154 28860
rect 3908 28806 3910 28858
rect 4090 28806 4092 28858
rect 3846 28804 3852 28806
rect 3908 28804 3932 28806
rect 3988 28804 4012 28806
rect 4068 28804 4092 28806
rect 4148 28804 4154 28806
rect 3846 28784 4154 28804
rect 2880 28316 3188 28336
rect 2880 28314 2886 28316
rect 2942 28314 2966 28316
rect 3022 28314 3046 28316
rect 3102 28314 3126 28316
rect 3182 28314 3188 28316
rect 2942 28262 2944 28314
rect 3124 28262 3126 28314
rect 2880 28260 2886 28262
rect 2942 28260 2966 28262
rect 3022 28260 3046 28262
rect 3102 28260 3126 28262
rect 3182 28260 3188 28262
rect 2880 28240 3188 28260
rect 2780 28076 2832 28082
rect 2780 28018 2832 28024
rect 2792 27577 2820 28018
rect 3846 27772 4154 27792
rect 3846 27770 3852 27772
rect 3908 27770 3932 27772
rect 3988 27770 4012 27772
rect 4068 27770 4092 27772
rect 4148 27770 4154 27772
rect 3908 27718 3910 27770
rect 4090 27718 4092 27770
rect 3846 27716 3852 27718
rect 3908 27716 3932 27718
rect 3988 27716 4012 27718
rect 4068 27716 4092 27718
rect 4148 27716 4154 27718
rect 3846 27696 4154 27716
rect 2778 27568 2834 27577
rect 2778 27503 2834 27512
rect 2880 27228 3188 27248
rect 2880 27226 2886 27228
rect 2942 27226 2966 27228
rect 3022 27226 3046 27228
rect 3102 27226 3126 27228
rect 3182 27226 3188 27228
rect 2942 27174 2944 27226
rect 3124 27174 3126 27226
rect 2880 27172 2886 27174
rect 2942 27172 2966 27174
rect 3022 27172 3046 27174
rect 3102 27172 3126 27174
rect 3182 27172 3188 27174
rect 2880 27152 3188 27172
rect 2504 27124 2556 27130
rect 2504 27066 2556 27072
rect 3846 26684 4154 26704
rect 3846 26682 3852 26684
rect 3908 26682 3932 26684
rect 3988 26682 4012 26684
rect 4068 26682 4092 26684
rect 4148 26682 4154 26684
rect 3908 26630 3910 26682
rect 4090 26630 4092 26682
rect 3846 26628 3852 26630
rect 3908 26628 3932 26630
rect 3988 26628 4012 26630
rect 4068 26628 4092 26630
rect 4148 26628 4154 26630
rect 3846 26608 4154 26628
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 1780 26206 2360 26234
rect 1582 26007 1638 26016
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1596 25401 1624 25842
rect 1582 25392 1638 25401
rect 1582 25327 1638 25336
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1596 24585 1624 24754
rect 1582 24576 1638 24585
rect 1582 24511 1638 24520
rect 1492 24404 1544 24410
rect 1492 24346 1544 24352
rect 1582 23896 1638 23905
rect 1582 23831 1638 23840
rect 1596 23730 1624 23831
rect 1584 23724 1636 23730
rect 1584 23666 1636 23672
rect 1584 23112 1636 23118
rect 1582 23080 1584 23089
rect 1636 23080 1638 23089
rect 1582 23015 1638 23024
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1596 22273 1624 22578
rect 1582 22264 1638 22273
rect 1582 22199 1638 22208
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21593 1624 21966
rect 1582 21584 1638 21593
rect 1582 21519 1638 21528
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1596 20777 1624 20878
rect 1582 20768 1638 20777
rect 1582 20703 1638 20712
rect 1780 20602 1808 26206
rect 2880 26140 3188 26160
rect 2880 26138 2886 26140
rect 2942 26138 2966 26140
rect 3022 26138 3046 26140
rect 3102 26138 3126 26140
rect 3182 26138 3188 26140
rect 2942 26086 2944 26138
rect 3124 26086 3126 26138
rect 2880 26084 2886 26086
rect 2942 26084 2966 26086
rect 3022 26084 3046 26086
rect 3102 26084 3126 26086
rect 3182 26084 3188 26086
rect 2880 26064 3188 26084
rect 3700 25968 3752 25974
rect 3700 25910 3752 25916
rect 3516 25900 3568 25906
rect 3516 25842 3568 25848
rect 1915 25596 2223 25616
rect 1915 25594 1921 25596
rect 1977 25594 2001 25596
rect 2057 25594 2081 25596
rect 2137 25594 2161 25596
rect 2217 25594 2223 25596
rect 1977 25542 1979 25594
rect 2159 25542 2161 25594
rect 1915 25540 1921 25542
rect 1977 25540 2001 25542
rect 2057 25540 2081 25542
rect 2137 25540 2161 25542
rect 2217 25540 2223 25542
rect 1915 25520 2223 25540
rect 2880 25052 3188 25072
rect 2880 25050 2886 25052
rect 2942 25050 2966 25052
rect 3022 25050 3046 25052
rect 3102 25050 3126 25052
rect 3182 25050 3188 25052
rect 2942 24998 2944 25050
rect 3124 24998 3126 25050
rect 2880 24996 2886 24998
rect 2942 24996 2966 24998
rect 3022 24996 3046 24998
rect 3102 24996 3126 24998
rect 3182 24996 3188 24998
rect 2880 24976 3188 24996
rect 1915 24508 2223 24528
rect 1915 24506 1921 24508
rect 1977 24506 2001 24508
rect 2057 24506 2081 24508
rect 2137 24506 2161 24508
rect 2217 24506 2223 24508
rect 1977 24454 1979 24506
rect 2159 24454 2161 24506
rect 1915 24452 1921 24454
rect 1977 24452 2001 24454
rect 2057 24452 2081 24454
rect 2137 24452 2161 24454
rect 2217 24452 2223 24454
rect 1915 24432 2223 24452
rect 2780 24132 2832 24138
rect 2780 24074 2832 24080
rect 1915 23420 2223 23440
rect 1915 23418 1921 23420
rect 1977 23418 2001 23420
rect 2057 23418 2081 23420
rect 2137 23418 2161 23420
rect 2217 23418 2223 23420
rect 1977 23366 1979 23418
rect 2159 23366 2161 23418
rect 1915 23364 1921 23366
rect 1977 23364 2001 23366
rect 2057 23364 2081 23366
rect 2137 23364 2161 23366
rect 2217 23364 2223 23366
rect 1915 23344 2223 23364
rect 1915 22332 2223 22352
rect 1915 22330 1921 22332
rect 1977 22330 2001 22332
rect 2057 22330 2081 22332
rect 2137 22330 2161 22332
rect 2217 22330 2223 22332
rect 1977 22278 1979 22330
rect 2159 22278 2161 22330
rect 1915 22276 1921 22278
rect 1977 22276 2001 22278
rect 2057 22276 2081 22278
rect 2137 22276 2161 22278
rect 2217 22276 2223 22278
rect 1915 22256 2223 22276
rect 2792 21894 2820 24074
rect 2880 23964 3188 23984
rect 2880 23962 2886 23964
rect 2942 23962 2966 23964
rect 3022 23962 3046 23964
rect 3102 23962 3126 23964
rect 3182 23962 3188 23964
rect 2942 23910 2944 23962
rect 3124 23910 3126 23962
rect 2880 23908 2886 23910
rect 2942 23908 2966 23910
rect 3022 23908 3046 23910
rect 3102 23908 3126 23910
rect 3182 23908 3188 23910
rect 2880 23888 3188 23908
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3424 23044 3476 23050
rect 3424 22986 3476 22992
rect 2880 22876 3188 22896
rect 2880 22874 2886 22876
rect 2942 22874 2966 22876
rect 3022 22874 3046 22876
rect 3102 22874 3126 22876
rect 3182 22874 3188 22876
rect 2942 22822 2944 22874
rect 3124 22822 3126 22874
rect 2880 22820 2886 22822
rect 2942 22820 2966 22822
rect 3022 22820 3046 22822
rect 3102 22820 3126 22822
rect 3182 22820 3188 22822
rect 2880 22800 3188 22820
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 2880 21788 3188 21808
rect 2880 21786 2886 21788
rect 2942 21786 2966 21788
rect 3022 21786 3046 21788
rect 3102 21786 3126 21788
rect 3182 21786 3188 21788
rect 2942 21734 2944 21786
rect 3124 21734 3126 21786
rect 2880 21732 2886 21734
rect 2942 21732 2966 21734
rect 3022 21732 3046 21734
rect 3102 21732 3126 21734
rect 3182 21732 3188 21734
rect 2880 21712 3188 21732
rect 1915 21244 2223 21264
rect 1915 21242 1921 21244
rect 1977 21242 2001 21244
rect 2057 21242 2081 21244
rect 2137 21242 2161 21244
rect 2217 21242 2223 21244
rect 1977 21190 1979 21242
rect 2159 21190 2161 21242
rect 1915 21188 1921 21190
rect 1977 21188 2001 21190
rect 2057 21188 2081 21190
rect 2137 21188 2161 21190
rect 2217 21188 2223 21190
rect 1915 21168 2223 21188
rect 2880 20700 3188 20720
rect 2880 20698 2886 20700
rect 2942 20698 2966 20700
rect 3022 20698 3046 20700
rect 3102 20698 3126 20700
rect 3182 20698 3188 20700
rect 2942 20646 2944 20698
rect 3124 20646 3126 20698
rect 2880 20644 2886 20646
rect 2942 20644 2966 20646
rect 3022 20644 3046 20646
rect 3102 20644 3126 20646
rect 3182 20644 3188 20646
rect 2880 20624 3188 20644
rect 1768 20596 1820 20602
rect 1768 20538 1820 20544
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1596 20097 1624 20402
rect 1915 20156 2223 20176
rect 1915 20154 1921 20156
rect 1977 20154 2001 20156
rect 2057 20154 2081 20156
rect 2137 20154 2161 20156
rect 2217 20154 2223 20156
rect 1977 20102 1979 20154
rect 2159 20102 2161 20154
rect 1915 20100 1921 20102
rect 1977 20100 2001 20102
rect 2057 20100 2081 20102
rect 2137 20100 2161 20102
rect 2217 20100 2223 20102
rect 1582 20088 1638 20097
rect 1915 20080 2223 20100
rect 1582 20023 1638 20032
rect 1400 19780 1452 19786
rect 1400 19722 1452 19728
rect 1412 17338 1440 19722
rect 2880 19612 3188 19632
rect 2880 19610 2886 19612
rect 2942 19610 2966 19612
rect 3022 19610 3046 19612
rect 3102 19610 3126 19612
rect 3182 19610 3188 19612
rect 2942 19558 2944 19610
rect 3124 19558 3126 19610
rect 2880 19556 2886 19558
rect 2942 19556 2966 19558
rect 3022 19556 3046 19558
rect 3102 19556 3126 19558
rect 3182 19556 3188 19558
rect 2880 19536 3188 19556
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1596 19281 1624 19314
rect 1582 19272 1638 19281
rect 1582 19207 1638 19216
rect 1915 19068 2223 19088
rect 1915 19066 1921 19068
rect 1977 19066 2001 19068
rect 2057 19066 2081 19068
rect 2137 19066 2161 19068
rect 2217 19066 2223 19068
rect 1977 19014 1979 19066
rect 2159 19014 2161 19066
rect 1915 19012 1921 19014
rect 1977 19012 2001 19014
rect 2057 19012 2081 19014
rect 2137 19012 2161 19014
rect 2217 19012 2223 19014
rect 1915 18992 2223 19012
rect 3252 18970 3280 22986
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1596 18465 1624 18702
rect 2880 18524 3188 18544
rect 2880 18522 2886 18524
rect 2942 18522 2966 18524
rect 3022 18522 3046 18524
rect 3102 18522 3126 18524
rect 3182 18522 3188 18524
rect 2942 18470 2944 18522
rect 3124 18470 3126 18522
rect 2880 18468 2886 18470
rect 2942 18468 2966 18470
rect 3022 18468 3046 18470
rect 3102 18468 3126 18470
rect 3182 18468 3188 18470
rect 1582 18456 1638 18465
rect 2880 18448 3188 18468
rect 3436 18426 3464 22986
rect 3528 22778 3556 25842
rect 3712 23322 3740 25910
rect 3846 25596 4154 25616
rect 3846 25594 3852 25596
rect 3908 25594 3932 25596
rect 3988 25594 4012 25596
rect 4068 25594 4092 25596
rect 4148 25594 4154 25596
rect 3908 25542 3910 25594
rect 4090 25542 4092 25594
rect 3846 25540 3852 25542
rect 3908 25540 3932 25542
rect 3988 25540 4012 25542
rect 4068 25540 4092 25542
rect 4148 25540 4154 25542
rect 3846 25520 4154 25540
rect 3846 24508 4154 24528
rect 3846 24506 3852 24508
rect 3908 24506 3932 24508
rect 3988 24506 4012 24508
rect 4068 24506 4092 24508
rect 4148 24506 4154 24508
rect 3908 24454 3910 24506
rect 4090 24454 4092 24506
rect 3846 24452 3852 24454
rect 3908 24452 3932 24454
rect 3988 24452 4012 24454
rect 4068 24452 4092 24454
rect 4148 24452 4154 24454
rect 3846 24432 4154 24452
rect 3846 23420 4154 23440
rect 3846 23418 3852 23420
rect 3908 23418 3932 23420
rect 3988 23418 4012 23420
rect 4068 23418 4092 23420
rect 4148 23418 4154 23420
rect 3908 23366 3910 23418
rect 4090 23366 4092 23418
rect 3846 23364 3852 23366
rect 3908 23364 3932 23366
rect 3988 23364 4012 23366
rect 4068 23364 4092 23366
rect 4148 23364 4154 23366
rect 3846 23344 4154 23364
rect 3700 23316 3752 23322
rect 3700 23258 3752 23264
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3846 22332 4154 22352
rect 3846 22330 3852 22332
rect 3908 22330 3932 22332
rect 3988 22330 4012 22332
rect 4068 22330 4092 22332
rect 4148 22330 4154 22332
rect 3908 22278 3910 22330
rect 4090 22278 4092 22330
rect 3846 22276 3852 22278
rect 3908 22276 3932 22278
rect 3988 22276 4012 22278
rect 4068 22276 4092 22278
rect 4148 22276 4154 22278
rect 3846 22256 4154 22276
rect 3846 21244 4154 21264
rect 3846 21242 3852 21244
rect 3908 21242 3932 21244
rect 3988 21242 4012 21244
rect 4068 21242 4092 21244
rect 4148 21242 4154 21244
rect 3908 21190 3910 21242
rect 4090 21190 4092 21242
rect 3846 21188 3852 21190
rect 3908 21188 3932 21190
rect 3988 21188 4012 21190
rect 4068 21188 4092 21190
rect 4148 21188 4154 21190
rect 3846 21168 4154 21188
rect 3846 20156 4154 20176
rect 3846 20154 3852 20156
rect 3908 20154 3932 20156
rect 3988 20154 4012 20156
rect 4068 20154 4092 20156
rect 4148 20154 4154 20156
rect 3908 20102 3910 20154
rect 4090 20102 4092 20154
rect 3846 20100 3852 20102
rect 3908 20100 3932 20102
rect 3988 20100 4012 20102
rect 4068 20100 4092 20102
rect 4148 20100 4154 20102
rect 3846 20080 4154 20100
rect 3846 19068 4154 19088
rect 3846 19066 3852 19068
rect 3908 19066 3932 19068
rect 3988 19066 4012 19068
rect 4068 19066 4092 19068
rect 4148 19066 4154 19068
rect 3908 19014 3910 19066
rect 4090 19014 4092 19066
rect 3846 19012 3852 19014
rect 3908 19012 3932 19014
rect 3988 19012 4012 19014
rect 4068 19012 4092 19014
rect 4148 19012 4154 19014
rect 3846 18992 4154 19012
rect 1582 18391 1638 18400
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17785 1624 18226
rect 1915 17980 2223 18000
rect 1915 17978 1921 17980
rect 1977 17978 2001 17980
rect 2057 17978 2081 17980
rect 2137 17978 2161 17980
rect 2217 17978 2223 17980
rect 1977 17926 1979 17978
rect 2159 17926 2161 17978
rect 1915 17924 1921 17926
rect 1977 17924 2001 17926
rect 2057 17924 2081 17926
rect 2137 17924 2161 17926
rect 2217 17924 2223 17926
rect 1915 17904 2223 17924
rect 3846 17980 4154 18000
rect 3846 17978 3852 17980
rect 3908 17978 3932 17980
rect 3988 17978 4012 17980
rect 4068 17978 4092 17980
rect 4148 17978 4154 17980
rect 3908 17926 3910 17978
rect 4090 17926 4092 17978
rect 3846 17924 3852 17926
rect 3908 17924 3932 17926
rect 3988 17924 4012 17926
rect 4068 17924 4092 17926
rect 4148 17924 4154 17926
rect 3846 17904 4154 17924
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 2880 17436 3188 17456
rect 2880 17434 2886 17436
rect 2942 17434 2966 17436
rect 3022 17434 3046 17436
rect 3102 17434 3126 17436
rect 3182 17434 3188 17436
rect 2942 17382 2944 17434
rect 3124 17382 3126 17434
rect 2880 17380 2886 17382
rect 2942 17380 2966 17382
rect 3022 17380 3046 17382
rect 3102 17380 3126 17382
rect 3182 17380 3188 17382
rect 2880 17360 3188 17380
rect 4264 17338 4292 40831
rect 4356 34678 4384 41262
rect 4434 41168 4490 41177
rect 4434 41103 4490 41112
rect 4344 34672 4396 34678
rect 4344 34614 4396 34620
rect 4342 34504 4398 34513
rect 4342 34439 4398 34448
rect 4356 31890 4384 34439
rect 4344 31884 4396 31890
rect 4344 31826 4396 31832
rect 4344 31792 4396 31798
rect 4344 31734 4396 31740
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1596 16969 1624 17138
rect 1582 16960 1638 16969
rect 1582 16895 1638 16904
rect 1915 16892 2223 16912
rect 1915 16890 1921 16892
rect 1977 16890 2001 16892
rect 2057 16890 2081 16892
rect 2137 16890 2161 16892
rect 2217 16890 2223 16892
rect 1977 16838 1979 16890
rect 2159 16838 2161 16890
rect 1915 16836 1921 16838
rect 1977 16836 2001 16838
rect 2057 16836 2081 16838
rect 2137 16836 2161 16838
rect 2217 16836 2223 16838
rect 1915 16816 2223 16836
rect 3846 16892 4154 16912
rect 3846 16890 3852 16892
rect 3908 16890 3932 16892
rect 3988 16890 4012 16892
rect 4068 16890 4092 16892
rect 4148 16890 4154 16892
rect 3908 16838 3910 16890
rect 4090 16838 4092 16890
rect 3846 16836 3852 16838
rect 3908 16836 3932 16838
rect 3988 16836 4012 16838
rect 4068 16836 4092 16838
rect 4148 16836 4154 16838
rect 3846 16816 4154 16836
rect 4356 16794 4384 31734
rect 4448 25838 4476 41103
rect 4436 25832 4488 25838
rect 4436 25774 4488 25780
rect 4540 24410 4568 41618
rect 4632 36650 4660 41647
rect 4620 36644 4672 36650
rect 4620 36586 4672 36592
rect 4724 36530 4752 41670
rect 4811 41372 5119 41392
rect 4811 41370 4817 41372
rect 4873 41370 4897 41372
rect 4953 41370 4977 41372
rect 5033 41370 5057 41372
rect 5113 41370 5119 41372
rect 4873 41318 4875 41370
rect 5055 41318 5057 41370
rect 4811 41316 4817 41318
rect 4873 41316 4897 41318
rect 4953 41316 4977 41318
rect 5033 41316 5057 41318
rect 5113 41316 5119 41318
rect 4811 41296 5119 41316
rect 5184 41290 5212 41670
rect 5264 41608 5316 41614
rect 5262 41576 5264 41585
rect 5316 41576 5318 41585
rect 5262 41511 5318 41520
rect 5184 41262 5304 41290
rect 4988 41064 5040 41070
rect 4986 41032 4988 41041
rect 5172 41064 5224 41070
rect 5040 41032 5042 41041
rect 5172 41006 5224 41012
rect 4986 40967 5042 40976
rect 4811 40284 5119 40304
rect 4811 40282 4817 40284
rect 4873 40282 4897 40284
rect 4953 40282 4977 40284
rect 5033 40282 5057 40284
rect 5113 40282 5119 40284
rect 4873 40230 4875 40282
rect 5055 40230 5057 40282
rect 4811 40228 4817 40230
rect 4873 40228 4897 40230
rect 4953 40228 4977 40230
rect 5033 40228 5057 40230
rect 5113 40228 5119 40230
rect 4811 40208 5119 40228
rect 4811 39196 5119 39216
rect 4811 39194 4817 39196
rect 4873 39194 4897 39196
rect 4953 39194 4977 39196
rect 5033 39194 5057 39196
rect 5113 39194 5119 39196
rect 4873 39142 4875 39194
rect 5055 39142 5057 39194
rect 4811 39140 4817 39142
rect 4873 39140 4897 39142
rect 4953 39140 4977 39142
rect 5033 39140 5057 39142
rect 5113 39140 5119 39142
rect 4811 39120 5119 39140
rect 5078 38992 5134 39001
rect 5078 38927 5134 38936
rect 5092 38321 5120 38927
rect 5078 38312 5134 38321
rect 5078 38247 5134 38256
rect 4811 38108 5119 38128
rect 4811 38106 4817 38108
rect 4873 38106 4897 38108
rect 4953 38106 4977 38108
rect 5033 38106 5057 38108
rect 5113 38106 5119 38108
rect 4873 38054 4875 38106
rect 5055 38054 5057 38106
rect 4811 38052 4817 38054
rect 4873 38052 4897 38054
rect 4953 38052 4977 38054
rect 5033 38052 5057 38054
rect 5113 38052 5119 38054
rect 4811 38032 5119 38052
rect 4988 37800 5040 37806
rect 4986 37768 4988 37777
rect 5040 37768 5042 37777
rect 4986 37703 5042 37712
rect 4811 37020 5119 37040
rect 4811 37018 4817 37020
rect 4873 37018 4897 37020
rect 4953 37018 4977 37020
rect 5033 37018 5057 37020
rect 5113 37018 5119 37020
rect 4873 36966 4875 37018
rect 5055 36966 5057 37018
rect 4811 36964 4817 36966
rect 4873 36964 4897 36966
rect 4953 36964 4977 36966
rect 5033 36964 5057 36966
rect 5113 36964 5119 36966
rect 4811 36944 5119 36964
rect 4988 36712 5040 36718
rect 4986 36680 4988 36689
rect 5040 36680 5042 36689
rect 4804 36644 4856 36650
rect 4986 36615 5042 36624
rect 4804 36586 4856 36592
rect 4632 36502 4752 36530
rect 4528 24404 4580 24410
rect 4528 24346 4580 24352
rect 4632 24290 4660 36502
rect 4816 36394 4844 36586
rect 4724 36366 4844 36394
rect 4724 26042 4752 36366
rect 4811 35932 5119 35952
rect 4811 35930 4817 35932
rect 4873 35930 4897 35932
rect 4953 35930 4977 35932
rect 5033 35930 5057 35932
rect 5113 35930 5119 35932
rect 4873 35878 4875 35930
rect 5055 35878 5057 35930
rect 4811 35876 4817 35878
rect 4873 35876 4897 35878
rect 4953 35876 4977 35878
rect 5033 35876 5057 35878
rect 5113 35876 5119 35878
rect 4811 35856 5119 35876
rect 5184 35850 5212 41006
rect 5276 37466 5304 41262
rect 5264 37460 5316 37466
rect 5264 37402 5316 37408
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 5276 37097 5304 37266
rect 5262 37088 5318 37097
rect 5262 37023 5318 37032
rect 5264 36168 5316 36174
rect 5264 36110 5316 36116
rect 5276 36009 5304 36110
rect 5262 36000 5318 36009
rect 5262 35935 5318 35944
rect 5184 35822 5304 35850
rect 5172 35760 5224 35766
rect 5172 35702 5224 35708
rect 4988 35624 5040 35630
rect 4986 35592 4988 35601
rect 5040 35592 5042 35601
rect 4986 35527 5042 35536
rect 4811 34844 5119 34864
rect 4811 34842 4817 34844
rect 4873 34842 4897 34844
rect 4953 34842 4977 34844
rect 5033 34842 5057 34844
rect 5113 34842 5119 34844
rect 4873 34790 4875 34842
rect 5055 34790 5057 34842
rect 4811 34788 4817 34790
rect 4873 34788 4897 34790
rect 4953 34788 4977 34790
rect 5033 34788 5057 34790
rect 5113 34788 5119 34790
rect 4811 34768 5119 34788
rect 4988 34536 5040 34542
rect 4986 34504 4988 34513
rect 5040 34504 5042 34513
rect 4986 34439 5042 34448
rect 4811 33756 5119 33776
rect 4811 33754 4817 33756
rect 4873 33754 4897 33756
rect 4953 33754 4977 33756
rect 5033 33754 5057 33756
rect 5113 33754 5119 33756
rect 4873 33702 4875 33754
rect 5055 33702 5057 33754
rect 4811 33700 4817 33702
rect 4873 33700 4897 33702
rect 4953 33700 4977 33702
rect 5033 33700 5057 33702
rect 5113 33700 5119 33702
rect 4811 33680 5119 33700
rect 4988 33448 5040 33454
rect 4988 33390 5040 33396
rect 5000 33017 5028 33390
rect 4986 33008 5042 33017
rect 4986 32943 5042 32952
rect 4811 32668 5119 32688
rect 4811 32666 4817 32668
rect 4873 32666 4897 32668
rect 4953 32666 4977 32668
rect 5033 32666 5057 32668
rect 5113 32666 5119 32668
rect 4873 32614 4875 32666
rect 5055 32614 5057 32666
rect 4811 32612 4817 32614
rect 4873 32612 4897 32614
rect 4953 32612 4977 32614
rect 5033 32612 5057 32614
rect 5113 32612 5119 32614
rect 4811 32592 5119 32612
rect 5184 32450 5212 35702
rect 5276 35222 5304 35822
rect 5264 35216 5316 35222
rect 5264 35158 5316 35164
rect 5264 35080 5316 35086
rect 5264 35022 5316 35028
rect 5276 34785 5304 35022
rect 5262 34776 5318 34785
rect 5262 34711 5318 34720
rect 5264 33992 5316 33998
rect 5264 33934 5316 33940
rect 5276 33697 5304 33934
rect 5262 33688 5318 33697
rect 5368 33658 5396 45766
rect 5460 42362 5488 51046
rect 6368 50720 6420 50726
rect 6366 50688 6368 50697
rect 6420 50688 6422 50697
rect 5776 50620 6084 50640
rect 6366 50623 6422 50632
rect 5776 50618 5782 50620
rect 5838 50618 5862 50620
rect 5918 50618 5942 50620
rect 5998 50618 6022 50620
rect 6078 50618 6084 50620
rect 5838 50566 5840 50618
rect 6020 50566 6022 50618
rect 5776 50564 5782 50566
rect 5838 50564 5862 50566
rect 5918 50564 5942 50566
rect 5998 50564 6022 50566
rect 6078 50564 6084 50566
rect 5776 50544 6084 50564
rect 5540 50312 5592 50318
rect 5540 50254 5592 50260
rect 5552 48346 5580 50254
rect 6000 50176 6052 50182
rect 5998 50144 6000 50153
rect 6052 50144 6054 50153
rect 5998 50079 6054 50088
rect 6184 49632 6236 49638
rect 6184 49574 6236 49580
rect 5776 49532 6084 49552
rect 5776 49530 5782 49532
rect 5838 49530 5862 49532
rect 5918 49530 5942 49532
rect 5998 49530 6022 49532
rect 6078 49530 6084 49532
rect 5838 49478 5840 49530
rect 6020 49478 6022 49530
rect 5776 49476 5782 49478
rect 5838 49476 5862 49478
rect 5918 49476 5942 49478
rect 5998 49476 6022 49478
rect 6078 49476 6084 49478
rect 5776 49456 6084 49476
rect 6196 49473 6224 49574
rect 6182 49464 6238 49473
rect 6182 49399 6238 49408
rect 6000 49088 6052 49094
rect 6000 49030 6052 49036
rect 6012 48929 6040 49030
rect 5998 48920 6054 48929
rect 5998 48855 6054 48864
rect 6184 48544 6236 48550
rect 6184 48486 6236 48492
rect 5776 48444 6084 48464
rect 5776 48442 5782 48444
rect 5838 48442 5862 48444
rect 5918 48442 5942 48444
rect 5998 48442 6022 48444
rect 6078 48442 6084 48444
rect 5838 48390 5840 48442
rect 6020 48390 6022 48442
rect 5776 48388 5782 48390
rect 5838 48388 5862 48390
rect 5918 48388 5942 48390
rect 5998 48388 6022 48390
rect 6078 48388 6084 48390
rect 5776 48368 6084 48388
rect 6196 48385 6224 48486
rect 6182 48376 6238 48385
rect 5540 48340 5592 48346
rect 6182 48311 6238 48320
rect 5540 48282 5592 48288
rect 6000 48000 6052 48006
rect 6000 47942 6052 47948
rect 6012 47841 6040 47942
rect 5998 47832 6054 47841
rect 5998 47767 6054 47776
rect 6184 47456 6236 47462
rect 6184 47398 6236 47404
rect 5776 47356 6084 47376
rect 5776 47354 5782 47356
rect 5838 47354 5862 47356
rect 5918 47354 5942 47356
rect 5998 47354 6022 47356
rect 6078 47354 6084 47356
rect 5838 47302 5840 47354
rect 6020 47302 6022 47354
rect 5776 47300 5782 47302
rect 5838 47300 5862 47302
rect 5918 47300 5942 47302
rect 5998 47300 6022 47302
rect 6078 47300 6084 47302
rect 5776 47280 6084 47300
rect 6196 47297 6224 47398
rect 6182 47288 6238 47297
rect 6182 47223 6238 47232
rect 6000 46912 6052 46918
rect 6000 46854 6052 46860
rect 6012 46753 6040 46854
rect 5998 46744 6054 46753
rect 5998 46679 6054 46688
rect 6276 46572 6328 46578
rect 6276 46514 6328 46520
rect 6184 46368 6236 46374
rect 6184 46310 6236 46316
rect 5776 46268 6084 46288
rect 5776 46266 5782 46268
rect 5838 46266 5862 46268
rect 5918 46266 5942 46268
rect 5998 46266 6022 46268
rect 6078 46266 6084 46268
rect 5838 46214 5840 46266
rect 6020 46214 6022 46266
rect 5776 46212 5782 46214
rect 5838 46212 5862 46214
rect 5918 46212 5942 46214
rect 5998 46212 6022 46214
rect 6078 46212 6084 46214
rect 5776 46192 6084 46212
rect 6196 46073 6224 46310
rect 6182 46064 6238 46073
rect 6182 45999 6238 46008
rect 5816 45960 5868 45966
rect 5816 45902 5868 45908
rect 5828 45393 5856 45902
rect 6000 45824 6052 45830
rect 6000 45766 6052 45772
rect 6012 45529 6040 45766
rect 5998 45520 6054 45529
rect 5998 45455 6054 45464
rect 5814 45384 5870 45393
rect 5814 45319 5870 45328
rect 6184 45280 6236 45286
rect 6184 45222 6236 45228
rect 5776 45180 6084 45200
rect 5776 45178 5782 45180
rect 5838 45178 5862 45180
rect 5918 45178 5942 45180
rect 5998 45178 6022 45180
rect 6078 45178 6084 45180
rect 5838 45126 5840 45178
rect 6020 45126 6022 45178
rect 5776 45124 5782 45126
rect 5838 45124 5862 45126
rect 5918 45124 5942 45126
rect 5998 45124 6022 45126
rect 6078 45124 6084 45126
rect 5776 45104 6084 45124
rect 6196 44985 6224 45222
rect 6182 44976 6238 44985
rect 6182 44911 6238 44920
rect 6000 44736 6052 44742
rect 6000 44678 6052 44684
rect 6012 44441 6040 44678
rect 5998 44432 6054 44441
rect 5540 44396 5592 44402
rect 5998 44367 6054 44376
rect 5540 44338 5592 44344
rect 5552 42650 5580 44338
rect 5632 44192 5684 44198
rect 5632 44134 5684 44140
rect 5644 43897 5672 44134
rect 5776 44092 6084 44112
rect 5776 44090 5782 44092
rect 5838 44090 5862 44092
rect 5918 44090 5942 44092
rect 5998 44090 6022 44092
rect 6078 44090 6084 44092
rect 5838 44038 5840 44090
rect 6020 44038 6022 44090
rect 5776 44036 5782 44038
rect 5838 44036 5862 44038
rect 5918 44036 5942 44038
rect 5998 44036 6022 44038
rect 6078 44036 6084 44038
rect 5776 44016 6084 44036
rect 6288 44010 6316 46514
rect 6196 43982 6316 44010
rect 5630 43888 5686 43897
rect 5630 43823 5686 43832
rect 6000 43648 6052 43654
rect 6000 43590 6052 43596
rect 6012 43353 6040 43590
rect 5998 43344 6054 43353
rect 5998 43279 6054 43288
rect 5632 43104 5684 43110
rect 5632 43046 5684 43052
rect 5644 42809 5672 43046
rect 5776 43004 6084 43024
rect 5776 43002 5782 43004
rect 5838 43002 5862 43004
rect 5918 43002 5942 43004
rect 5998 43002 6022 43004
rect 6078 43002 6084 43004
rect 5838 42950 5840 43002
rect 6020 42950 6022 43002
rect 5776 42948 5782 42950
rect 5838 42948 5862 42950
rect 5918 42948 5942 42950
rect 5998 42948 6022 42950
rect 6078 42948 6084 42950
rect 5776 42928 6084 42948
rect 5630 42800 5686 42809
rect 5630 42735 5686 42744
rect 5552 42622 5672 42650
rect 5448 42356 5500 42362
rect 5448 42298 5500 42304
rect 5448 42220 5500 42226
rect 5448 42162 5500 42168
rect 5460 42022 5488 42162
rect 5448 42016 5500 42022
rect 5448 41958 5500 41964
rect 5262 33623 5318 33632
rect 5356 33652 5408 33658
rect 5356 33594 5408 33600
rect 5264 32904 5316 32910
rect 5264 32846 5316 32852
rect 5276 32609 5304 32846
rect 5262 32600 5318 32609
rect 5262 32535 5318 32544
rect 5184 32422 5304 32450
rect 4988 32360 5040 32366
rect 4988 32302 5040 32308
rect 5172 32360 5224 32366
rect 5172 32302 5224 32308
rect 5000 31929 5028 32302
rect 4986 31920 5042 31929
rect 4986 31855 5042 31864
rect 4811 31580 5119 31600
rect 4811 31578 4817 31580
rect 4873 31578 4897 31580
rect 4953 31578 4977 31580
rect 5033 31578 5057 31580
rect 5113 31578 5119 31580
rect 4873 31526 4875 31578
rect 5055 31526 5057 31578
rect 4811 31524 4817 31526
rect 4873 31524 4897 31526
rect 4953 31524 4977 31526
rect 5033 31524 5057 31526
rect 5113 31524 5119 31526
rect 4811 31504 5119 31524
rect 5184 30954 5212 32302
rect 5092 30926 5212 30954
rect 5276 30938 5304 32422
rect 5460 32366 5488 41958
rect 5540 41472 5592 41478
rect 5540 41414 5592 41420
rect 5552 40186 5580 41414
rect 5540 40180 5592 40186
rect 5540 40122 5592 40128
rect 5644 40066 5672 42622
rect 5722 42120 5778 42129
rect 5722 42055 5724 42064
rect 5776 42055 5778 42064
rect 5724 42026 5776 42032
rect 5776 41916 6084 41936
rect 5776 41914 5782 41916
rect 5838 41914 5862 41916
rect 5918 41914 5942 41916
rect 5998 41914 6022 41916
rect 6078 41914 6084 41916
rect 5838 41862 5840 41914
rect 6020 41862 6022 41914
rect 5776 41860 5782 41862
rect 5838 41860 5862 41862
rect 5918 41860 5942 41862
rect 5998 41860 6022 41862
rect 6078 41860 6084 41862
rect 5776 41840 6084 41860
rect 5776 40828 6084 40848
rect 5776 40826 5782 40828
rect 5838 40826 5862 40828
rect 5918 40826 5942 40828
rect 5998 40826 6022 40828
rect 6078 40826 6084 40828
rect 5838 40774 5840 40826
rect 6020 40774 6022 40826
rect 5776 40772 5782 40774
rect 5838 40772 5862 40774
rect 5918 40772 5942 40774
rect 5998 40772 6022 40774
rect 6078 40772 6084 40774
rect 5776 40752 6084 40772
rect 5724 40520 5776 40526
rect 5722 40488 5724 40497
rect 5776 40488 5778 40497
rect 5722 40423 5778 40432
rect 5552 40038 5672 40066
rect 5816 40044 5868 40050
rect 5552 36378 5580 40038
rect 5816 39986 5868 39992
rect 5632 39976 5684 39982
rect 5828 39953 5856 39986
rect 5632 39918 5684 39924
rect 5814 39944 5870 39953
rect 5644 39642 5672 39918
rect 5814 39879 5870 39888
rect 5776 39740 6084 39760
rect 5776 39738 5782 39740
rect 5838 39738 5862 39740
rect 5918 39738 5942 39740
rect 5998 39738 6022 39740
rect 6078 39738 6084 39740
rect 5838 39686 5840 39738
rect 6020 39686 6022 39738
rect 5776 39684 5782 39686
rect 5838 39684 5862 39686
rect 5918 39684 5942 39686
rect 5998 39684 6022 39686
rect 6078 39684 6084 39686
rect 5776 39664 6084 39684
rect 5632 39636 5684 39642
rect 5632 39578 5684 39584
rect 6092 39432 6144 39438
rect 6090 39400 6092 39409
rect 6144 39400 6146 39409
rect 6090 39335 6146 39344
rect 6196 39098 6224 43982
rect 6276 43784 6328 43790
rect 6276 43726 6328 43732
rect 6184 39092 6236 39098
rect 6184 39034 6236 39040
rect 6184 38956 6236 38962
rect 6184 38898 6236 38904
rect 6196 38729 6224 38898
rect 6182 38720 6238 38729
rect 5776 38652 6084 38672
rect 6182 38655 6238 38664
rect 5776 38650 5782 38652
rect 5838 38650 5862 38652
rect 5918 38650 5942 38652
rect 5998 38650 6022 38652
rect 6078 38650 6084 38652
rect 5838 38598 5840 38650
rect 6020 38598 6022 38650
rect 5776 38596 5782 38598
rect 5838 38596 5862 38598
rect 5918 38596 5942 38598
rect 5998 38596 6022 38598
rect 6078 38596 6084 38598
rect 5776 38576 6084 38596
rect 5630 38448 5686 38457
rect 5630 38383 5686 38392
rect 5540 36372 5592 36378
rect 5540 36314 5592 36320
rect 5540 35216 5592 35222
rect 5540 35158 5592 35164
rect 5448 32360 5500 32366
rect 5354 32328 5410 32337
rect 5448 32302 5500 32308
rect 5354 32263 5410 32272
rect 5368 32178 5396 32263
rect 5368 32150 5488 32178
rect 5354 31784 5410 31793
rect 5354 31719 5410 31728
rect 5264 30932 5316 30938
rect 5092 30666 5120 30926
rect 5264 30874 5316 30880
rect 5172 30864 5224 30870
rect 5172 30806 5224 30812
rect 5080 30660 5132 30666
rect 5080 30602 5132 30608
rect 4811 30492 5119 30512
rect 4811 30490 4817 30492
rect 4873 30490 4897 30492
rect 4953 30490 4977 30492
rect 5033 30490 5057 30492
rect 5113 30490 5119 30492
rect 4873 30438 4875 30490
rect 5055 30438 5057 30490
rect 4811 30436 4817 30438
rect 4873 30436 4897 30438
rect 4953 30436 4977 30438
rect 5033 30436 5057 30438
rect 5113 30436 5119 30438
rect 4811 30416 5119 30436
rect 4811 29404 5119 29424
rect 4811 29402 4817 29404
rect 4873 29402 4897 29404
rect 4953 29402 4977 29404
rect 5033 29402 5057 29404
rect 5113 29402 5119 29404
rect 4873 29350 4875 29402
rect 5055 29350 5057 29402
rect 4811 29348 4817 29350
rect 4873 29348 4897 29350
rect 4953 29348 4977 29350
rect 5033 29348 5057 29350
rect 5113 29348 5119 29350
rect 4811 29328 5119 29348
rect 4988 29096 5040 29102
rect 4988 29038 5040 29044
rect 5000 28665 5028 29038
rect 5184 28762 5212 30806
rect 5368 30410 5396 31719
rect 5460 30870 5488 32150
rect 5448 30864 5500 30870
rect 5448 30806 5500 30812
rect 5552 30818 5580 35158
rect 5644 32434 5672 38383
rect 6092 38344 6144 38350
rect 6092 38286 6144 38292
rect 6104 38185 6132 38286
rect 6090 38176 6146 38185
rect 6090 38111 6146 38120
rect 5776 37564 6084 37584
rect 5776 37562 5782 37564
rect 5838 37562 5862 37564
rect 5918 37562 5942 37564
rect 5998 37562 6022 37564
rect 6078 37562 6084 37564
rect 5838 37510 5840 37562
rect 6020 37510 6022 37562
rect 5776 37508 5782 37510
rect 5838 37508 5862 37510
rect 5918 37508 5942 37510
rect 5998 37508 6022 37510
rect 6078 37508 6084 37510
rect 5776 37488 6084 37508
rect 5776 36476 6084 36496
rect 5776 36474 5782 36476
rect 5838 36474 5862 36476
rect 5918 36474 5942 36476
rect 5998 36474 6022 36476
rect 6078 36474 6084 36476
rect 5838 36422 5840 36474
rect 6020 36422 6022 36474
rect 5776 36420 5782 36422
rect 5838 36420 5862 36422
rect 5918 36420 5942 36422
rect 5998 36420 6022 36422
rect 6078 36420 6084 36422
rect 5776 36400 6084 36420
rect 5776 35388 6084 35408
rect 5776 35386 5782 35388
rect 5838 35386 5862 35388
rect 5918 35386 5942 35388
rect 5998 35386 6022 35388
rect 6078 35386 6084 35388
rect 5838 35334 5840 35386
rect 6020 35334 6022 35386
rect 5776 35332 5782 35334
rect 5838 35332 5862 35334
rect 5918 35332 5942 35334
rect 5998 35332 6022 35334
rect 6078 35332 6084 35334
rect 5776 35312 6084 35332
rect 5776 34300 6084 34320
rect 5776 34298 5782 34300
rect 5838 34298 5862 34300
rect 5918 34298 5942 34300
rect 5998 34298 6022 34300
rect 6078 34298 6084 34300
rect 5838 34246 5840 34298
rect 6020 34246 6022 34298
rect 5776 34244 5782 34246
rect 5838 34244 5862 34246
rect 5918 34244 5942 34246
rect 5998 34244 6022 34246
rect 6078 34244 6084 34246
rect 5776 34224 6084 34244
rect 5776 33212 6084 33232
rect 5776 33210 5782 33212
rect 5838 33210 5862 33212
rect 5918 33210 5942 33212
rect 5998 33210 6022 33212
rect 6078 33210 6084 33212
rect 5838 33158 5840 33210
rect 6020 33158 6022 33210
rect 5776 33156 5782 33158
rect 5838 33156 5862 33158
rect 5918 33156 5942 33158
rect 5998 33156 6022 33158
rect 6078 33156 6084 33158
rect 5776 33136 6084 33156
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 5776 32124 6084 32144
rect 5776 32122 5782 32124
rect 5838 32122 5862 32124
rect 5918 32122 5942 32124
rect 5998 32122 6022 32124
rect 6078 32122 6084 32124
rect 5838 32070 5840 32122
rect 6020 32070 6022 32122
rect 5776 32068 5782 32070
rect 5838 32068 5862 32070
rect 5918 32068 5942 32070
rect 5998 32068 6022 32070
rect 6078 32068 6084 32070
rect 5776 32048 6084 32068
rect 6184 31340 6236 31346
rect 6184 31282 6236 31288
rect 5776 31036 6084 31056
rect 5776 31034 5782 31036
rect 5838 31034 5862 31036
rect 5918 31034 5942 31036
rect 5998 31034 6022 31036
rect 6078 31034 6084 31036
rect 5838 30982 5840 31034
rect 6020 30982 6022 31034
rect 5776 30980 5782 30982
rect 5838 30980 5862 30982
rect 5918 30980 5942 30982
rect 5998 30980 6022 30982
rect 6078 30980 6084 30982
rect 5776 30960 6084 30980
rect 6196 30841 6224 31282
rect 6182 30832 6238 30841
rect 5552 30790 5672 30818
rect 5448 30728 5500 30734
rect 5448 30670 5500 30676
rect 5276 30382 5396 30410
rect 5276 29782 5304 30382
rect 5460 30297 5488 30670
rect 5540 30660 5592 30666
rect 5540 30602 5592 30608
rect 5446 30288 5502 30297
rect 5356 30252 5408 30258
rect 5446 30223 5502 30232
rect 5356 30194 5408 30200
rect 5264 29776 5316 29782
rect 5264 29718 5316 29724
rect 5264 29640 5316 29646
rect 5264 29582 5316 29588
rect 5276 29209 5304 29582
rect 5368 29306 5396 30194
rect 5552 30138 5580 30602
rect 5460 30110 5580 30138
rect 5356 29300 5408 29306
rect 5356 29242 5408 29248
rect 5262 29200 5318 29209
rect 5460 29186 5488 30110
rect 5262 29135 5318 29144
rect 5368 29158 5488 29186
rect 5264 29028 5316 29034
rect 5264 28970 5316 28976
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 4986 28656 5042 28665
rect 4986 28591 5042 28600
rect 4811 28316 5119 28336
rect 4811 28314 4817 28316
rect 4873 28314 4897 28316
rect 4953 28314 4977 28316
rect 5033 28314 5057 28316
rect 5113 28314 5119 28316
rect 4873 28262 4875 28314
rect 5055 28262 5057 28314
rect 4811 28260 4817 28262
rect 4873 28260 4897 28262
rect 4953 28260 4977 28262
rect 5033 28260 5057 28262
rect 5113 28260 5119 28262
rect 4811 28240 5119 28260
rect 5172 28008 5224 28014
rect 5172 27950 5224 27956
rect 4811 27228 5119 27248
rect 4811 27226 4817 27228
rect 4873 27226 4897 27228
rect 4953 27226 4977 27228
rect 5033 27226 5057 27228
rect 5113 27226 5119 27228
rect 4873 27174 4875 27226
rect 5055 27174 5057 27226
rect 4811 27172 4817 27174
rect 4873 27172 4897 27174
rect 4953 27172 4977 27174
rect 5033 27172 5057 27174
rect 5113 27172 5119 27174
rect 4811 27152 5119 27172
rect 5184 27130 5212 27950
rect 5172 27124 5224 27130
rect 5172 27066 5224 27072
rect 5080 26988 5132 26994
rect 5080 26930 5132 26936
rect 5092 26897 5120 26930
rect 5078 26888 5134 26897
rect 5078 26823 5134 26832
rect 5172 26852 5224 26858
rect 5172 26794 5224 26800
rect 4811 26140 5119 26160
rect 4811 26138 4817 26140
rect 4873 26138 4897 26140
rect 4953 26138 4977 26140
rect 5033 26138 5057 26140
rect 5113 26138 5119 26140
rect 4873 26086 4875 26138
rect 5055 26086 5057 26138
rect 4811 26084 4817 26086
rect 4873 26084 4897 26086
rect 4953 26084 4977 26086
rect 5033 26084 5057 26086
rect 5113 26084 5119 26086
rect 4811 26064 5119 26084
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 4448 24262 4660 24290
rect 4448 22098 4476 24262
rect 4436 22092 4488 22098
rect 4724 22094 4752 25774
rect 5184 25362 5212 26794
rect 5276 26586 5304 28970
rect 5264 26580 5316 26586
rect 5264 26522 5316 26528
rect 5264 26444 5316 26450
rect 5264 26386 5316 26392
rect 5172 25356 5224 25362
rect 5172 25298 5224 25304
rect 5172 25220 5224 25226
rect 5172 25162 5224 25168
rect 4811 25052 5119 25072
rect 4811 25050 4817 25052
rect 4873 25050 4897 25052
rect 4953 25050 4977 25052
rect 5033 25050 5057 25052
rect 5113 25050 5119 25052
rect 4873 24998 4875 25050
rect 5055 24998 5057 25050
rect 4811 24996 4817 24998
rect 4873 24996 4897 24998
rect 4953 24996 4977 24998
rect 5033 24996 5057 24998
rect 5113 24996 5119 24998
rect 4811 24976 5119 24996
rect 4811 23964 5119 23984
rect 4811 23962 4817 23964
rect 4873 23962 4897 23964
rect 4953 23962 4977 23964
rect 5033 23962 5057 23964
rect 5113 23962 5119 23964
rect 4873 23910 4875 23962
rect 5055 23910 5057 23962
rect 4811 23908 4817 23910
rect 4873 23908 4897 23910
rect 4953 23908 4977 23910
rect 5033 23908 5057 23910
rect 5113 23908 5119 23910
rect 4811 23888 5119 23908
rect 5184 23866 5212 25162
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 4811 22876 5119 22896
rect 4811 22874 4817 22876
rect 4873 22874 4897 22876
rect 4953 22874 4977 22876
rect 5033 22874 5057 22876
rect 5113 22874 5119 22876
rect 4873 22822 4875 22874
rect 5055 22822 5057 22874
rect 4811 22820 4817 22822
rect 4873 22820 4897 22822
rect 4953 22820 4977 22822
rect 5033 22820 5057 22822
rect 5113 22820 5119 22822
rect 4811 22800 5119 22820
rect 5184 22778 5212 23666
rect 5276 23254 5304 26386
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5276 22953 5304 23054
rect 5262 22944 5318 22953
rect 5262 22879 5318 22888
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5184 22545 5212 22578
rect 5170 22536 5226 22545
rect 5170 22471 5226 22480
rect 5368 22094 5396 29158
rect 5644 29050 5672 30790
rect 6182 30767 6238 30776
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 5776 29948 6084 29968
rect 5776 29946 5782 29948
rect 5838 29946 5862 29948
rect 5918 29946 5942 29948
rect 5998 29946 6022 29948
rect 6078 29946 6084 29948
rect 5838 29894 5840 29946
rect 6020 29894 6022 29946
rect 5776 29892 5782 29894
rect 5838 29892 5862 29894
rect 5918 29892 5942 29894
rect 5998 29892 6022 29894
rect 6078 29892 6084 29894
rect 5776 29872 6084 29892
rect 6196 29753 6224 30670
rect 6182 29744 6238 29753
rect 6182 29679 6238 29688
rect 5460 29022 5672 29050
rect 5460 26518 5488 29022
rect 5776 28860 6084 28880
rect 5776 28858 5782 28860
rect 5838 28858 5862 28860
rect 5918 28858 5942 28860
rect 5998 28858 6022 28860
rect 6078 28858 6084 28860
rect 5838 28806 5840 28858
rect 6020 28806 6022 28858
rect 5776 28804 5782 28806
rect 5838 28804 5862 28806
rect 5918 28804 5942 28806
rect 5998 28804 6022 28806
rect 6078 28804 6084 28806
rect 5776 28784 6084 28804
rect 6092 28552 6144 28558
rect 6092 28494 6144 28500
rect 6104 27985 6132 28494
rect 6184 28076 6236 28082
rect 6184 28018 6236 28024
rect 6090 27976 6146 27985
rect 6090 27911 6146 27920
rect 5540 27872 5592 27878
rect 5540 27814 5592 27820
rect 5552 27062 5580 27814
rect 5776 27772 6084 27792
rect 5776 27770 5782 27772
rect 5838 27770 5862 27772
rect 5918 27770 5942 27772
rect 5998 27770 6022 27772
rect 6078 27770 6084 27772
rect 5838 27718 5840 27770
rect 6020 27718 6022 27770
rect 5776 27716 5782 27718
rect 5838 27716 5862 27718
rect 5918 27716 5942 27718
rect 5998 27716 6022 27718
rect 6078 27716 6084 27718
rect 5776 27696 6084 27716
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5816 27464 5868 27470
rect 6196 27441 6224 28018
rect 5816 27406 5868 27412
rect 6182 27432 6238 27441
rect 5540 27056 5592 27062
rect 5540 26998 5592 27004
rect 5540 26920 5592 26926
rect 5540 26862 5592 26868
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 5448 26376 5500 26382
rect 5446 26344 5448 26353
rect 5500 26344 5502 26353
rect 5446 26279 5502 26288
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 5460 24290 5488 25298
rect 5552 24682 5580 26862
rect 5540 24676 5592 24682
rect 5540 24618 5592 24624
rect 5460 24262 5580 24290
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5460 24041 5488 24142
rect 5446 24032 5502 24041
rect 5446 23967 5502 23976
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 4436 22034 4488 22040
rect 4632 22066 4752 22094
rect 5276 22066 5396 22094
rect 4528 21956 4580 21962
rect 4528 21898 4580 21904
rect 4540 21146 4568 21898
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4632 17882 4660 22066
rect 4811 21788 5119 21808
rect 4811 21786 4817 21788
rect 4873 21786 4897 21788
rect 4953 21786 4977 21788
rect 5033 21786 5057 21788
rect 5113 21786 5119 21788
rect 4873 21734 4875 21786
rect 5055 21734 5057 21786
rect 4811 21732 4817 21734
rect 4873 21732 4897 21734
rect 4953 21732 4977 21734
rect 5033 21732 5057 21734
rect 5113 21732 5119 21734
rect 4811 21712 5119 21732
rect 5276 21434 5304 22066
rect 5460 21690 5488 23462
rect 5552 23322 5580 24262
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 5644 22778 5672 27406
rect 5828 26858 5856 27406
rect 6182 27367 6238 27376
rect 6288 27010 6316 43726
rect 6368 43308 6420 43314
rect 6368 43250 6420 43256
rect 6196 26982 6316 27010
rect 5816 26852 5868 26858
rect 5816 26794 5868 26800
rect 5776 26684 6084 26704
rect 5776 26682 5782 26684
rect 5838 26682 5862 26684
rect 5918 26682 5942 26684
rect 5998 26682 6022 26684
rect 6078 26682 6084 26684
rect 5838 26630 5840 26682
rect 6020 26630 6022 26682
rect 5776 26628 5782 26630
rect 5838 26628 5862 26630
rect 5918 26628 5942 26630
rect 5998 26628 6022 26630
rect 6078 26628 6084 26630
rect 5776 26608 6084 26628
rect 6196 26586 6224 26982
rect 6380 26874 6408 43250
rect 6472 27538 6500 52430
rect 6644 48136 6696 48142
rect 6644 48078 6696 48084
rect 6552 47524 6604 47530
rect 6552 47466 6604 47472
rect 6564 41070 6592 47466
rect 6552 41064 6604 41070
rect 6552 41006 6604 41012
rect 6656 36530 6684 48078
rect 7748 46776 7800 46782
rect 7748 46718 7800 46724
rect 6828 44872 6880 44878
rect 6828 44814 6880 44820
rect 6736 39092 6788 39098
rect 6736 39034 6788 39040
rect 6564 36502 6684 36530
rect 6460 27532 6512 27538
rect 6460 27474 6512 27480
rect 6288 26846 6408 26874
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 5776 25596 6084 25616
rect 5776 25594 5782 25596
rect 5838 25594 5862 25596
rect 5918 25594 5942 25596
rect 5998 25594 6022 25596
rect 6078 25594 6084 25596
rect 5838 25542 5840 25594
rect 6020 25542 6022 25594
rect 5776 25540 5782 25542
rect 5838 25540 5862 25542
rect 5918 25540 5942 25542
rect 5998 25540 6022 25542
rect 6078 25540 6084 25542
rect 5776 25520 6084 25540
rect 6092 25288 6144 25294
rect 6090 25256 6092 25265
rect 6144 25256 6146 25265
rect 6090 25191 6146 25200
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 6196 24585 6224 24754
rect 6182 24576 6238 24585
rect 5776 24508 6084 24528
rect 6182 24511 6238 24520
rect 5776 24506 5782 24508
rect 5838 24506 5862 24508
rect 5918 24506 5942 24508
rect 5998 24506 6022 24508
rect 6078 24506 6084 24508
rect 5838 24454 5840 24506
rect 6020 24454 6022 24506
rect 5776 24452 5782 24454
rect 5838 24452 5862 24454
rect 5918 24452 5942 24454
rect 5998 24452 6022 24454
rect 6078 24452 6084 24454
rect 5776 24432 6084 24452
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 6196 23497 6224 24142
rect 6182 23488 6238 23497
rect 5776 23420 6084 23440
rect 6182 23423 6238 23432
rect 5776 23418 5782 23420
rect 5838 23418 5862 23420
rect 5918 23418 5942 23420
rect 5998 23418 6022 23420
rect 6078 23418 6084 23420
rect 5838 23366 5840 23418
rect 6020 23366 6022 23418
rect 5776 23364 5782 23366
rect 5838 23364 5862 23366
rect 5918 23364 5942 23366
rect 5998 23364 6022 23366
rect 6078 23364 6084 23366
rect 5776 23344 6084 23364
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 6184 22636 6236 22642
rect 6184 22578 6236 22584
rect 5776 22332 6084 22352
rect 5776 22330 5782 22332
rect 5838 22330 5862 22332
rect 5918 22330 5942 22332
rect 5998 22330 6022 22332
rect 6078 22330 6084 22332
rect 5838 22278 5840 22330
rect 6020 22278 6022 22330
rect 5776 22276 5782 22278
rect 5838 22276 5862 22278
rect 5918 22276 5942 22278
rect 5998 22276 6022 22278
rect 6078 22276 6084 22278
rect 5776 22256 6084 22276
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5184 21406 5304 21434
rect 4811 20700 5119 20720
rect 4811 20698 4817 20700
rect 4873 20698 4897 20700
rect 4953 20698 4977 20700
rect 5033 20698 5057 20700
rect 5113 20698 5119 20700
rect 4873 20646 4875 20698
rect 5055 20646 5057 20698
rect 4811 20644 4817 20646
rect 4873 20644 4897 20646
rect 4953 20644 4977 20646
rect 5033 20644 5057 20646
rect 5113 20644 5119 20646
rect 4811 20624 5119 20644
rect 4811 19612 5119 19632
rect 4811 19610 4817 19612
rect 4873 19610 4897 19612
rect 4953 19610 4977 19612
rect 5033 19610 5057 19612
rect 5113 19610 5119 19612
rect 4873 19558 4875 19610
rect 5055 19558 5057 19610
rect 4811 19556 4817 19558
rect 4873 19556 4897 19558
rect 4953 19556 4977 19558
rect 5033 19556 5057 19558
rect 5113 19556 5119 19558
rect 4811 19536 5119 19556
rect 4811 18524 5119 18544
rect 4811 18522 4817 18524
rect 4873 18522 4897 18524
rect 4953 18522 4977 18524
rect 5033 18522 5057 18524
rect 5113 18522 5119 18524
rect 4873 18470 4875 18522
rect 5055 18470 5057 18522
rect 4811 18468 4817 18470
rect 4873 18468 4897 18470
rect 4953 18468 4977 18470
rect 5033 18468 5057 18470
rect 5113 18468 5119 18470
rect 4811 18448 5119 18468
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4528 17604 4580 17610
rect 4528 17546 4580 17552
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1596 16289 1624 16526
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 2880 16348 3188 16368
rect 2880 16346 2886 16348
rect 2942 16346 2966 16348
rect 3022 16346 3046 16348
rect 3102 16346 3126 16348
rect 3182 16346 3188 16348
rect 2942 16294 2944 16346
rect 3124 16294 3126 16346
rect 2880 16292 2886 16294
rect 2942 16292 2966 16294
rect 3022 16292 3046 16294
rect 3102 16292 3126 16294
rect 3182 16292 3188 16294
rect 1582 16280 1638 16289
rect 2880 16272 3188 16292
rect 1582 16215 1638 16224
rect 1915 15804 2223 15824
rect 1915 15802 1921 15804
rect 1977 15802 2001 15804
rect 2057 15802 2081 15804
rect 2137 15802 2161 15804
rect 2217 15802 2223 15804
rect 1977 15750 1979 15802
rect 2159 15750 2161 15802
rect 1915 15748 1921 15750
rect 1977 15748 2001 15750
rect 2057 15748 2081 15750
rect 2137 15748 2161 15750
rect 2217 15748 2223 15750
rect 1915 15728 2223 15748
rect 3846 15804 4154 15824
rect 3846 15802 3852 15804
rect 3908 15802 3932 15804
rect 3988 15802 4012 15804
rect 4068 15802 4092 15804
rect 4148 15802 4154 15804
rect 3908 15750 3910 15802
rect 4090 15750 4092 15802
rect 3846 15748 3852 15750
rect 3908 15748 3932 15750
rect 3988 15748 4012 15750
rect 4068 15748 4092 15750
rect 4148 15748 4154 15750
rect 3846 15728 4154 15748
rect 1584 15496 1636 15502
rect 1582 15464 1584 15473
rect 1636 15464 1638 15473
rect 1582 15399 1638 15408
rect 2880 15260 3188 15280
rect 2880 15258 2886 15260
rect 2942 15258 2966 15260
rect 3022 15258 3046 15260
rect 3102 15258 3126 15260
rect 3182 15258 3188 15260
rect 2942 15206 2944 15258
rect 3124 15206 3126 15258
rect 2880 15204 2886 15206
rect 2942 15204 2966 15206
rect 3022 15204 3046 15206
rect 3102 15204 3126 15206
rect 3182 15204 3188 15206
rect 2880 15184 3188 15204
rect 4264 15162 4292 16458
rect 4448 16454 4476 17138
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 14793 1624 14962
rect 1582 14784 1638 14793
rect 1582 14719 1638 14728
rect 1915 14716 2223 14736
rect 1915 14714 1921 14716
rect 1977 14714 2001 14716
rect 2057 14714 2081 14716
rect 2137 14714 2161 14716
rect 2217 14714 2223 14716
rect 1977 14662 1979 14714
rect 2159 14662 2161 14714
rect 1915 14660 1921 14662
rect 1977 14660 2001 14662
rect 2057 14660 2081 14662
rect 2137 14660 2161 14662
rect 2217 14660 2223 14662
rect 1915 14640 2223 14660
rect 3846 14716 4154 14736
rect 3846 14714 3852 14716
rect 3908 14714 3932 14716
rect 3988 14714 4012 14716
rect 4068 14714 4092 14716
rect 4148 14714 4154 14716
rect 3908 14662 3910 14714
rect 4090 14662 4092 14714
rect 3846 14660 3852 14662
rect 3908 14660 3932 14662
rect 3988 14660 4012 14662
rect 4068 14660 4092 14662
rect 4148 14660 4154 14662
rect 3846 14640 4154 14660
rect 4356 14618 4384 16050
rect 4540 15706 4568 17546
rect 4811 17436 5119 17456
rect 4811 17434 4817 17436
rect 4873 17434 4897 17436
rect 4953 17434 4977 17436
rect 5033 17434 5057 17436
rect 5113 17434 5119 17436
rect 4873 17382 4875 17434
rect 5055 17382 5057 17434
rect 4811 17380 4817 17382
rect 4873 17380 4897 17382
rect 4953 17380 4977 17382
rect 5033 17380 5057 17382
rect 5113 17380 5119 17382
rect 4811 17360 5119 17380
rect 4811 16348 5119 16368
rect 4811 16346 4817 16348
rect 4873 16346 4897 16348
rect 4953 16346 4977 16348
rect 5033 16346 5057 16348
rect 5113 16346 5119 16348
rect 4873 16294 4875 16346
rect 5055 16294 5057 16346
rect 4811 16292 4817 16294
rect 4873 16292 4897 16294
rect 4953 16292 4977 16294
rect 5033 16292 5057 16294
rect 5113 16292 5119 16294
rect 4811 16272 5119 16292
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4811 15260 5119 15280
rect 4811 15258 4817 15260
rect 4873 15258 4897 15260
rect 4953 15258 4977 15260
rect 5033 15258 5057 15260
rect 5113 15258 5119 15260
rect 4873 15206 4875 15258
rect 5055 15206 5057 15258
rect 4811 15204 4817 15206
rect 4873 15204 4897 15206
rect 4953 15204 4977 15206
rect 5033 15204 5057 15206
rect 5113 15204 5119 15206
rect 4811 15184 5119 15204
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13977 1624 14350
rect 2880 14172 3188 14192
rect 2880 14170 2886 14172
rect 2942 14170 2966 14172
rect 3022 14170 3046 14172
rect 3102 14170 3126 14172
rect 3182 14170 3188 14172
rect 2942 14118 2944 14170
rect 3124 14118 3126 14170
rect 2880 14116 2886 14118
rect 2942 14116 2966 14118
rect 3022 14116 3046 14118
rect 3102 14116 3126 14118
rect 3182 14116 3188 14118
rect 2880 14096 3188 14116
rect 4811 14172 5119 14192
rect 4811 14170 4817 14172
rect 4873 14170 4897 14172
rect 4953 14170 4977 14172
rect 5033 14170 5057 14172
rect 5113 14170 5119 14172
rect 4873 14118 4875 14170
rect 5055 14118 5057 14170
rect 4811 14116 4817 14118
rect 4873 14116 4897 14118
rect 4953 14116 4977 14118
rect 5033 14116 5057 14118
rect 5113 14116 5119 14118
rect 4811 14096 5119 14116
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 1915 13628 2223 13648
rect 1915 13626 1921 13628
rect 1977 13626 2001 13628
rect 2057 13626 2081 13628
rect 2137 13626 2161 13628
rect 2217 13626 2223 13628
rect 1977 13574 1979 13626
rect 2159 13574 2161 13626
rect 1915 13572 1921 13574
rect 1977 13572 2001 13574
rect 2057 13572 2081 13574
rect 2137 13572 2161 13574
rect 2217 13572 2223 13574
rect 1915 13552 2223 13572
rect 3160 13530 3188 13874
rect 3846 13628 4154 13648
rect 3846 13626 3852 13628
rect 3908 13626 3932 13628
rect 3988 13626 4012 13628
rect 4068 13626 4092 13628
rect 4148 13626 4154 13628
rect 3908 13574 3910 13626
rect 4090 13574 4092 13626
rect 3846 13572 3852 13574
rect 3908 13572 3932 13574
rect 3988 13572 4012 13574
rect 4068 13572 4092 13574
rect 4148 13572 4154 13574
rect 3846 13552 4154 13572
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1412 12986 1440 13194
rect 1596 13161 1624 13262
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 2880 13084 3188 13104
rect 2880 13082 2886 13084
rect 2942 13082 2966 13084
rect 3022 13082 3046 13084
rect 3102 13082 3126 13084
rect 3182 13082 3188 13084
rect 2942 13030 2944 13082
rect 3124 13030 3126 13082
rect 2880 13028 2886 13030
rect 2942 13028 2966 13030
rect 3022 13028 3046 13030
rect 3102 13028 3126 13030
rect 3182 13028 3188 13030
rect 2880 13008 3188 13028
rect 4811 13084 5119 13104
rect 4811 13082 4817 13084
rect 4873 13082 4897 13084
rect 4953 13082 4977 13084
rect 5033 13082 5057 13084
rect 5113 13082 5119 13084
rect 4873 13030 4875 13082
rect 5055 13030 5057 13082
rect 4811 13028 4817 13030
rect 4873 13028 4897 13030
rect 4953 13028 4977 13030
rect 5033 13028 5057 13030
rect 5113 13028 5119 13030
rect 4811 13008 5119 13028
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 5184 12918 5212 21406
rect 5552 19514 5580 22170
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5644 20602 5672 21898
rect 6196 21865 6224 22578
rect 6182 21856 6238 21865
rect 6182 21791 6238 21800
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 5776 21244 6084 21264
rect 5776 21242 5782 21244
rect 5838 21242 5862 21244
rect 5918 21242 5942 21244
rect 5998 21242 6022 21244
rect 6078 21242 6084 21244
rect 5838 21190 5840 21242
rect 6020 21190 6022 21242
rect 5776 21188 5782 21190
rect 5838 21188 5862 21190
rect 5918 21188 5942 21190
rect 5998 21188 6022 21190
rect 6078 21188 6084 21190
rect 5776 21168 6084 21188
rect 6196 21185 6224 21490
rect 6182 21176 6238 21185
rect 6182 21111 6238 21120
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 6104 20641 6132 20878
rect 6090 20632 6146 20641
rect 5632 20596 5684 20602
rect 6090 20567 6146 20576
rect 5632 20538 5684 20544
rect 6184 20460 6236 20466
rect 6184 20402 6236 20408
rect 5776 20156 6084 20176
rect 5776 20154 5782 20156
rect 5838 20154 5862 20156
rect 5918 20154 5942 20156
rect 5998 20154 6022 20156
rect 6078 20154 6084 20156
rect 5838 20102 5840 20154
rect 6020 20102 6022 20154
rect 5776 20100 5782 20102
rect 5838 20100 5862 20102
rect 5918 20100 5942 20102
rect 5998 20100 6022 20102
rect 6078 20100 6084 20102
rect 5776 20080 6084 20100
rect 6196 20097 6224 20402
rect 6182 20088 6238 20097
rect 6182 20023 6238 20032
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6104 19553 6132 19790
rect 6090 19544 6146 19553
rect 5540 19508 5592 19514
rect 6090 19479 6146 19488
rect 5540 19450 5592 19456
rect 5776 19068 6084 19088
rect 5776 19066 5782 19068
rect 5838 19066 5862 19068
rect 5918 19066 5942 19068
rect 5998 19066 6022 19068
rect 6078 19066 6084 19068
rect 5838 19014 5840 19066
rect 6020 19014 6022 19066
rect 5776 19012 5782 19014
rect 5838 19012 5862 19014
rect 5918 19012 5942 19014
rect 5998 19012 6022 19014
rect 6078 19012 6084 19014
rect 5776 18992 6084 19012
rect 6288 18850 6316 26846
rect 6564 26738 6592 36502
rect 6644 36372 6696 36378
rect 6644 36314 6696 36320
rect 6380 26710 6592 26738
rect 6380 19242 6408 26710
rect 6552 26580 6604 26586
rect 6552 26522 6604 26528
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6472 22234 6500 23258
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6472 19009 6500 19246
rect 6458 19000 6514 19009
rect 6458 18935 6514 18944
rect 6288 18822 6500 18850
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6104 18465 6132 18702
rect 6090 18456 6146 18465
rect 6090 18391 6146 18400
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5460 17241 5488 17614
rect 5446 17232 5502 17241
rect 5446 17167 5502 17176
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5276 15706 5304 16526
rect 5552 16522 5580 18022
rect 5776 17980 6084 18000
rect 5776 17978 5782 17980
rect 5838 17978 5862 17980
rect 5918 17978 5942 17980
rect 5998 17978 6022 17980
rect 6078 17978 6084 17980
rect 5838 17926 5840 17978
rect 6020 17926 6022 17978
rect 5776 17924 5782 17926
rect 5838 17924 5862 17926
rect 5918 17924 5942 17926
rect 5998 17924 6022 17926
rect 6078 17924 6084 17926
rect 5776 17904 6084 17924
rect 6196 17785 6224 18226
rect 6182 17776 6238 17785
rect 6182 17711 6238 17720
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5644 16658 5672 16934
rect 5776 16892 6084 16912
rect 5776 16890 5782 16892
rect 5838 16890 5862 16892
rect 5918 16890 5942 16892
rect 5998 16890 6022 16892
rect 6078 16890 6084 16892
rect 5838 16838 5840 16890
rect 6020 16838 6022 16890
rect 5776 16836 5782 16838
rect 5838 16836 5862 16838
rect 5918 16836 5942 16838
rect 5998 16836 6022 16838
rect 6078 16836 6084 16838
rect 5776 16816 6084 16836
rect 5816 16720 5868 16726
rect 6196 16697 6224 17614
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 5816 16662 5868 16668
rect 6182 16688 6238 16697
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5828 16250 5856 16662
rect 6182 16623 6238 16632
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 15065 5488 15438
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5446 15056 5502 15065
rect 5356 15020 5408 15026
rect 5446 14991 5502 15000
rect 5356 14962 5408 14968
rect 5368 14550 5396 14962
rect 5552 14618 5580 15302
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5644 14414 5672 15846
rect 5776 15804 6084 15824
rect 5776 15802 5782 15804
rect 5838 15802 5862 15804
rect 5918 15802 5942 15804
rect 5998 15802 6022 15804
rect 6078 15802 6084 15804
rect 5838 15750 5840 15802
rect 6020 15750 6022 15802
rect 5776 15748 5782 15750
rect 5838 15748 5862 15750
rect 5918 15748 5942 15750
rect 5998 15748 6022 15750
rect 6078 15748 6084 15750
rect 5776 15728 6084 15748
rect 6196 15609 6224 16050
rect 6182 15600 6238 15609
rect 6182 15535 6238 15544
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 5776 14716 6084 14736
rect 5776 14714 5782 14716
rect 5838 14714 5862 14716
rect 5918 14714 5942 14716
rect 5998 14714 6022 14716
rect 6078 14714 6084 14716
rect 5838 14662 5840 14714
rect 6020 14662 6022 14714
rect 5776 14660 5782 14662
rect 5838 14660 5862 14662
rect 5918 14660 5942 14662
rect 5998 14660 6022 14662
rect 6078 14660 6084 14662
rect 5776 14640 6084 14660
rect 6196 14521 6224 15438
rect 6288 14958 6316 16390
rect 6380 16153 6408 17138
rect 6366 16144 6422 16153
rect 6366 16079 6422 16088
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6182 14512 6238 14521
rect 6182 14447 6238 14456
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 1596 12481 1624 12786
rect 1915 12540 2223 12560
rect 1915 12538 1921 12540
rect 1977 12538 2001 12540
rect 2057 12538 2081 12540
rect 2137 12538 2161 12540
rect 2217 12538 2223 12540
rect 1977 12486 1979 12538
rect 2159 12486 2161 12538
rect 1915 12484 1921 12486
rect 1977 12484 2001 12486
rect 2057 12484 2081 12486
rect 2137 12484 2161 12486
rect 2217 12484 2223 12486
rect 1582 12472 1638 12481
rect 1915 12464 2223 12484
rect 3846 12540 4154 12560
rect 3846 12538 3852 12540
rect 3908 12538 3932 12540
rect 3988 12538 4012 12540
rect 4068 12538 4092 12540
rect 4148 12538 4154 12540
rect 3908 12486 3910 12538
rect 4090 12486 4092 12538
rect 3846 12484 3852 12486
rect 3908 12484 3932 12486
rect 3988 12484 4012 12486
rect 4068 12484 4092 12486
rect 4148 12484 4154 12486
rect 3846 12464 4154 12484
rect 1582 12407 1638 12416
rect 2880 11996 3188 12016
rect 2880 11994 2886 11996
rect 2942 11994 2966 11996
rect 3022 11994 3046 11996
rect 3102 11994 3126 11996
rect 3182 11994 3188 11996
rect 2942 11942 2944 11994
rect 3124 11942 3126 11994
rect 2880 11940 2886 11942
rect 2942 11940 2966 11942
rect 3022 11940 3046 11942
rect 3102 11940 3126 11942
rect 3182 11940 3188 11942
rect 2880 11920 3188 11940
rect 4264 11898 4292 12786
rect 4811 11996 5119 12016
rect 4811 11994 4817 11996
rect 4873 11994 4897 11996
rect 4953 11994 4977 11996
rect 5033 11994 5057 11996
rect 5113 11994 5119 11996
rect 4873 11942 4875 11994
rect 5055 11942 5057 11994
rect 4811 11940 4817 11942
rect 4873 11940 4897 11942
rect 4953 11940 4977 11942
rect 5033 11940 5057 11942
rect 5113 11940 5119 11942
rect 4811 11920 5119 11940
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 5552 11830 5580 13126
rect 5644 12986 5672 14214
rect 5828 14074 5856 14350
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5828 13841 5856 13874
rect 5814 13832 5870 13841
rect 5814 13767 5870 13776
rect 5776 13628 6084 13648
rect 5776 13626 5782 13628
rect 5838 13626 5862 13628
rect 5918 13626 5942 13628
rect 5998 13626 6022 13628
rect 6078 13626 6084 13628
rect 5838 13574 5840 13626
rect 6020 13574 6022 13626
rect 5776 13572 5782 13574
rect 5838 13572 5862 13574
rect 5918 13572 5942 13574
rect 5998 13572 6022 13574
rect 6078 13572 6084 13574
rect 5776 13552 6084 13572
rect 6472 13462 6500 18822
rect 6564 14006 6592 26522
rect 6656 16726 6684 36314
rect 6748 19990 6776 39034
rect 6840 31890 6868 44814
rect 7472 42288 7524 42294
rect 7472 42230 7524 42236
rect 7484 41432 7512 42230
rect 7656 41540 7708 41546
rect 7656 41482 7708 41488
rect 7472 41426 7524 41432
rect 7472 41368 7524 41374
rect 7668 41206 7696 41482
rect 7656 41200 7708 41206
rect 7656 41142 7708 41148
rect 7760 40458 7788 46718
rect 7932 41404 7984 41410
rect 7932 41346 7984 41352
rect 7748 40452 7800 40458
rect 7748 40394 7800 40400
rect 7944 36514 7972 41346
rect 7932 36508 7984 36514
rect 7932 36450 7984 36456
rect 6828 31884 6880 31890
rect 6828 31826 6880 31832
rect 6828 31748 6880 31754
rect 6828 31690 6880 31696
rect 6840 31385 6868 31690
rect 6826 31376 6882 31385
rect 6826 31311 6882 31320
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6840 25809 6868 26182
rect 6826 25800 6882 25809
rect 6826 25735 6882 25744
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6840 23118 6868 23462
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6092 13320 6144 13326
rect 6090 13288 6092 13297
rect 6144 13288 6146 13297
rect 6090 13223 6146 13232
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12753 5856 12786
rect 5814 12744 5870 12753
rect 5814 12679 5870 12688
rect 5776 12540 6084 12560
rect 5776 12538 5782 12540
rect 5838 12538 5862 12540
rect 5918 12538 5942 12540
rect 5998 12538 6022 12540
rect 6078 12538 6084 12540
rect 5838 12486 5840 12538
rect 6020 12486 6022 12538
rect 5776 12484 5782 12486
rect 5838 12484 5862 12486
rect 5918 12484 5942 12486
rect 5998 12484 6022 12486
rect 6078 12484 6084 12486
rect 5776 12464 6084 12484
rect 6092 12232 6144 12238
rect 6090 12200 6092 12209
rect 6144 12200 6146 12209
rect 6090 12135 6146 12144
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 1596 11665 1624 11698
rect 1582 11656 1638 11665
rect 1582 11591 1638 11600
rect 1915 11452 2223 11472
rect 1915 11450 1921 11452
rect 1977 11450 2001 11452
rect 2057 11450 2081 11452
rect 2137 11450 2161 11452
rect 2217 11450 2223 11452
rect 1977 11398 1979 11450
rect 2159 11398 2161 11450
rect 1915 11396 1921 11398
rect 1977 11396 2001 11398
rect 2057 11396 2081 11398
rect 2137 11396 2161 11398
rect 2217 11396 2223 11398
rect 1915 11376 2223 11396
rect 3846 11452 4154 11472
rect 3846 11450 3852 11452
rect 3908 11450 3932 11452
rect 3988 11450 4012 11452
rect 4068 11450 4092 11452
rect 4148 11450 4154 11452
rect 3908 11398 3910 11450
rect 4090 11398 4092 11450
rect 3846 11396 3852 11398
rect 3908 11396 3932 11398
rect 3988 11396 4012 11398
rect 4068 11396 4092 11398
rect 4148 11396 4154 11398
rect 3846 11376 4154 11396
rect 5460 11354 5488 11698
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 11354 5580 11630
rect 5644 11558 5672 12038
rect 6182 11656 6238 11665
rect 6182 11591 6238 11600
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5776 11452 6084 11472
rect 5776 11450 5782 11452
rect 5838 11450 5862 11452
rect 5918 11450 5942 11452
rect 5998 11450 6022 11452
rect 6078 11450 6084 11452
rect 5838 11398 5840 11450
rect 6020 11398 6022 11450
rect 5776 11396 5782 11398
rect 5838 11396 5862 11398
rect 5918 11396 5942 11398
rect 5998 11396 6022 11398
rect 6078 11396 6084 11398
rect 5776 11376 6084 11396
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6196 11150 6224 11591
rect 4252 11144 4304 11150
rect 4804 11144 4856 11150
rect 4252 11086 4304 11092
rect 4802 11112 4804 11121
rect 5356 11144 5408 11150
rect 4856 11112 4858 11121
rect 1584 11008 1636 11014
rect 1582 10976 1584 10985
rect 1636 10976 1638 10985
rect 1582 10911 1638 10920
rect 2880 10908 3188 10928
rect 2880 10906 2886 10908
rect 2942 10906 2966 10908
rect 3022 10906 3046 10908
rect 3102 10906 3126 10908
rect 3182 10906 3188 10908
rect 2942 10854 2944 10906
rect 3124 10854 3126 10906
rect 2880 10852 2886 10854
rect 2942 10852 2966 10854
rect 3022 10852 3046 10854
rect 3102 10852 3126 10854
rect 3182 10852 3188 10854
rect 2880 10832 3188 10852
rect 4264 10810 4292 11086
rect 5356 11086 5408 11092
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 4802 11047 4858 11056
rect 4811 10908 5119 10928
rect 4811 10906 4817 10908
rect 4873 10906 4897 10908
rect 4953 10906 4977 10908
rect 5033 10906 5057 10908
rect 5113 10906 5119 10908
rect 4873 10854 4875 10906
rect 5055 10854 5057 10906
rect 4811 10852 4817 10854
rect 4873 10852 4897 10854
rect 4953 10852 4977 10854
rect 5033 10852 5057 10854
rect 5113 10852 5119 10854
rect 4811 10832 5119 10852
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10266 1440 10610
rect 5368 10577 5396 11086
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5354 10568 5410 10577
rect 5354 10503 5410 10512
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1596 10169 1624 10406
rect 1915 10364 2223 10384
rect 1915 10362 1921 10364
rect 1977 10362 2001 10364
rect 2057 10362 2081 10364
rect 2137 10362 2161 10364
rect 2217 10362 2223 10364
rect 1977 10310 1979 10362
rect 2159 10310 2161 10362
rect 1915 10308 1921 10310
rect 1977 10308 2001 10310
rect 2057 10308 2081 10310
rect 2137 10308 2161 10310
rect 2217 10308 2223 10310
rect 1915 10288 2223 10308
rect 3846 10364 4154 10384
rect 3846 10362 3852 10364
rect 3908 10362 3932 10364
rect 3988 10362 4012 10364
rect 4068 10362 4092 10364
rect 4148 10362 4154 10364
rect 3908 10310 3910 10362
rect 4090 10310 4092 10362
rect 3846 10308 3852 10310
rect 3908 10308 3932 10310
rect 3988 10308 4012 10310
rect 4068 10308 4092 10310
rect 4148 10308 4154 10310
rect 3846 10288 4154 10308
rect 1582 10160 1638 10169
rect 1582 10095 1638 10104
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 2880 9820 3188 9840
rect 2880 9818 2886 9820
rect 2942 9818 2966 9820
rect 3022 9818 3046 9820
rect 3102 9818 3126 9820
rect 3182 9818 3188 9820
rect 2942 9766 2944 9818
rect 3124 9766 3126 9818
rect 2880 9764 2886 9766
rect 2942 9764 2966 9766
rect 3022 9764 3046 9766
rect 3102 9764 3126 9766
rect 3182 9764 3188 9766
rect 2880 9744 3188 9764
rect 4811 9820 5119 9840
rect 4811 9818 4817 9820
rect 4873 9818 4897 9820
rect 4953 9818 4977 9820
rect 5033 9818 5057 9820
rect 5113 9818 5119 9820
rect 4873 9766 4875 9818
rect 5055 9766 5057 9818
rect 4811 9764 4817 9766
rect 4873 9764 4897 9766
rect 4953 9764 4977 9766
rect 5033 9764 5057 9766
rect 5113 9764 5119 9766
rect 4811 9744 5119 9764
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9178 1440 9522
rect 5184 9489 5212 9998
rect 5460 9897 5488 10610
rect 5776 10364 6084 10384
rect 5776 10362 5782 10364
rect 5838 10362 5862 10364
rect 5918 10362 5942 10364
rect 5998 10362 6022 10364
rect 6078 10362 6084 10364
rect 5838 10310 5840 10362
rect 6020 10310 6022 10362
rect 5776 10308 5782 10310
rect 5838 10308 5862 10310
rect 5918 10308 5942 10310
rect 5998 10308 6022 10310
rect 6078 10308 6084 10310
rect 5776 10288 6084 10308
rect 5632 9920 5684 9926
rect 5446 9888 5502 9897
rect 5632 9862 5684 9868
rect 5446 9823 5502 9832
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5170 9480 5226 9489
rect 5170 9415 5226 9424
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 4252 9376 4304 9382
rect 1636 9344 1638 9353
rect 4252 9318 4304 9324
rect 1582 9279 1638 9288
rect 1915 9276 2223 9296
rect 1915 9274 1921 9276
rect 1977 9274 2001 9276
rect 2057 9274 2081 9276
rect 2137 9274 2161 9276
rect 2217 9274 2223 9276
rect 1977 9222 1979 9274
rect 2159 9222 2161 9274
rect 1915 9220 1921 9222
rect 1977 9220 2001 9222
rect 2057 9220 2081 9222
rect 2137 9220 2161 9222
rect 2217 9220 2223 9222
rect 1915 9200 2223 9220
rect 3846 9276 4154 9296
rect 3846 9274 3852 9276
rect 3908 9274 3932 9276
rect 3988 9274 4012 9276
rect 4068 9274 4092 9276
rect 4148 9274 4154 9276
rect 3908 9222 3910 9274
rect 4090 9222 4092 9274
rect 3846 9220 3852 9222
rect 3908 9220 3932 9222
rect 3988 9220 4012 9222
rect 4068 9220 4092 9222
rect 4148 9220 4154 9222
rect 3846 9200 4154 9220
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8634 1440 8910
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8673 1624 8774
rect 2880 8732 3188 8752
rect 2880 8730 2886 8732
rect 2942 8730 2966 8732
rect 3022 8730 3046 8732
rect 3102 8730 3126 8732
rect 3182 8730 3188 8732
rect 2942 8678 2944 8730
rect 3124 8678 3126 8730
rect 2880 8676 2886 8678
rect 2942 8676 2966 8678
rect 3022 8676 3046 8678
rect 3102 8676 3126 8678
rect 3182 8676 3188 8678
rect 1582 8664 1638 8673
rect 1400 8628 1452 8634
rect 2880 8656 3188 8676
rect 1582 8599 1638 8608
rect 1400 8570 1452 8576
rect 4264 8498 4292 9318
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 1915 8188 2223 8208
rect 1915 8186 1921 8188
rect 1977 8186 2001 8188
rect 2057 8186 2081 8188
rect 2137 8186 2161 8188
rect 2217 8186 2223 8188
rect 1977 8134 1979 8186
rect 2159 8134 2161 8186
rect 1915 8132 1921 8134
rect 1977 8132 2001 8134
rect 2057 8132 2081 8134
rect 2137 8132 2161 8134
rect 2217 8132 2223 8134
rect 1915 8112 2223 8132
rect 3846 8188 4154 8208
rect 3846 8186 3852 8188
rect 3908 8186 3932 8188
rect 3988 8186 4012 8188
rect 4068 8186 4092 8188
rect 4148 8186 4154 8188
rect 3908 8134 3910 8186
rect 4090 8134 4092 8186
rect 3846 8132 3852 8134
rect 3908 8132 3932 8134
rect 3988 8132 4012 8134
rect 4068 8132 4092 8134
rect 4148 8132 4154 8134
rect 3846 8112 4154 8132
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1582 7848 1638 7857
rect 1412 7546 1440 7822
rect 1582 7783 1638 7792
rect 1596 7750 1624 7783
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 2880 7644 3188 7664
rect 2880 7642 2886 7644
rect 2942 7642 2966 7644
rect 3022 7642 3046 7644
rect 3102 7642 3126 7644
rect 3182 7642 3188 7644
rect 2942 7590 2944 7642
rect 3124 7590 3126 7642
rect 2880 7588 2886 7590
rect 2942 7588 2966 7590
rect 3022 7588 3046 7590
rect 3102 7588 3126 7590
rect 3182 7588 3188 7590
rect 2880 7568 3188 7588
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 1584 7200 1636 7206
rect 1582 7168 1584 7177
rect 1636 7168 1638 7177
rect 1582 7103 1638 7112
rect 1915 7100 2223 7120
rect 1915 7098 1921 7100
rect 1977 7098 2001 7100
rect 2057 7098 2081 7100
rect 2137 7098 2161 7100
rect 2217 7098 2223 7100
rect 1977 7046 1979 7098
rect 2159 7046 2161 7098
rect 1915 7044 1921 7046
rect 1977 7044 2001 7046
rect 2057 7044 2081 7046
rect 2137 7044 2161 7046
rect 2217 7044 2223 7046
rect 1915 7024 2223 7044
rect 3252 7002 3280 7346
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6458 1440 6734
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1596 6361 1624 6598
rect 2880 6556 3188 6576
rect 2880 6554 2886 6556
rect 2942 6554 2966 6556
rect 3022 6554 3046 6556
rect 3102 6554 3126 6556
rect 3182 6554 3188 6556
rect 2942 6502 2944 6554
rect 3124 6502 3126 6554
rect 2880 6500 2886 6502
rect 2942 6500 2966 6502
rect 3022 6500 3046 6502
rect 3102 6500 3126 6502
rect 3182 6500 3188 6502
rect 2880 6480 3188 6500
rect 1582 6352 1638 6361
rect 3712 6322 3740 7142
rect 3846 7100 4154 7120
rect 3846 7098 3852 7100
rect 3908 7098 3932 7100
rect 3988 7098 4012 7100
rect 4068 7098 4092 7100
rect 4148 7098 4154 7100
rect 3908 7046 3910 7098
rect 4090 7046 4092 7098
rect 3846 7044 3852 7046
rect 3908 7044 3932 7046
rect 3988 7044 4012 7046
rect 4068 7044 4092 7046
rect 4148 7044 4154 7046
rect 3846 7024 4154 7044
rect 4264 7002 4292 7346
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4356 6390 4384 7686
rect 4448 7546 4476 8366
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4540 7478 4568 8774
rect 4811 8732 5119 8752
rect 4811 8730 4817 8732
rect 4873 8730 4897 8732
rect 4953 8730 4977 8732
rect 5033 8730 5057 8732
rect 5113 8730 5119 8732
rect 4873 8678 4875 8730
rect 5055 8678 5057 8730
rect 4811 8676 4817 8678
rect 4873 8676 4897 8678
rect 4953 8676 4977 8678
rect 5033 8676 5057 8678
rect 5113 8676 5119 8678
rect 4811 8656 5119 8676
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5276 8090 5304 8434
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4811 7644 5119 7664
rect 4811 7642 4817 7644
rect 4873 7642 4897 7644
rect 4953 7642 4977 7644
rect 5033 7642 5057 7644
rect 5113 7642 5119 7644
rect 4873 7590 4875 7642
rect 5055 7590 5057 7642
rect 4811 7588 4817 7590
rect 4873 7588 4897 7590
rect 4953 7588 4977 7590
rect 5033 7588 5057 7590
rect 5113 7588 5119 7590
rect 4811 7568 5119 7588
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4448 6458 4476 7346
rect 5184 6914 5212 7822
rect 5368 7721 5396 8910
rect 5460 8401 5488 9522
rect 5644 9042 5672 9862
rect 5776 9276 6084 9296
rect 5776 9274 5782 9276
rect 5838 9274 5862 9276
rect 5918 9274 5942 9276
rect 5998 9274 6022 9276
rect 6078 9274 6084 9276
rect 5838 9222 5840 9274
rect 6020 9222 6022 9274
rect 5776 9220 5782 9222
rect 5838 9220 5862 9222
rect 5918 9220 5942 9222
rect 5998 9220 6022 9222
rect 6078 9220 6084 9222
rect 5776 9200 6084 9220
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 6184 8832 6236 8838
rect 6920 8832 6972 8838
rect 6184 8774 6236 8780
rect 6918 8800 6920 8809
rect 6972 8800 6974 8809
rect 5446 8392 5502 8401
rect 5446 8327 5502 8336
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 7886 5488 8230
rect 5776 8188 6084 8208
rect 5776 8186 5782 8188
rect 5838 8186 5862 8188
rect 5918 8186 5942 8188
rect 5998 8186 6022 8188
rect 6078 8186 6084 8188
rect 5838 8134 5840 8186
rect 6020 8134 6022 8186
rect 5776 8132 5782 8134
rect 5838 8132 5862 8134
rect 5918 8132 5942 8134
rect 5998 8132 6022 8134
rect 6078 8132 6084 8134
rect 5776 8112 6084 8132
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5354 7712 5410 7721
rect 5354 7647 5410 7656
rect 5460 7410 5488 7822
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5184 6886 5304 6914
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 1582 6287 1638 6296
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 1915 6012 2223 6032
rect 1915 6010 1921 6012
rect 1977 6010 2001 6012
rect 2057 6010 2081 6012
rect 2137 6010 2161 6012
rect 2217 6010 2223 6012
rect 1977 5958 1979 6010
rect 2159 5958 2161 6010
rect 1915 5956 1921 5958
rect 1977 5956 2001 5958
rect 2057 5956 2081 5958
rect 2137 5956 2161 5958
rect 2217 5956 2223 5958
rect 1915 5936 2223 5956
rect 3846 6012 4154 6032
rect 3846 6010 3852 6012
rect 3908 6010 3932 6012
rect 3988 6010 4012 6012
rect 4068 6010 4092 6012
rect 4148 6010 4154 6012
rect 3908 5958 3910 6010
rect 4090 5958 4092 6010
rect 3846 5956 3852 5958
rect 3908 5956 3932 5958
rect 3988 5956 4012 5958
rect 4068 5956 4092 5958
rect 4148 5956 4154 5958
rect 3846 5936 4154 5956
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 4252 5636 4304 5642
rect 1596 5574 1624 5607
rect 4252 5578 4304 5584
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 2880 5468 3188 5488
rect 2880 5466 2886 5468
rect 2942 5466 2966 5468
rect 3022 5466 3046 5468
rect 3102 5466 3126 5468
rect 3182 5466 3188 5468
rect 2942 5414 2944 5466
rect 3124 5414 3126 5466
rect 2880 5412 2886 5414
rect 2942 5412 2966 5414
rect 3022 5412 3046 5414
rect 3102 5412 3126 5414
rect 3182 5412 3188 5414
rect 2880 5392 3188 5412
rect 3606 5264 3662 5273
rect 3606 5199 3608 5208
rect 3660 5199 3662 5208
rect 3608 5170 3660 5176
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4865 1624 4966
rect 1915 4924 2223 4944
rect 1915 4922 1921 4924
rect 1977 4922 2001 4924
rect 2057 4922 2081 4924
rect 2137 4922 2161 4924
rect 2217 4922 2223 4924
rect 1977 4870 1979 4922
rect 2159 4870 2161 4922
rect 1915 4868 1921 4870
rect 1977 4868 2001 4870
rect 2057 4868 2081 4870
rect 2137 4868 2161 4870
rect 2217 4868 2223 4870
rect 1582 4856 1638 4865
rect 1915 4848 2223 4868
rect 3846 4924 4154 4944
rect 3846 4922 3852 4924
rect 3908 4922 3932 4924
rect 3988 4922 4012 4924
rect 4068 4922 4092 4924
rect 4148 4922 4154 4924
rect 3908 4870 3910 4922
rect 4090 4870 4092 4922
rect 3846 4868 3852 4870
rect 3908 4868 3932 4870
rect 3988 4868 4012 4870
rect 4068 4868 4092 4870
rect 4148 4868 4154 4870
rect 3846 4848 4154 4868
rect 1582 4791 1638 4800
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 1398 4040 1454 4049
rect 1398 3975 1400 3984
rect 1452 3975 1454 3984
rect 1400 3946 1452 3952
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1400 3392 1452 3398
rect 1596 3369 1624 3878
rect 1915 3836 2223 3856
rect 1915 3834 1921 3836
rect 1977 3834 2001 3836
rect 2057 3834 2081 3836
rect 2137 3834 2161 3836
rect 2217 3834 2223 3836
rect 1977 3782 1979 3834
rect 2159 3782 2161 3834
rect 1915 3780 1921 3782
rect 1977 3780 2001 3782
rect 2057 3780 2081 3782
rect 2137 3780 2161 3782
rect 2217 3780 2223 3782
rect 1915 3760 2223 3780
rect 1400 3334 1452 3340
rect 1582 3360 1638 3369
rect 1412 2553 1440 3334
rect 1582 3295 1638 3304
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1398 2544 1454 2553
rect 1398 2479 1454 2488
rect 1504 1873 1532 2790
rect 1915 2748 2223 2768
rect 1915 2746 1921 2748
rect 1977 2746 2001 2748
rect 2057 2746 2081 2748
rect 2137 2746 2161 2748
rect 2217 2746 2223 2748
rect 1977 2694 1979 2746
rect 2159 2694 2161 2746
rect 1915 2692 1921 2694
rect 1977 2692 2001 2694
rect 2057 2692 2081 2694
rect 2137 2692 2161 2694
rect 2217 2692 2223 2694
rect 1915 2672 2223 2692
rect 2332 2446 2360 4422
rect 2608 3058 2636 4422
rect 2792 3534 2820 4422
rect 2880 4380 3188 4400
rect 2880 4378 2886 4380
rect 2942 4378 2966 4380
rect 3022 4378 3046 4380
rect 3102 4378 3126 4380
rect 3182 4378 3188 4380
rect 2942 4326 2944 4378
rect 3124 4326 3126 4378
rect 2880 4324 2886 4326
rect 2942 4324 2966 4326
rect 3022 4324 3046 4326
rect 3102 4324 3126 4326
rect 3182 4324 3188 4326
rect 2880 4304 3188 4324
rect 3846 3836 4154 3856
rect 3846 3834 3852 3836
rect 3908 3834 3932 3836
rect 3988 3834 4012 3836
rect 4068 3834 4092 3836
rect 4148 3834 4154 3836
rect 3908 3782 3910 3834
rect 4090 3782 4092 3834
rect 3846 3780 3852 3782
rect 3908 3780 3932 3782
rect 3988 3780 4012 3782
rect 4068 3780 4092 3782
rect 4148 3780 4154 3782
rect 3846 3760 4154 3780
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2880 3292 3188 3312
rect 2880 3290 2886 3292
rect 2942 3290 2966 3292
rect 3022 3290 3046 3292
rect 3102 3290 3126 3292
rect 3182 3290 3188 3292
rect 2942 3238 2944 3290
rect 3124 3238 3126 3290
rect 2880 3236 2886 3238
rect 2942 3236 2966 3238
rect 3022 3236 3046 3238
rect 3102 3236 3126 3238
rect 3182 3236 3188 3238
rect 2880 3216 3188 3236
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 3846 2748 4154 2768
rect 3846 2746 3852 2748
rect 3908 2746 3932 2748
rect 3988 2746 4012 2748
rect 4068 2746 4092 2748
rect 4148 2746 4154 2748
rect 3908 2694 3910 2746
rect 4090 2694 4092 2746
rect 3846 2692 3852 2694
rect 3908 2692 3932 2694
rect 3988 2692 4012 2694
rect 4068 2692 4092 2694
rect 4148 2692 4154 2694
rect 3846 2672 4154 2692
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 1490 1864 1546 1873
rect 1490 1799 1546 1808
rect 1596 1057 1624 2246
rect 1582 1048 1638 1057
rect 1582 983 1638 992
rect 2792 377 2820 2246
rect 2880 2204 3188 2224
rect 2880 2202 2886 2204
rect 2942 2202 2966 2204
rect 3022 2202 3046 2204
rect 3102 2202 3126 2204
rect 3182 2202 3188 2204
rect 2942 2150 2944 2202
rect 3124 2150 3126 2202
rect 2880 2148 2886 2150
rect 2942 2148 2966 2150
rect 3022 2148 3046 2150
rect 3102 2148 3126 2150
rect 3182 2148 3188 2150
rect 2880 2128 3188 2148
rect 4264 377 4292 5578
rect 4448 5234 4476 6054
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4356 3738 4384 4558
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4448 3194 4476 4626
rect 4540 4146 4568 6122
rect 4632 4554 4660 6258
rect 4724 5574 4752 6666
rect 4811 6556 5119 6576
rect 4811 6554 4817 6556
rect 4873 6554 4897 6556
rect 4953 6554 4977 6556
rect 5033 6554 5057 6556
rect 5113 6554 5119 6556
rect 4873 6502 4875 6554
rect 5055 6502 5057 6554
rect 4811 6500 4817 6502
rect 4873 6500 4897 6502
rect 4953 6500 4977 6502
rect 5033 6500 5057 6502
rect 5113 6500 5119 6502
rect 4811 6480 5119 6500
rect 5276 6497 5304 6886
rect 5262 6488 5318 6497
rect 5262 6423 5318 6432
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4526 3632 4582 3641
rect 4526 3567 4582 3576
rect 4540 3534 4568 3567
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4632 3126 4660 4490
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4724 3058 4752 5510
rect 4811 5468 5119 5488
rect 4811 5466 4817 5468
rect 4873 5466 4897 5468
rect 4953 5466 4977 5468
rect 5033 5466 5057 5468
rect 5113 5466 5119 5468
rect 4873 5414 4875 5466
rect 5055 5414 5057 5466
rect 4811 5412 4817 5414
rect 4873 5412 4897 5414
rect 4953 5412 4977 5414
rect 5033 5412 5057 5414
rect 5113 5412 5119 5414
rect 4811 5392 5119 5412
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4816 4826 4844 5238
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5368 4690 5396 7142
rect 5776 7100 6084 7120
rect 5776 7098 5782 7100
rect 5838 7098 5862 7100
rect 5918 7098 5942 7100
rect 5998 7098 6022 7100
rect 6078 7098 6084 7100
rect 5838 7046 5840 7098
rect 6020 7046 6022 7098
rect 5776 7044 5782 7046
rect 5838 7044 5862 7046
rect 5918 7044 5942 7046
rect 5998 7044 6022 7046
rect 6078 7044 6084 7046
rect 5776 7024 6084 7044
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5460 5137 5488 6258
rect 5644 5370 5672 6870
rect 6196 6730 6224 8774
rect 6918 8735 6974 8744
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 5776 6012 6084 6032
rect 5776 6010 5782 6012
rect 5838 6010 5862 6012
rect 5918 6010 5942 6012
rect 5998 6010 6022 6012
rect 6078 6010 6084 6012
rect 5838 5958 5840 6010
rect 6020 5958 6022 6010
rect 5776 5956 5782 5958
rect 5838 5956 5862 5958
rect 5918 5956 5942 5958
rect 5998 5956 6022 5958
rect 6078 5956 6084 5958
rect 5776 5936 6084 5956
rect 6288 5710 6316 7686
rect 7012 7064 7064 7070
rect 7010 7032 7012 7041
rect 7064 7032 7066 7041
rect 7010 6967 7066 6976
rect 7012 5976 7064 5982
rect 7010 5944 7012 5953
rect 7064 5944 7066 5953
rect 7010 5879 7066 5888
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5446 5128 5502 5137
rect 5446 5063 5502 5072
rect 5776 4924 6084 4944
rect 5776 4922 5782 4924
rect 5838 4922 5862 4924
rect 5918 4922 5942 4924
rect 5998 4922 6022 4924
rect 6078 4922 6084 4924
rect 5838 4870 5840 4922
rect 6020 4870 6022 4922
rect 5776 4868 5782 4870
rect 5838 4868 5862 4870
rect 5918 4868 5942 4870
rect 5998 4868 6022 4870
rect 6078 4868 6084 4870
rect 5776 4848 6084 4868
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4811 4380 5119 4400
rect 4811 4378 4817 4380
rect 4873 4378 4897 4380
rect 4953 4378 4977 4380
rect 5033 4378 5057 4380
rect 5113 4378 5119 4380
rect 4873 4326 4875 4378
rect 5055 4326 5057 4378
rect 4811 4324 4817 4326
rect 4873 4324 4897 4326
rect 4953 4324 4977 4326
rect 5033 4324 5057 4326
rect 5113 4324 5119 4326
rect 4811 4304 5119 4324
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 3738 5028 4082
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5184 3346 5212 4626
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5262 4312 5318 4321
rect 5262 4247 5318 4256
rect 5276 3534 5304 4247
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5184 3318 5304 3346
rect 4811 3292 5119 3312
rect 4811 3290 4817 3292
rect 4873 3290 4897 3292
rect 4953 3290 4977 3292
rect 5033 3290 5057 3292
rect 5113 3290 5119 3292
rect 4873 3238 4875 3290
rect 5055 3238 5057 3290
rect 4811 3236 4817 3238
rect 4873 3236 4897 3238
rect 4953 3236 4977 3238
rect 5033 3236 5057 3238
rect 5113 3236 5119 3238
rect 4811 3216 5119 3236
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5184 2553 5212 2994
rect 5170 2544 5226 2553
rect 5276 2514 5304 3318
rect 5368 2582 5396 4490
rect 5460 2650 5488 4558
rect 5552 3194 5580 4558
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 3534 5672 3878
rect 5776 3836 6084 3856
rect 5776 3834 5782 3836
rect 5838 3834 5862 3836
rect 5918 3834 5942 3836
rect 5998 3834 6022 3836
rect 6078 3834 6084 3836
rect 5838 3782 5840 3834
rect 6020 3782 6022 3834
rect 5776 3780 5782 3782
rect 5838 3780 5862 3782
rect 5918 3780 5942 3782
rect 5998 3780 6022 3782
rect 6078 3780 6084 3782
rect 5776 3760 6084 3780
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6012 3097 6040 3334
rect 5998 3088 6054 3097
rect 5998 3023 6054 3032
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 5776 2748 6084 2768
rect 5776 2746 5782 2748
rect 5838 2746 5862 2748
rect 5918 2746 5942 2748
rect 5998 2746 6022 2748
rect 6078 2746 6084 2748
rect 5838 2694 5840 2746
rect 6020 2694 6022 2746
rect 5776 2692 5782 2694
rect 5838 2692 5862 2694
rect 5918 2692 5942 2694
rect 5998 2692 6022 2694
rect 6078 2692 6084 2694
rect 5776 2672 6084 2692
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 5170 2479 5226 2488
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 4811 2204 5119 2224
rect 4811 2202 4817 2204
rect 4873 2202 4897 2204
rect 4953 2202 4977 2204
rect 5033 2202 5057 2204
rect 5113 2202 5119 2204
rect 4873 2150 4875 2202
rect 5055 2150 5057 2202
rect 4811 2148 4817 2150
rect 4873 2148 4897 2150
rect 4953 2148 4977 2150
rect 5033 2148 5057 2150
rect 5113 2148 5119 2150
rect 4811 2128 5119 2148
rect 5184 1465 5212 2382
rect 5170 1456 5226 1465
rect 5170 1391 5226 1400
rect 5828 921 5856 2382
rect 6196 2009 6224 2994
rect 6182 2000 6238 2009
rect 6182 1935 6238 1944
rect 5814 912 5870 921
rect 5814 847 5870 856
rect 2778 368 2834 377
rect 2778 303 2834 312
rect 4250 368 4306 377
rect 4250 303 4306 312
<< via2 >>
rect 4526 59608 4582 59664
rect 3330 59472 3386 59528
rect 3238 58656 3294 58712
rect 2778 57976 2834 58032
rect 2886 57690 2942 57692
rect 2966 57690 3022 57692
rect 3046 57690 3102 57692
rect 3126 57690 3182 57692
rect 2886 57638 2932 57690
rect 2932 57638 2942 57690
rect 2966 57638 2996 57690
rect 2996 57638 3008 57690
rect 3008 57638 3022 57690
rect 3046 57638 3060 57690
rect 3060 57638 3072 57690
rect 3072 57638 3102 57690
rect 3126 57638 3136 57690
rect 3136 57638 3182 57690
rect 2886 57636 2942 57638
rect 2966 57636 3022 57638
rect 3046 57636 3102 57638
rect 3126 57636 3182 57638
rect 1582 57196 1584 57216
rect 1584 57196 1636 57216
rect 1636 57196 1638 57216
rect 1582 57160 1638 57196
rect 1921 57146 1977 57148
rect 2001 57146 2057 57148
rect 2081 57146 2137 57148
rect 2161 57146 2217 57148
rect 1921 57094 1967 57146
rect 1967 57094 1977 57146
rect 2001 57094 2031 57146
rect 2031 57094 2043 57146
rect 2043 57094 2057 57146
rect 2081 57094 2095 57146
rect 2095 57094 2107 57146
rect 2107 57094 2137 57146
rect 2161 57094 2171 57146
rect 2171 57094 2217 57146
rect 1921 57092 1977 57094
rect 2001 57092 2057 57094
rect 2081 57092 2137 57094
rect 2161 57092 2217 57094
rect 1582 56480 1638 56536
rect 1921 56058 1977 56060
rect 2001 56058 2057 56060
rect 2081 56058 2137 56060
rect 2161 56058 2217 56060
rect 1921 56006 1967 56058
rect 1967 56006 1977 56058
rect 2001 56006 2031 56058
rect 2031 56006 2043 56058
rect 2043 56006 2057 56058
rect 2081 56006 2095 56058
rect 2095 56006 2107 56058
rect 2107 56006 2137 56058
rect 2161 56006 2171 56058
rect 2171 56006 2217 56058
rect 1921 56004 1977 56006
rect 2001 56004 2057 56006
rect 2081 56004 2137 56006
rect 2161 56004 2217 56006
rect 1582 55664 1638 55720
rect 2886 56602 2942 56604
rect 2966 56602 3022 56604
rect 3046 56602 3102 56604
rect 3126 56602 3182 56604
rect 2886 56550 2932 56602
rect 2932 56550 2942 56602
rect 2966 56550 2996 56602
rect 2996 56550 3008 56602
rect 3008 56550 3022 56602
rect 3046 56550 3060 56602
rect 3060 56550 3072 56602
rect 3072 56550 3102 56602
rect 3126 56550 3136 56602
rect 3136 56550 3182 56602
rect 2886 56548 2942 56550
rect 2966 56548 3022 56550
rect 3046 56548 3102 56550
rect 3126 56548 3182 56550
rect 2886 55514 2942 55516
rect 2966 55514 3022 55516
rect 3046 55514 3102 55516
rect 3126 55514 3182 55516
rect 2886 55462 2932 55514
rect 2932 55462 2942 55514
rect 2966 55462 2996 55514
rect 2996 55462 3008 55514
rect 3008 55462 3022 55514
rect 3046 55462 3060 55514
rect 3060 55462 3072 55514
rect 3072 55462 3102 55514
rect 3126 55462 3136 55514
rect 3136 55462 3182 55514
rect 2886 55460 2942 55462
rect 2966 55460 3022 55462
rect 3046 55460 3102 55462
rect 3126 55460 3182 55462
rect 4250 59064 4306 59120
rect 1921 54970 1977 54972
rect 2001 54970 2057 54972
rect 2081 54970 2137 54972
rect 2161 54970 2217 54972
rect 1921 54918 1967 54970
rect 1967 54918 1977 54970
rect 2001 54918 2031 54970
rect 2031 54918 2043 54970
rect 2043 54918 2057 54970
rect 2081 54918 2095 54970
rect 2095 54918 2107 54970
rect 2107 54918 2137 54970
rect 2161 54918 2171 54970
rect 2171 54918 2217 54970
rect 1921 54916 1977 54918
rect 2001 54916 2057 54918
rect 2081 54916 2137 54918
rect 2161 54916 2217 54918
rect 1582 54848 1638 54904
rect 1582 54168 1638 54224
rect 1582 53388 1584 53408
rect 1584 53388 1636 53408
rect 1636 53388 1638 53408
rect 1582 53352 1638 53388
rect 1582 52672 1638 52728
rect 1582 51876 1638 51912
rect 1582 51856 1584 51876
rect 1584 51856 1636 51876
rect 1636 51856 1638 51876
rect 1582 51212 1584 51232
rect 1584 51212 1636 51232
rect 1636 51212 1638 51232
rect 1582 51176 1638 51212
rect 1582 50360 1638 50416
rect 1582 49580 1584 49600
rect 1584 49580 1636 49600
rect 1636 49580 1638 49600
rect 1582 49544 1638 49580
rect 1582 48864 1638 48920
rect 1582 48048 1638 48104
rect 1582 47404 1584 47424
rect 1584 47404 1636 47424
rect 1636 47404 1638 47424
rect 1582 47368 1638 47404
rect 1582 46552 1638 46608
rect 1582 45772 1584 45792
rect 1584 45772 1636 45792
rect 1636 45772 1638 45792
rect 1582 45736 1638 45772
rect 1582 45056 1638 45112
rect 1582 44260 1638 44296
rect 1582 44240 1584 44260
rect 1584 44240 1636 44260
rect 1636 44240 1638 44260
rect 1582 43596 1584 43616
rect 1584 43596 1636 43616
rect 1636 43596 1638 43616
rect 1582 43560 1638 43596
rect 1582 42744 1638 42800
rect 1582 42084 1638 42120
rect 1582 42064 1584 42084
rect 1584 42064 1636 42084
rect 1636 42064 1638 42084
rect 1490 41792 1546 41848
rect 1490 41384 1546 41440
rect 1306 35980 1308 36000
rect 1308 35980 1360 36000
rect 1360 35980 1362 36000
rect 1306 35944 1362 35980
rect 1582 41248 1638 41304
rect 1582 40432 1638 40488
rect 1582 39752 1638 39808
rect 1582 38936 1638 38992
rect 1582 38256 1638 38312
rect 1582 37440 1638 37496
rect 1921 53882 1977 53884
rect 2001 53882 2057 53884
rect 2081 53882 2137 53884
rect 2161 53882 2217 53884
rect 1921 53830 1967 53882
rect 1967 53830 1977 53882
rect 2001 53830 2031 53882
rect 2031 53830 2043 53882
rect 2043 53830 2057 53882
rect 2081 53830 2095 53882
rect 2095 53830 2107 53882
rect 2107 53830 2137 53882
rect 2161 53830 2171 53882
rect 2171 53830 2217 53882
rect 1921 53828 1977 53830
rect 2001 53828 2057 53830
rect 2081 53828 2137 53830
rect 2161 53828 2217 53830
rect 1921 52794 1977 52796
rect 2001 52794 2057 52796
rect 2081 52794 2137 52796
rect 2161 52794 2217 52796
rect 1921 52742 1967 52794
rect 1967 52742 1977 52794
rect 2001 52742 2031 52794
rect 2031 52742 2043 52794
rect 2043 52742 2057 52794
rect 2081 52742 2095 52794
rect 2095 52742 2107 52794
rect 2107 52742 2137 52794
rect 2161 52742 2171 52794
rect 2171 52742 2217 52794
rect 1921 52740 1977 52742
rect 2001 52740 2057 52742
rect 2081 52740 2137 52742
rect 2161 52740 2217 52742
rect 1921 51706 1977 51708
rect 2001 51706 2057 51708
rect 2081 51706 2137 51708
rect 2161 51706 2217 51708
rect 1921 51654 1967 51706
rect 1967 51654 1977 51706
rect 2001 51654 2031 51706
rect 2031 51654 2043 51706
rect 2043 51654 2057 51706
rect 2081 51654 2095 51706
rect 2095 51654 2107 51706
rect 2107 51654 2137 51706
rect 2161 51654 2171 51706
rect 2171 51654 2217 51706
rect 1921 51652 1977 51654
rect 2001 51652 2057 51654
rect 2081 51652 2137 51654
rect 2161 51652 2217 51654
rect 2886 54426 2942 54428
rect 2966 54426 3022 54428
rect 3046 54426 3102 54428
rect 3126 54426 3182 54428
rect 2886 54374 2932 54426
rect 2932 54374 2942 54426
rect 2966 54374 2996 54426
rect 2996 54374 3008 54426
rect 3008 54374 3022 54426
rect 3046 54374 3060 54426
rect 3060 54374 3072 54426
rect 3072 54374 3102 54426
rect 3126 54374 3136 54426
rect 3136 54374 3182 54426
rect 2886 54372 2942 54374
rect 2966 54372 3022 54374
rect 3046 54372 3102 54374
rect 3126 54372 3182 54374
rect 3852 57146 3908 57148
rect 3932 57146 3988 57148
rect 4012 57146 4068 57148
rect 4092 57146 4148 57148
rect 3852 57094 3898 57146
rect 3898 57094 3908 57146
rect 3932 57094 3962 57146
rect 3962 57094 3974 57146
rect 3974 57094 3988 57146
rect 4012 57094 4026 57146
rect 4026 57094 4038 57146
rect 4038 57094 4068 57146
rect 4092 57094 4102 57146
rect 4102 57094 4148 57146
rect 3852 57092 3908 57094
rect 3932 57092 3988 57094
rect 4012 57092 4068 57094
rect 4092 57092 4148 57094
rect 3852 56058 3908 56060
rect 3932 56058 3988 56060
rect 4012 56058 4068 56060
rect 4092 56058 4148 56060
rect 3852 56006 3898 56058
rect 3898 56006 3908 56058
rect 3932 56006 3962 56058
rect 3962 56006 3974 56058
rect 3974 56006 3988 56058
rect 4012 56006 4026 56058
rect 4026 56006 4038 56058
rect 4038 56006 4068 56058
rect 4092 56006 4102 56058
rect 4102 56006 4148 56058
rect 3852 56004 3908 56006
rect 3932 56004 3988 56006
rect 4012 56004 4068 56006
rect 4092 56004 4148 56006
rect 5262 58520 5318 58576
rect 4817 57690 4873 57692
rect 4897 57690 4953 57692
rect 4977 57690 5033 57692
rect 5057 57690 5113 57692
rect 4817 57638 4863 57690
rect 4863 57638 4873 57690
rect 4897 57638 4927 57690
rect 4927 57638 4939 57690
rect 4939 57638 4953 57690
rect 4977 57638 4991 57690
rect 4991 57638 5003 57690
rect 5003 57638 5033 57690
rect 5057 57638 5067 57690
rect 5067 57638 5113 57690
rect 4817 57636 4873 57638
rect 4897 57636 4953 57638
rect 4977 57636 5033 57638
rect 5057 57636 5113 57638
rect 4250 55276 4306 55312
rect 4250 55256 4252 55276
rect 4252 55256 4304 55276
rect 4304 55256 4306 55276
rect 3852 54970 3908 54972
rect 3932 54970 3988 54972
rect 4012 54970 4068 54972
rect 4092 54970 4148 54972
rect 3852 54918 3898 54970
rect 3898 54918 3908 54970
rect 3932 54918 3962 54970
rect 3962 54918 3974 54970
rect 3974 54918 3988 54970
rect 4012 54918 4026 54970
rect 4026 54918 4038 54970
rect 4038 54918 4068 54970
rect 4092 54918 4102 54970
rect 4102 54918 4148 54970
rect 3852 54916 3908 54918
rect 3932 54916 3988 54918
rect 4012 54916 4068 54918
rect 4092 54916 4148 54918
rect 2886 53338 2942 53340
rect 2966 53338 3022 53340
rect 3046 53338 3102 53340
rect 3126 53338 3182 53340
rect 2886 53286 2932 53338
rect 2932 53286 2942 53338
rect 2966 53286 2996 53338
rect 2996 53286 3008 53338
rect 3008 53286 3022 53338
rect 3046 53286 3060 53338
rect 3060 53286 3072 53338
rect 3072 53286 3102 53338
rect 3126 53286 3136 53338
rect 3136 53286 3182 53338
rect 2886 53284 2942 53286
rect 2966 53284 3022 53286
rect 3046 53284 3102 53286
rect 3126 53284 3182 53286
rect 1921 50618 1977 50620
rect 2001 50618 2057 50620
rect 2081 50618 2137 50620
rect 2161 50618 2217 50620
rect 1921 50566 1967 50618
rect 1967 50566 1977 50618
rect 2001 50566 2031 50618
rect 2031 50566 2043 50618
rect 2043 50566 2057 50618
rect 2081 50566 2095 50618
rect 2095 50566 2107 50618
rect 2107 50566 2137 50618
rect 2161 50566 2171 50618
rect 2171 50566 2217 50618
rect 1921 50564 1977 50566
rect 2001 50564 2057 50566
rect 2081 50564 2137 50566
rect 2161 50564 2217 50566
rect 1921 49530 1977 49532
rect 2001 49530 2057 49532
rect 2081 49530 2137 49532
rect 2161 49530 2217 49532
rect 1921 49478 1967 49530
rect 1967 49478 1977 49530
rect 2001 49478 2031 49530
rect 2031 49478 2043 49530
rect 2043 49478 2057 49530
rect 2081 49478 2095 49530
rect 2095 49478 2107 49530
rect 2107 49478 2137 49530
rect 2161 49478 2171 49530
rect 2171 49478 2217 49530
rect 1921 49476 1977 49478
rect 2001 49476 2057 49478
rect 2081 49476 2137 49478
rect 2161 49476 2217 49478
rect 1921 48442 1977 48444
rect 2001 48442 2057 48444
rect 2081 48442 2137 48444
rect 2161 48442 2217 48444
rect 1921 48390 1967 48442
rect 1967 48390 1977 48442
rect 2001 48390 2031 48442
rect 2031 48390 2043 48442
rect 2043 48390 2057 48442
rect 2081 48390 2095 48442
rect 2095 48390 2107 48442
rect 2107 48390 2137 48442
rect 2161 48390 2171 48442
rect 2171 48390 2217 48442
rect 1921 48388 1977 48390
rect 2001 48388 2057 48390
rect 2081 48388 2137 48390
rect 2161 48388 2217 48390
rect 1921 47354 1977 47356
rect 2001 47354 2057 47356
rect 2081 47354 2137 47356
rect 2161 47354 2217 47356
rect 1921 47302 1967 47354
rect 1967 47302 1977 47354
rect 2001 47302 2031 47354
rect 2031 47302 2043 47354
rect 2043 47302 2057 47354
rect 2081 47302 2095 47354
rect 2095 47302 2107 47354
rect 2107 47302 2137 47354
rect 2161 47302 2171 47354
rect 2171 47302 2217 47354
rect 1921 47300 1977 47302
rect 2001 47300 2057 47302
rect 2081 47300 2137 47302
rect 2161 47300 2217 47302
rect 1921 46266 1977 46268
rect 2001 46266 2057 46268
rect 2081 46266 2137 46268
rect 2161 46266 2217 46268
rect 1921 46214 1967 46266
rect 1967 46214 1977 46266
rect 2001 46214 2031 46266
rect 2031 46214 2043 46266
rect 2043 46214 2057 46266
rect 2081 46214 2095 46266
rect 2095 46214 2107 46266
rect 2107 46214 2137 46266
rect 2161 46214 2171 46266
rect 2171 46214 2217 46266
rect 1921 46212 1977 46214
rect 2001 46212 2057 46214
rect 2081 46212 2137 46214
rect 2161 46212 2217 46214
rect 1921 45178 1977 45180
rect 2001 45178 2057 45180
rect 2081 45178 2137 45180
rect 2161 45178 2217 45180
rect 1921 45126 1967 45178
rect 1967 45126 1977 45178
rect 2001 45126 2031 45178
rect 2031 45126 2043 45178
rect 2043 45126 2057 45178
rect 2081 45126 2095 45178
rect 2095 45126 2107 45178
rect 2107 45126 2137 45178
rect 2161 45126 2171 45178
rect 2171 45126 2217 45178
rect 1921 45124 1977 45126
rect 2001 45124 2057 45126
rect 2081 45124 2137 45126
rect 2161 45124 2217 45126
rect 1921 44090 1977 44092
rect 2001 44090 2057 44092
rect 2081 44090 2137 44092
rect 2161 44090 2217 44092
rect 1921 44038 1967 44090
rect 1967 44038 1977 44090
rect 2001 44038 2031 44090
rect 2031 44038 2043 44090
rect 2043 44038 2057 44090
rect 2081 44038 2095 44090
rect 2095 44038 2107 44090
rect 2107 44038 2137 44090
rect 2161 44038 2171 44090
rect 2171 44038 2217 44090
rect 1921 44036 1977 44038
rect 2001 44036 2057 44038
rect 2081 44036 2137 44038
rect 2161 44036 2217 44038
rect 1921 43002 1977 43004
rect 2001 43002 2057 43004
rect 2081 43002 2137 43004
rect 2161 43002 2217 43004
rect 1921 42950 1967 43002
rect 1967 42950 1977 43002
rect 2001 42950 2031 43002
rect 2031 42950 2043 43002
rect 2043 42950 2057 43002
rect 2081 42950 2095 43002
rect 2095 42950 2107 43002
rect 2107 42950 2137 43002
rect 2161 42950 2171 43002
rect 2171 42950 2217 43002
rect 1921 42948 1977 42950
rect 2001 42948 2057 42950
rect 2081 42948 2137 42950
rect 2161 42948 2217 42950
rect 1921 41914 1977 41916
rect 2001 41914 2057 41916
rect 2081 41914 2137 41916
rect 2161 41914 2217 41916
rect 1921 41862 1967 41914
rect 1967 41862 1977 41914
rect 2001 41862 2031 41914
rect 2031 41862 2043 41914
rect 2043 41862 2057 41914
rect 2081 41862 2095 41914
rect 2095 41862 2107 41914
rect 2107 41862 2137 41914
rect 2161 41862 2171 41914
rect 2171 41862 2217 41914
rect 1921 41860 1977 41862
rect 2001 41860 2057 41862
rect 2081 41860 2137 41862
rect 2161 41860 2217 41862
rect 1921 40826 1977 40828
rect 2001 40826 2057 40828
rect 2081 40826 2137 40828
rect 2161 40826 2217 40828
rect 1921 40774 1967 40826
rect 1967 40774 1977 40826
rect 2001 40774 2031 40826
rect 2031 40774 2043 40826
rect 2043 40774 2057 40826
rect 2081 40774 2095 40826
rect 2095 40774 2107 40826
rect 2107 40774 2137 40826
rect 2161 40774 2171 40826
rect 2171 40774 2217 40826
rect 1921 40772 1977 40774
rect 2001 40772 2057 40774
rect 2081 40772 2137 40774
rect 2161 40772 2217 40774
rect 1921 39738 1977 39740
rect 2001 39738 2057 39740
rect 2081 39738 2137 39740
rect 2161 39738 2217 39740
rect 1921 39686 1967 39738
rect 1967 39686 1977 39738
rect 2001 39686 2031 39738
rect 2031 39686 2043 39738
rect 2043 39686 2057 39738
rect 2081 39686 2095 39738
rect 2095 39686 2107 39738
rect 2107 39686 2137 39738
rect 2161 39686 2171 39738
rect 2171 39686 2217 39738
rect 1921 39684 1977 39686
rect 2001 39684 2057 39686
rect 2081 39684 2137 39686
rect 2161 39684 2217 39686
rect 1921 38650 1977 38652
rect 2001 38650 2057 38652
rect 2081 38650 2137 38652
rect 2161 38650 2217 38652
rect 1921 38598 1967 38650
rect 1967 38598 1977 38650
rect 2001 38598 2031 38650
rect 2031 38598 2043 38650
rect 2043 38598 2057 38650
rect 2081 38598 2095 38650
rect 2095 38598 2107 38650
rect 2107 38598 2137 38650
rect 2161 38598 2171 38650
rect 2171 38598 2217 38650
rect 1921 38596 1977 38598
rect 2001 38596 2057 38598
rect 2081 38596 2137 38598
rect 2161 38596 2217 38598
rect 2886 52250 2942 52252
rect 2966 52250 3022 52252
rect 3046 52250 3102 52252
rect 3126 52250 3182 52252
rect 2886 52198 2932 52250
rect 2932 52198 2942 52250
rect 2966 52198 2996 52250
rect 2996 52198 3008 52250
rect 3008 52198 3022 52250
rect 3046 52198 3060 52250
rect 3060 52198 3072 52250
rect 3072 52198 3102 52250
rect 3126 52198 3136 52250
rect 3136 52198 3182 52250
rect 2886 52196 2942 52198
rect 2966 52196 3022 52198
rect 3046 52196 3102 52198
rect 3126 52196 3182 52198
rect 2886 51162 2942 51164
rect 2966 51162 3022 51164
rect 3046 51162 3102 51164
rect 3126 51162 3182 51164
rect 2886 51110 2932 51162
rect 2932 51110 2942 51162
rect 2966 51110 2996 51162
rect 2996 51110 3008 51162
rect 3008 51110 3022 51162
rect 3046 51110 3060 51162
rect 3060 51110 3072 51162
rect 3072 51110 3102 51162
rect 3126 51110 3136 51162
rect 3136 51110 3182 51162
rect 2886 51108 2942 51110
rect 2966 51108 3022 51110
rect 3046 51108 3102 51110
rect 3126 51108 3182 51110
rect 2410 38664 2466 38720
rect 2594 38392 2650 38448
rect 1921 37562 1977 37564
rect 2001 37562 2057 37564
rect 2081 37562 2137 37564
rect 2161 37562 2217 37564
rect 1921 37510 1967 37562
rect 1967 37510 1977 37562
rect 2001 37510 2031 37562
rect 2031 37510 2043 37562
rect 2043 37510 2057 37562
rect 2081 37510 2095 37562
rect 2095 37510 2107 37562
rect 2107 37510 2137 37562
rect 2161 37510 2171 37562
rect 2171 37510 2217 37562
rect 1921 37508 1977 37510
rect 2001 37508 2057 37510
rect 2081 37508 2137 37510
rect 2161 37508 2217 37510
rect 1582 36644 1638 36680
rect 1582 36624 1584 36644
rect 1584 36624 1636 36644
rect 1636 36624 1638 36644
rect 1398 35128 1454 35184
rect 1398 32952 1454 33008
rect 1398 32136 1454 32192
rect 1398 30676 1400 30696
rect 1400 30676 1452 30696
rect 1452 30676 1454 30696
rect 1398 30640 1454 30676
rect 1398 29824 1454 29880
rect 1398 28328 1454 28384
rect 1674 34312 1730 34368
rect 1582 34040 1638 34096
rect 1582 29144 1638 29200
rect 1921 36474 1977 36476
rect 2001 36474 2057 36476
rect 2081 36474 2137 36476
rect 2161 36474 2217 36476
rect 1921 36422 1967 36474
rect 1967 36422 1977 36474
rect 2001 36422 2031 36474
rect 2031 36422 2043 36474
rect 2043 36422 2057 36474
rect 2081 36422 2095 36474
rect 2095 36422 2107 36474
rect 2107 36422 2137 36474
rect 2161 36422 2171 36474
rect 2171 36422 2217 36474
rect 1921 36420 1977 36422
rect 2001 36420 2057 36422
rect 2081 36420 2137 36422
rect 2161 36420 2217 36422
rect 1921 35386 1977 35388
rect 2001 35386 2057 35388
rect 2081 35386 2137 35388
rect 2161 35386 2217 35388
rect 1921 35334 1967 35386
rect 1967 35334 1977 35386
rect 2001 35334 2031 35386
rect 2031 35334 2043 35386
rect 2043 35334 2057 35386
rect 2081 35334 2095 35386
rect 2095 35334 2107 35386
rect 2107 35334 2137 35386
rect 2161 35334 2171 35386
rect 2171 35334 2217 35386
rect 1921 35332 1977 35334
rect 2001 35332 2057 35334
rect 2081 35332 2137 35334
rect 2161 35332 2217 35334
rect 1858 34448 1914 34504
rect 1921 34298 1977 34300
rect 2001 34298 2057 34300
rect 2081 34298 2137 34300
rect 2161 34298 2217 34300
rect 1921 34246 1967 34298
rect 1967 34246 1977 34298
rect 2001 34246 2031 34298
rect 2031 34246 2043 34298
rect 2043 34246 2057 34298
rect 2081 34246 2095 34298
rect 2095 34246 2107 34298
rect 2107 34246 2137 34298
rect 2161 34246 2171 34298
rect 2171 34246 2217 34298
rect 1921 34244 1977 34246
rect 2001 34244 2057 34246
rect 2081 34244 2137 34246
rect 2161 34244 2217 34246
rect 1858 33632 1914 33688
rect 1921 33210 1977 33212
rect 2001 33210 2057 33212
rect 2081 33210 2137 33212
rect 2161 33210 2217 33212
rect 1921 33158 1967 33210
rect 1967 33158 1977 33210
rect 2001 33158 2031 33210
rect 2031 33158 2043 33210
rect 2043 33158 2057 33210
rect 2081 33158 2095 33210
rect 2095 33158 2107 33210
rect 2107 33158 2137 33210
rect 2161 33158 2171 33210
rect 2171 33158 2217 33210
rect 1921 33156 1977 33158
rect 2001 33156 2057 33158
rect 2081 33156 2137 33158
rect 2161 33156 2217 33158
rect 2042 32816 2098 32872
rect 1921 32122 1977 32124
rect 2001 32122 2057 32124
rect 2081 32122 2137 32124
rect 2161 32122 2217 32124
rect 1921 32070 1967 32122
rect 1967 32070 1977 32122
rect 2001 32070 2031 32122
rect 2031 32070 2043 32122
rect 2043 32070 2057 32122
rect 2081 32070 2095 32122
rect 2095 32070 2107 32122
rect 2107 32070 2137 32122
rect 2161 32070 2171 32122
rect 2171 32070 2217 32122
rect 1921 32068 1977 32070
rect 2001 32068 2057 32070
rect 2081 32068 2137 32070
rect 2161 32068 2217 32070
rect 2686 36896 2742 36952
rect 2886 50074 2942 50076
rect 2966 50074 3022 50076
rect 3046 50074 3102 50076
rect 3126 50074 3182 50076
rect 2886 50022 2932 50074
rect 2932 50022 2942 50074
rect 2966 50022 2996 50074
rect 2996 50022 3008 50074
rect 3008 50022 3022 50074
rect 3046 50022 3060 50074
rect 3060 50022 3072 50074
rect 3072 50022 3102 50074
rect 3126 50022 3136 50074
rect 3136 50022 3182 50074
rect 2886 50020 2942 50022
rect 2966 50020 3022 50022
rect 3046 50020 3102 50022
rect 3126 50020 3182 50022
rect 2886 48986 2942 48988
rect 2966 48986 3022 48988
rect 3046 48986 3102 48988
rect 3126 48986 3182 48988
rect 2886 48934 2932 48986
rect 2932 48934 2942 48986
rect 2966 48934 2996 48986
rect 2996 48934 3008 48986
rect 3008 48934 3022 48986
rect 3046 48934 3060 48986
rect 3060 48934 3072 48986
rect 3072 48934 3102 48986
rect 3126 48934 3136 48986
rect 3136 48934 3182 48986
rect 2886 48932 2942 48934
rect 2966 48932 3022 48934
rect 3046 48932 3102 48934
rect 3126 48932 3182 48934
rect 2870 48084 2872 48104
rect 2872 48084 2924 48104
rect 2924 48084 2926 48104
rect 2870 48048 2926 48084
rect 2886 47898 2942 47900
rect 2966 47898 3022 47900
rect 3046 47898 3102 47900
rect 3126 47898 3182 47900
rect 2886 47846 2932 47898
rect 2932 47846 2942 47898
rect 2966 47846 2996 47898
rect 2996 47846 3008 47898
rect 3008 47846 3022 47898
rect 3046 47846 3060 47898
rect 3060 47846 3072 47898
rect 3072 47846 3102 47898
rect 3126 47846 3136 47898
rect 3136 47846 3182 47898
rect 2886 47844 2942 47846
rect 2966 47844 3022 47846
rect 3046 47844 3102 47846
rect 3126 47844 3182 47846
rect 2886 46810 2942 46812
rect 2966 46810 3022 46812
rect 3046 46810 3102 46812
rect 3126 46810 3182 46812
rect 2886 46758 2932 46810
rect 2932 46758 2942 46810
rect 2966 46758 2996 46810
rect 2996 46758 3008 46810
rect 3008 46758 3022 46810
rect 3046 46758 3060 46810
rect 3060 46758 3072 46810
rect 3072 46758 3102 46810
rect 3126 46758 3136 46810
rect 3136 46758 3182 46810
rect 2886 46756 2942 46758
rect 2966 46756 3022 46758
rect 3046 46756 3102 46758
rect 3126 46756 3182 46758
rect 3852 53882 3908 53884
rect 3932 53882 3988 53884
rect 4012 53882 4068 53884
rect 4092 53882 4148 53884
rect 3852 53830 3898 53882
rect 3898 53830 3908 53882
rect 3932 53830 3962 53882
rect 3962 53830 3974 53882
rect 3974 53830 3988 53882
rect 4012 53830 4026 53882
rect 4026 53830 4038 53882
rect 4038 53830 4068 53882
rect 4092 53830 4102 53882
rect 4102 53830 4148 53882
rect 3852 53828 3908 53830
rect 3932 53828 3988 53830
rect 4012 53828 4068 53830
rect 4092 53828 4148 53830
rect 3852 52794 3908 52796
rect 3932 52794 3988 52796
rect 4012 52794 4068 52796
rect 4092 52794 4148 52796
rect 3852 52742 3898 52794
rect 3898 52742 3908 52794
rect 3932 52742 3962 52794
rect 3962 52742 3974 52794
rect 3974 52742 3988 52794
rect 4012 52742 4026 52794
rect 4026 52742 4038 52794
rect 4038 52742 4068 52794
rect 4092 52742 4102 52794
rect 4102 52742 4148 52794
rect 3852 52740 3908 52742
rect 3932 52740 3988 52742
rect 4012 52740 4068 52742
rect 4092 52740 4148 52742
rect 2886 45722 2942 45724
rect 2966 45722 3022 45724
rect 3046 45722 3102 45724
rect 3126 45722 3182 45724
rect 2886 45670 2932 45722
rect 2932 45670 2942 45722
rect 2966 45670 2996 45722
rect 2996 45670 3008 45722
rect 3008 45670 3022 45722
rect 3046 45670 3060 45722
rect 3060 45670 3072 45722
rect 3072 45670 3102 45722
rect 3126 45670 3136 45722
rect 3136 45670 3182 45722
rect 2886 45668 2942 45670
rect 2966 45668 3022 45670
rect 3046 45668 3102 45670
rect 3126 45668 3182 45670
rect 2886 44634 2942 44636
rect 2966 44634 3022 44636
rect 3046 44634 3102 44636
rect 3126 44634 3182 44636
rect 2886 44582 2932 44634
rect 2932 44582 2942 44634
rect 2966 44582 2996 44634
rect 2996 44582 3008 44634
rect 3008 44582 3022 44634
rect 3046 44582 3060 44634
rect 3060 44582 3072 44634
rect 3072 44582 3102 44634
rect 3126 44582 3136 44634
rect 3136 44582 3182 44634
rect 2886 44580 2942 44582
rect 2966 44580 3022 44582
rect 3046 44580 3102 44582
rect 3126 44580 3182 44582
rect 3146 43696 3202 43752
rect 2886 43546 2942 43548
rect 2966 43546 3022 43548
rect 3046 43546 3102 43548
rect 3126 43546 3182 43548
rect 2886 43494 2932 43546
rect 2932 43494 2942 43546
rect 2966 43494 2996 43546
rect 2996 43494 3008 43546
rect 3008 43494 3022 43546
rect 3046 43494 3060 43546
rect 3060 43494 3072 43546
rect 3072 43494 3102 43546
rect 3126 43494 3136 43546
rect 3136 43494 3182 43546
rect 2886 43492 2942 43494
rect 2966 43492 3022 43494
rect 3046 43492 3102 43494
rect 3126 43492 3182 43494
rect 2886 42458 2942 42460
rect 2966 42458 3022 42460
rect 3046 42458 3102 42460
rect 3126 42458 3182 42460
rect 2886 42406 2932 42458
rect 2932 42406 2942 42458
rect 2966 42406 2996 42458
rect 2996 42406 3008 42458
rect 3008 42406 3022 42458
rect 3046 42406 3060 42458
rect 3060 42406 3072 42458
rect 3072 42406 3102 42458
rect 3126 42406 3136 42458
rect 3136 42406 3182 42458
rect 2886 42404 2942 42406
rect 2966 42404 3022 42406
rect 3046 42404 3102 42406
rect 3126 42404 3182 42406
rect 2886 41370 2942 41372
rect 2966 41370 3022 41372
rect 3046 41370 3102 41372
rect 3126 41370 3182 41372
rect 2886 41318 2932 41370
rect 2932 41318 2942 41370
rect 2966 41318 2996 41370
rect 2996 41318 3008 41370
rect 3008 41318 3022 41370
rect 3046 41318 3060 41370
rect 3060 41318 3072 41370
rect 3072 41318 3102 41370
rect 3126 41318 3136 41370
rect 3136 41318 3182 41370
rect 2886 41316 2942 41318
rect 2966 41316 3022 41318
rect 3046 41316 3102 41318
rect 3126 41316 3182 41318
rect 3238 41112 3294 41168
rect 2886 40282 2942 40284
rect 2966 40282 3022 40284
rect 3046 40282 3102 40284
rect 3126 40282 3182 40284
rect 2886 40230 2932 40282
rect 2932 40230 2942 40282
rect 2966 40230 2996 40282
rect 2996 40230 3008 40282
rect 3008 40230 3022 40282
rect 3046 40230 3060 40282
rect 3060 40230 3072 40282
rect 3072 40230 3102 40282
rect 3126 40230 3136 40282
rect 3136 40230 3182 40282
rect 2886 40228 2942 40230
rect 2966 40228 3022 40230
rect 3046 40228 3102 40230
rect 3126 40228 3182 40230
rect 2886 39194 2942 39196
rect 2966 39194 3022 39196
rect 3046 39194 3102 39196
rect 3126 39194 3182 39196
rect 2886 39142 2932 39194
rect 2932 39142 2942 39194
rect 2966 39142 2996 39194
rect 2996 39142 3008 39194
rect 3008 39142 3022 39194
rect 3046 39142 3060 39194
rect 3060 39142 3072 39194
rect 3072 39142 3102 39194
rect 3126 39142 3136 39194
rect 3136 39142 3182 39194
rect 2886 39140 2942 39142
rect 2966 39140 3022 39142
rect 3046 39140 3102 39142
rect 3126 39140 3182 39142
rect 3146 38936 3202 38992
rect 2886 38106 2942 38108
rect 2966 38106 3022 38108
rect 3046 38106 3102 38108
rect 3126 38106 3182 38108
rect 2886 38054 2932 38106
rect 2932 38054 2942 38106
rect 2966 38054 2996 38106
rect 2996 38054 3008 38106
rect 3008 38054 3022 38106
rect 3046 38054 3060 38106
rect 3060 38054 3072 38106
rect 3072 38054 3102 38106
rect 3126 38054 3136 38106
rect 3136 38054 3182 38106
rect 2886 38052 2942 38054
rect 2966 38052 3022 38054
rect 3046 38052 3102 38054
rect 3126 38052 3182 38054
rect 2886 37018 2942 37020
rect 2966 37018 3022 37020
rect 3046 37018 3102 37020
rect 3126 37018 3182 37020
rect 2886 36966 2932 37018
rect 2932 36966 2942 37018
rect 2966 36966 2996 37018
rect 2996 36966 3008 37018
rect 3008 36966 3022 37018
rect 3046 36966 3060 37018
rect 3060 36966 3072 37018
rect 3072 36966 3102 37018
rect 3126 36966 3136 37018
rect 3136 36966 3182 37018
rect 2886 36964 2942 36966
rect 2966 36964 3022 36966
rect 3046 36964 3102 36966
rect 3126 36964 3182 36966
rect 2886 35930 2942 35932
rect 2966 35930 3022 35932
rect 3046 35930 3102 35932
rect 3126 35930 3182 35932
rect 2886 35878 2932 35930
rect 2932 35878 2942 35930
rect 2966 35878 2996 35930
rect 2996 35878 3008 35930
rect 3008 35878 3022 35930
rect 3046 35878 3060 35930
rect 3060 35878 3072 35930
rect 3072 35878 3102 35930
rect 3126 35878 3136 35930
rect 3136 35878 3182 35930
rect 2886 35876 2942 35878
rect 2966 35876 3022 35878
rect 3046 35876 3102 35878
rect 3126 35876 3182 35878
rect 3514 41520 3570 41576
rect 3514 38612 3570 38668
rect 2886 34842 2942 34844
rect 2966 34842 3022 34844
rect 3046 34842 3102 34844
rect 3126 34842 3182 34844
rect 2886 34790 2932 34842
rect 2932 34790 2942 34842
rect 2966 34790 2996 34842
rect 2996 34790 3008 34842
rect 3008 34790 3022 34842
rect 3046 34790 3060 34842
rect 3060 34790 3072 34842
rect 3072 34790 3102 34842
rect 3126 34790 3136 34842
rect 3136 34790 3182 34842
rect 2886 34788 2942 34790
rect 2966 34788 3022 34790
rect 3046 34788 3102 34790
rect 3126 34788 3182 34790
rect 2886 33754 2942 33756
rect 2966 33754 3022 33756
rect 3046 33754 3102 33756
rect 3126 33754 3182 33756
rect 2886 33702 2932 33754
rect 2932 33702 2942 33754
rect 2966 33702 2996 33754
rect 2996 33702 3008 33754
rect 3008 33702 3022 33754
rect 3046 33702 3060 33754
rect 3060 33702 3072 33754
rect 3072 33702 3102 33754
rect 3126 33702 3136 33754
rect 3136 33702 3182 33754
rect 2886 33700 2942 33702
rect 2966 33700 3022 33702
rect 3046 33700 3102 33702
rect 3126 33700 3182 33702
rect 1858 31320 1914 31376
rect 2410 31184 2466 31240
rect 1921 31034 1977 31036
rect 2001 31034 2057 31036
rect 2081 31034 2137 31036
rect 2161 31034 2217 31036
rect 1921 30982 1967 31034
rect 1967 30982 1977 31034
rect 2001 30982 2031 31034
rect 2031 30982 2043 31034
rect 2043 30982 2057 31034
rect 2081 30982 2095 31034
rect 2095 30982 2107 31034
rect 2107 30982 2137 31034
rect 2161 30982 2171 31034
rect 2171 30982 2217 31034
rect 1921 30980 1977 30982
rect 2001 30980 2057 30982
rect 2081 30980 2137 30982
rect 2161 30980 2217 30982
rect 1921 29946 1977 29948
rect 2001 29946 2057 29948
rect 2081 29946 2137 29948
rect 2161 29946 2217 29948
rect 1921 29894 1967 29946
rect 1967 29894 1977 29946
rect 2001 29894 2031 29946
rect 2031 29894 2043 29946
rect 2043 29894 2057 29946
rect 2081 29894 2095 29946
rect 2095 29894 2107 29946
rect 2107 29894 2137 29946
rect 2161 29894 2171 29946
rect 2171 29894 2217 29946
rect 1921 29892 1977 29894
rect 2001 29892 2057 29894
rect 2081 29892 2137 29894
rect 2161 29892 2217 29894
rect 1921 28858 1977 28860
rect 2001 28858 2057 28860
rect 2081 28858 2137 28860
rect 2161 28858 2217 28860
rect 1921 28806 1967 28858
rect 1967 28806 1977 28858
rect 2001 28806 2031 28858
rect 2031 28806 2043 28858
rect 2043 28806 2057 28858
rect 2081 28806 2095 28858
rect 2095 28806 2107 28858
rect 2107 28806 2137 28858
rect 2161 28806 2171 28858
rect 2171 28806 2217 28858
rect 1921 28804 1977 28806
rect 2001 28804 2057 28806
rect 2081 28804 2137 28806
rect 2161 28804 2217 28806
rect 1921 27770 1977 27772
rect 2001 27770 2057 27772
rect 2081 27770 2137 27772
rect 2161 27770 2217 27772
rect 1921 27718 1967 27770
rect 1967 27718 1977 27770
rect 2001 27718 2031 27770
rect 2031 27718 2043 27770
rect 2043 27718 2057 27770
rect 2081 27718 2095 27770
rect 2095 27718 2107 27770
rect 2107 27718 2137 27770
rect 2161 27718 2171 27770
rect 2171 27718 2217 27770
rect 1921 27716 1977 27718
rect 2001 27716 2057 27718
rect 2081 27716 2137 27718
rect 2161 27716 2217 27718
rect 1582 26832 1638 26888
rect 1582 26016 1638 26072
rect 1921 26682 1977 26684
rect 2001 26682 2057 26684
rect 2081 26682 2137 26684
rect 2161 26682 2217 26684
rect 1921 26630 1967 26682
rect 1967 26630 1977 26682
rect 2001 26630 2031 26682
rect 2031 26630 2043 26682
rect 2043 26630 2057 26682
rect 2081 26630 2095 26682
rect 2095 26630 2107 26682
rect 2107 26630 2137 26682
rect 2161 26630 2171 26682
rect 2171 26630 2217 26682
rect 1921 26628 1977 26630
rect 2001 26628 2057 26630
rect 2081 26628 2137 26630
rect 2161 26628 2217 26630
rect 2886 32666 2942 32668
rect 2966 32666 3022 32668
rect 3046 32666 3102 32668
rect 3126 32666 3182 32668
rect 2886 32614 2932 32666
rect 2932 32614 2942 32666
rect 2966 32614 2996 32666
rect 2996 32614 3008 32666
rect 3008 32614 3022 32666
rect 3046 32614 3060 32666
rect 3060 32614 3072 32666
rect 3072 32614 3102 32666
rect 3126 32614 3136 32666
rect 3136 32614 3182 32666
rect 2886 32612 2942 32614
rect 2966 32612 3022 32614
rect 3046 32612 3102 32614
rect 3126 32612 3182 32614
rect 2886 31578 2942 31580
rect 2966 31578 3022 31580
rect 3046 31578 3102 31580
rect 3126 31578 3182 31580
rect 2886 31526 2932 31578
rect 2932 31526 2942 31578
rect 2966 31526 2996 31578
rect 2996 31526 3008 31578
rect 3008 31526 3022 31578
rect 3046 31526 3060 31578
rect 3060 31526 3072 31578
rect 3072 31526 3102 31578
rect 3126 31526 3136 31578
rect 3136 31526 3182 31578
rect 2886 31524 2942 31526
rect 2966 31524 3022 31526
rect 3046 31524 3102 31526
rect 3126 31524 3182 31526
rect 2886 30490 2942 30492
rect 2966 30490 3022 30492
rect 3046 30490 3102 30492
rect 3126 30490 3182 30492
rect 2886 30438 2932 30490
rect 2932 30438 2942 30490
rect 2966 30438 2996 30490
rect 2996 30438 3008 30490
rect 3008 30438 3022 30490
rect 3046 30438 3060 30490
rect 3060 30438 3072 30490
rect 3072 30438 3102 30490
rect 3126 30438 3136 30490
rect 3136 30438 3182 30490
rect 2886 30436 2942 30438
rect 2966 30436 3022 30438
rect 3046 30436 3102 30438
rect 3126 30436 3182 30438
rect 2870 29824 2926 29880
rect 2886 29402 2942 29404
rect 2966 29402 3022 29404
rect 3046 29402 3102 29404
rect 3126 29402 3182 29404
rect 2886 29350 2932 29402
rect 2932 29350 2942 29402
rect 2966 29350 2996 29402
rect 2996 29350 3008 29402
rect 3008 29350 3022 29402
rect 3046 29350 3060 29402
rect 3060 29350 3072 29402
rect 3072 29350 3102 29402
rect 3126 29350 3136 29402
rect 3136 29350 3182 29402
rect 2886 29348 2942 29350
rect 2966 29348 3022 29350
rect 3046 29348 3102 29350
rect 3126 29348 3182 29350
rect 3514 37848 3570 37904
rect 3852 51706 3908 51708
rect 3932 51706 3988 51708
rect 4012 51706 4068 51708
rect 4092 51706 4148 51708
rect 3852 51654 3898 51706
rect 3898 51654 3908 51706
rect 3932 51654 3962 51706
rect 3962 51654 3974 51706
rect 3974 51654 3988 51706
rect 4012 51654 4026 51706
rect 4026 51654 4038 51706
rect 4038 51654 4068 51706
rect 4092 51654 4102 51706
rect 4102 51654 4148 51706
rect 3852 51652 3908 51654
rect 3932 51652 3988 51654
rect 4012 51652 4068 51654
rect 4092 51652 4148 51654
rect 3852 50618 3908 50620
rect 3932 50618 3988 50620
rect 4012 50618 4068 50620
rect 4092 50618 4148 50620
rect 3852 50566 3898 50618
rect 3898 50566 3908 50618
rect 3932 50566 3962 50618
rect 3962 50566 3974 50618
rect 3974 50566 3988 50618
rect 4012 50566 4026 50618
rect 4026 50566 4038 50618
rect 4038 50566 4068 50618
rect 4092 50566 4102 50618
rect 4102 50566 4148 50618
rect 3852 50564 3908 50566
rect 3932 50564 3988 50566
rect 4012 50564 4068 50566
rect 4092 50564 4148 50566
rect 3852 49530 3908 49532
rect 3932 49530 3988 49532
rect 4012 49530 4068 49532
rect 4092 49530 4148 49532
rect 3852 49478 3898 49530
rect 3898 49478 3908 49530
rect 3932 49478 3962 49530
rect 3962 49478 3974 49530
rect 3974 49478 3988 49530
rect 4012 49478 4026 49530
rect 4026 49478 4038 49530
rect 4038 49478 4068 49530
rect 4092 49478 4102 49530
rect 4102 49478 4148 49530
rect 3852 49476 3908 49478
rect 3932 49476 3988 49478
rect 4012 49476 4068 49478
rect 4092 49476 4148 49478
rect 3852 48442 3908 48444
rect 3932 48442 3988 48444
rect 4012 48442 4068 48444
rect 4092 48442 4148 48444
rect 3852 48390 3898 48442
rect 3898 48390 3908 48442
rect 3932 48390 3962 48442
rect 3962 48390 3974 48442
rect 3974 48390 3988 48442
rect 4012 48390 4026 48442
rect 4026 48390 4038 48442
rect 4038 48390 4068 48442
rect 4092 48390 4102 48442
rect 4102 48390 4148 48442
rect 3852 48388 3908 48390
rect 3932 48388 3988 48390
rect 4012 48388 4068 48390
rect 4092 48388 4148 48390
rect 3852 47354 3908 47356
rect 3932 47354 3988 47356
rect 4012 47354 4068 47356
rect 4092 47354 4148 47356
rect 3852 47302 3898 47354
rect 3898 47302 3908 47354
rect 3932 47302 3962 47354
rect 3962 47302 3974 47354
rect 3974 47302 3988 47354
rect 4012 47302 4026 47354
rect 4026 47302 4038 47354
rect 4038 47302 4068 47354
rect 4092 47302 4102 47354
rect 4102 47302 4148 47354
rect 3852 47300 3908 47302
rect 3932 47300 3988 47302
rect 4012 47300 4068 47302
rect 4092 47300 4148 47302
rect 3852 46266 3908 46268
rect 3932 46266 3988 46268
rect 4012 46266 4068 46268
rect 4092 46266 4148 46268
rect 3852 46214 3898 46266
rect 3898 46214 3908 46266
rect 3932 46214 3962 46266
rect 3962 46214 3974 46266
rect 3974 46214 3988 46266
rect 4012 46214 4026 46266
rect 4026 46214 4038 46266
rect 4038 46214 4068 46266
rect 4092 46214 4102 46266
rect 4102 46214 4148 46266
rect 3852 46212 3908 46214
rect 3932 46212 3988 46214
rect 4012 46212 4068 46214
rect 4092 46212 4148 46214
rect 5446 57976 5502 58032
rect 6274 57432 6330 57488
rect 4817 56602 4873 56604
rect 4897 56602 4953 56604
rect 4977 56602 5033 56604
rect 5057 56602 5113 56604
rect 4817 56550 4863 56602
rect 4863 56550 4873 56602
rect 4897 56550 4927 56602
rect 4927 56550 4939 56602
rect 4939 56550 4953 56602
rect 4977 56550 4991 56602
rect 4991 56550 5003 56602
rect 5003 56550 5033 56602
rect 5057 56550 5067 56602
rect 5067 56550 5113 56602
rect 4817 56548 4873 56550
rect 4897 56548 4953 56550
rect 4977 56548 5033 56550
rect 5057 56548 5113 56550
rect 4817 55514 4873 55516
rect 4897 55514 4953 55516
rect 4977 55514 5033 55516
rect 5057 55514 5113 55516
rect 4817 55462 4863 55514
rect 4863 55462 4873 55514
rect 4897 55462 4927 55514
rect 4927 55462 4939 55514
rect 4939 55462 4953 55514
rect 4977 55462 4991 55514
rect 4991 55462 5003 55514
rect 5003 55462 5033 55514
rect 5057 55462 5067 55514
rect 5067 55462 5113 55514
rect 4817 55460 4873 55462
rect 4897 55460 4953 55462
rect 4977 55460 5033 55462
rect 5057 55460 5113 55462
rect 5782 57146 5838 57148
rect 5862 57146 5918 57148
rect 5942 57146 5998 57148
rect 6022 57146 6078 57148
rect 5782 57094 5828 57146
rect 5828 57094 5838 57146
rect 5862 57094 5892 57146
rect 5892 57094 5904 57146
rect 5904 57094 5918 57146
rect 5942 57094 5956 57146
rect 5956 57094 5968 57146
rect 5968 57094 5998 57146
rect 6022 57094 6032 57146
rect 6032 57094 6078 57146
rect 5782 57092 5838 57094
rect 5862 57092 5918 57094
rect 5942 57092 5998 57094
rect 6022 57092 6078 57094
rect 6182 56888 6238 56944
rect 5722 56228 5778 56264
rect 5722 56208 5724 56228
rect 5724 56208 5776 56228
rect 5776 56208 5778 56228
rect 5782 56058 5838 56060
rect 5862 56058 5918 56060
rect 5942 56058 5998 56060
rect 6022 56058 6078 56060
rect 5782 56006 5828 56058
rect 5828 56006 5838 56058
rect 5862 56006 5892 56058
rect 5892 56006 5904 56058
rect 5904 56006 5918 56058
rect 5942 56006 5956 56058
rect 5956 56006 5968 56058
rect 5968 56006 5998 56058
rect 6022 56006 6032 56058
rect 6032 56006 6078 56058
rect 5782 56004 5838 56006
rect 5862 56004 5918 56006
rect 5942 56004 5998 56006
rect 6022 56004 6078 56006
rect 5998 55664 6054 55720
rect 4342 47776 4398 47832
rect 3852 45178 3908 45180
rect 3932 45178 3988 45180
rect 4012 45178 4068 45180
rect 4092 45178 4148 45180
rect 3852 45126 3898 45178
rect 3898 45126 3908 45178
rect 3932 45126 3962 45178
rect 3962 45126 3974 45178
rect 3974 45126 3988 45178
rect 4012 45126 4026 45178
rect 4026 45126 4038 45178
rect 4038 45126 4068 45178
rect 4092 45126 4102 45178
rect 4102 45126 4148 45178
rect 3852 45124 3908 45126
rect 3932 45124 3988 45126
rect 4012 45124 4068 45126
rect 4092 45124 4148 45126
rect 3852 44090 3908 44092
rect 3932 44090 3988 44092
rect 4012 44090 4068 44092
rect 4092 44090 4148 44092
rect 3852 44038 3898 44090
rect 3898 44038 3908 44090
rect 3932 44038 3962 44090
rect 3962 44038 3974 44090
rect 3974 44038 3988 44090
rect 4012 44038 4026 44090
rect 4026 44038 4038 44090
rect 4038 44038 4068 44090
rect 4092 44038 4102 44090
rect 4102 44038 4148 44090
rect 3852 44036 3908 44038
rect 3932 44036 3988 44038
rect 4012 44036 4068 44038
rect 4092 44036 4148 44038
rect 3852 43002 3908 43004
rect 3932 43002 3988 43004
rect 4012 43002 4068 43004
rect 4092 43002 4148 43004
rect 3852 42950 3898 43002
rect 3898 42950 3908 43002
rect 3932 42950 3962 43002
rect 3962 42950 3974 43002
rect 3974 42950 3988 43002
rect 4012 42950 4026 43002
rect 4026 42950 4038 43002
rect 4038 42950 4068 43002
rect 4092 42950 4102 43002
rect 4102 42950 4148 43002
rect 3852 42948 3908 42950
rect 3932 42948 3988 42950
rect 4012 42948 4068 42950
rect 4092 42948 4148 42950
rect 3852 41914 3908 41916
rect 3932 41914 3988 41916
rect 4012 41914 4068 41916
rect 4092 41914 4148 41916
rect 3852 41862 3898 41914
rect 3898 41862 3908 41914
rect 3932 41862 3962 41914
rect 3962 41862 3974 41914
rect 3974 41862 3988 41914
rect 4012 41862 4026 41914
rect 4026 41862 4038 41914
rect 4038 41862 4068 41914
rect 4092 41862 4102 41914
rect 4102 41862 4148 41914
rect 3852 41860 3908 41862
rect 3932 41860 3988 41862
rect 4012 41860 4068 41862
rect 4092 41860 4148 41862
rect 4342 41656 4398 41712
rect 4817 54426 4873 54428
rect 4897 54426 4953 54428
rect 4977 54426 5033 54428
rect 5057 54426 5113 54428
rect 4817 54374 4863 54426
rect 4863 54374 4873 54426
rect 4897 54374 4927 54426
rect 4927 54374 4939 54426
rect 4939 54374 4953 54426
rect 4977 54374 4991 54426
rect 4991 54374 5003 54426
rect 5003 54374 5033 54426
rect 5057 54374 5067 54426
rect 5067 54374 5113 54426
rect 4817 54372 4873 54374
rect 4897 54372 4953 54374
rect 4977 54372 5033 54374
rect 5057 54372 5113 54374
rect 4817 53338 4873 53340
rect 4897 53338 4953 53340
rect 4977 53338 5033 53340
rect 5057 53338 5113 53340
rect 4817 53286 4863 53338
rect 4863 53286 4873 53338
rect 4897 53286 4927 53338
rect 4927 53286 4939 53338
rect 4939 53286 4953 53338
rect 4977 53286 4991 53338
rect 4991 53286 5003 53338
rect 5003 53286 5033 53338
rect 5057 53286 5067 53338
rect 5067 53286 5113 53338
rect 4817 53284 4873 53286
rect 4897 53284 4953 53286
rect 4977 53284 5033 53286
rect 5057 53284 5113 53286
rect 4817 52250 4873 52252
rect 4897 52250 4953 52252
rect 4977 52250 5033 52252
rect 5057 52250 5113 52252
rect 4817 52198 4863 52250
rect 4863 52198 4873 52250
rect 4897 52198 4927 52250
rect 4927 52198 4939 52250
rect 4939 52198 4953 52250
rect 4977 52198 4991 52250
rect 4991 52198 5003 52250
rect 5003 52198 5033 52250
rect 5057 52198 5067 52250
rect 5067 52198 5113 52250
rect 4817 52196 4873 52198
rect 4897 52196 4953 52198
rect 4977 52196 5033 52198
rect 5057 52196 5113 52198
rect 4817 51162 4873 51164
rect 4897 51162 4953 51164
rect 4977 51162 5033 51164
rect 5057 51162 5113 51164
rect 4817 51110 4863 51162
rect 4863 51110 4873 51162
rect 4897 51110 4927 51162
rect 4927 51110 4939 51162
rect 4939 51110 4953 51162
rect 4977 51110 4991 51162
rect 4991 51110 5003 51162
rect 5003 51110 5033 51162
rect 5057 51110 5067 51162
rect 5067 51110 5113 51162
rect 4817 51108 4873 51110
rect 4897 51108 4953 51110
rect 4977 51108 5033 51110
rect 5057 51108 5113 51110
rect 4817 50074 4873 50076
rect 4897 50074 4953 50076
rect 4977 50074 5033 50076
rect 5057 50074 5113 50076
rect 4817 50022 4863 50074
rect 4863 50022 4873 50074
rect 4897 50022 4927 50074
rect 4927 50022 4939 50074
rect 4939 50022 4953 50074
rect 4977 50022 4991 50074
rect 4991 50022 5003 50074
rect 5003 50022 5033 50074
rect 5057 50022 5067 50074
rect 5067 50022 5113 50074
rect 4817 50020 4873 50022
rect 4897 50020 4953 50022
rect 4977 50020 5033 50022
rect 5057 50020 5113 50022
rect 4817 48986 4873 48988
rect 4897 48986 4953 48988
rect 4977 48986 5033 48988
rect 5057 48986 5113 48988
rect 4817 48934 4863 48986
rect 4863 48934 4873 48986
rect 4897 48934 4927 48986
rect 4927 48934 4939 48986
rect 4939 48934 4953 48986
rect 4977 48934 4991 48986
rect 4991 48934 5003 48986
rect 5003 48934 5033 48986
rect 5057 48934 5067 48986
rect 5067 48934 5113 48986
rect 4817 48932 4873 48934
rect 4897 48932 4953 48934
rect 4977 48932 5033 48934
rect 5057 48932 5113 48934
rect 4802 48048 4858 48104
rect 4817 47898 4873 47900
rect 4897 47898 4953 47900
rect 4977 47898 5033 47900
rect 5057 47898 5113 47900
rect 4817 47846 4863 47898
rect 4863 47846 4873 47898
rect 4897 47846 4927 47898
rect 4927 47846 4939 47898
rect 4939 47846 4953 47898
rect 4977 47846 4991 47898
rect 4991 47846 5003 47898
rect 5003 47846 5033 47898
rect 5057 47846 5067 47898
rect 5067 47846 5113 47898
rect 4817 47844 4873 47846
rect 4897 47844 4953 47846
rect 4977 47844 5033 47846
rect 5057 47844 5113 47846
rect 4817 46810 4873 46812
rect 4897 46810 4953 46812
rect 4977 46810 5033 46812
rect 5057 46810 5113 46812
rect 4817 46758 4863 46810
rect 4863 46758 4873 46810
rect 4897 46758 4927 46810
rect 4927 46758 4939 46810
rect 4939 46758 4953 46810
rect 4977 46758 4991 46810
rect 4991 46758 5003 46810
rect 5003 46758 5033 46810
rect 5057 46758 5067 46810
rect 5067 46758 5113 46810
rect 4817 46756 4873 46758
rect 4897 46756 4953 46758
rect 4977 46756 5033 46758
rect 5057 46756 5113 46758
rect 4817 45722 4873 45724
rect 4897 45722 4953 45724
rect 4977 45722 5033 45724
rect 5057 45722 5113 45724
rect 4817 45670 4863 45722
rect 4863 45670 4873 45722
rect 4897 45670 4927 45722
rect 4927 45670 4939 45722
rect 4939 45670 4953 45722
rect 4977 45670 4991 45722
rect 4991 45670 5003 45722
rect 5003 45670 5033 45722
rect 5057 45670 5067 45722
rect 5067 45670 5113 45722
rect 4817 45668 4873 45670
rect 4897 45668 4953 45670
rect 4977 45668 5033 45670
rect 5057 45668 5113 45670
rect 4618 43288 4674 43344
rect 4817 44634 4873 44636
rect 4897 44634 4953 44636
rect 4977 44634 5033 44636
rect 5057 44634 5113 44636
rect 4817 44582 4863 44634
rect 4863 44582 4873 44634
rect 4897 44582 4927 44634
rect 4927 44582 4939 44634
rect 4939 44582 4953 44634
rect 4977 44582 4991 44634
rect 4991 44582 5003 44634
rect 5003 44582 5033 44634
rect 5057 44582 5067 44634
rect 5067 44582 5113 44634
rect 4817 44580 4873 44582
rect 4897 44580 4953 44582
rect 4977 44580 5033 44582
rect 5057 44580 5113 44582
rect 4817 43546 4873 43548
rect 4897 43546 4953 43548
rect 4977 43546 5033 43548
rect 5057 43546 5113 43548
rect 4817 43494 4863 43546
rect 4863 43494 4873 43546
rect 4897 43494 4927 43546
rect 4927 43494 4939 43546
rect 4939 43494 4953 43546
rect 4977 43494 4991 43546
rect 4991 43494 5003 43546
rect 5003 43494 5033 43546
rect 5057 43494 5067 43546
rect 5067 43494 5113 43546
rect 4817 43492 4873 43494
rect 4897 43492 4953 43494
rect 4977 43492 5033 43494
rect 5057 43492 5113 43494
rect 4817 42458 4873 42460
rect 4897 42458 4953 42460
rect 4977 42458 5033 42460
rect 5057 42458 5113 42460
rect 4817 42406 4863 42458
rect 4863 42406 4873 42458
rect 4897 42406 4927 42458
rect 4927 42406 4939 42458
rect 4939 42406 4953 42458
rect 4977 42406 4991 42458
rect 4991 42406 5003 42458
rect 5003 42406 5033 42458
rect 5057 42406 5067 42458
rect 5067 42406 5113 42458
rect 4817 42404 4873 42406
rect 4897 42404 4953 42406
rect 4977 42404 5033 42406
rect 5057 42404 5113 42406
rect 4802 42200 4858 42256
rect 4710 41928 4766 41984
rect 4526 41792 4582 41848
rect 4618 41656 4674 41712
rect 5722 55140 5778 55176
rect 5722 55120 5724 55140
rect 5724 55120 5776 55140
rect 5776 55120 5778 55140
rect 5782 54970 5838 54972
rect 5862 54970 5918 54972
rect 5942 54970 5998 54972
rect 6022 54970 6078 54972
rect 5782 54918 5828 54970
rect 5828 54918 5838 54970
rect 5862 54918 5892 54970
rect 5892 54918 5904 54970
rect 5904 54918 5918 54970
rect 5942 54918 5956 54970
rect 5956 54918 5968 54970
rect 5968 54918 5998 54970
rect 6022 54918 6032 54970
rect 6032 54918 6078 54970
rect 5782 54916 5838 54918
rect 5862 54916 5918 54918
rect 5942 54916 5998 54918
rect 6022 54916 6078 54918
rect 5998 54576 6054 54632
rect 5722 54052 5778 54088
rect 5722 54032 5724 54052
rect 5724 54032 5776 54052
rect 5776 54032 5778 54052
rect 5782 53882 5838 53884
rect 5862 53882 5918 53884
rect 5942 53882 5998 53884
rect 6022 53882 6078 53884
rect 5782 53830 5828 53882
rect 5828 53830 5838 53882
rect 5862 53830 5892 53882
rect 5892 53830 5904 53882
rect 5904 53830 5918 53882
rect 5942 53830 5956 53882
rect 5956 53830 5968 53882
rect 5968 53830 5998 53882
rect 6022 53830 6032 53882
rect 6032 53830 6078 53882
rect 5782 53828 5838 53830
rect 5862 53828 5918 53830
rect 5942 53828 5998 53830
rect 6022 53828 6078 53830
rect 5998 53488 6054 53544
rect 6182 52844 6184 52864
rect 6184 52844 6236 52864
rect 6236 52844 6238 52864
rect 6182 52808 6238 52844
rect 5782 52794 5838 52796
rect 5862 52794 5918 52796
rect 5942 52794 5998 52796
rect 6022 52794 6078 52796
rect 5782 52742 5828 52794
rect 5828 52742 5838 52794
rect 5862 52742 5892 52794
rect 5892 52742 5904 52794
rect 5904 52742 5918 52794
rect 5942 52742 5956 52794
rect 5956 52742 5968 52794
rect 5968 52742 5998 52794
rect 6022 52742 6032 52794
rect 6032 52742 6078 52794
rect 5782 52740 5838 52742
rect 5862 52740 5918 52742
rect 5942 52740 5998 52742
rect 6022 52740 6078 52742
rect 5998 52300 6000 52320
rect 6000 52300 6052 52320
rect 6052 52300 6054 52320
rect 5998 52264 6054 52300
rect 6182 51756 6184 51776
rect 6184 51756 6236 51776
rect 6236 51756 6238 51776
rect 6182 51720 6238 51756
rect 5782 51706 5838 51708
rect 5862 51706 5918 51708
rect 5942 51706 5998 51708
rect 6022 51706 6078 51708
rect 5782 51654 5828 51706
rect 5828 51654 5838 51706
rect 5862 51654 5892 51706
rect 5892 51654 5904 51706
rect 5904 51654 5918 51706
rect 5942 51654 5956 51706
rect 5956 51654 5968 51706
rect 5968 51654 5998 51706
rect 6022 51654 6032 51706
rect 6032 51654 6078 51706
rect 5782 51652 5838 51654
rect 5862 51652 5918 51654
rect 5942 51652 5998 51654
rect 6022 51652 6078 51654
rect 5998 51212 6000 51232
rect 6000 51212 6052 51232
rect 6052 51212 6054 51232
rect 5998 51176 6054 51212
rect 5262 42064 5318 42120
rect 4250 40840 4306 40896
rect 3852 40826 3908 40828
rect 3932 40826 3988 40828
rect 4012 40826 4068 40828
rect 4092 40826 4148 40828
rect 3852 40774 3898 40826
rect 3898 40774 3908 40826
rect 3932 40774 3962 40826
rect 3962 40774 3974 40826
rect 3974 40774 3988 40826
rect 4012 40774 4026 40826
rect 4026 40774 4038 40826
rect 4038 40774 4068 40826
rect 4092 40774 4102 40826
rect 4102 40774 4148 40826
rect 3852 40772 3908 40774
rect 3932 40772 3988 40774
rect 4012 40772 4068 40774
rect 4092 40772 4148 40774
rect 3852 39738 3908 39740
rect 3932 39738 3988 39740
rect 4012 39738 4068 39740
rect 4092 39738 4148 39740
rect 3852 39686 3898 39738
rect 3898 39686 3908 39738
rect 3932 39686 3962 39738
rect 3962 39686 3974 39738
rect 3974 39686 3988 39738
rect 4012 39686 4026 39738
rect 4026 39686 4038 39738
rect 4038 39686 4068 39738
rect 4092 39686 4102 39738
rect 4102 39686 4148 39738
rect 3852 39684 3908 39686
rect 3932 39684 3988 39686
rect 4012 39684 4068 39686
rect 4092 39684 4148 39686
rect 3852 38650 3908 38652
rect 3932 38650 3988 38652
rect 4012 38650 4068 38652
rect 4092 38650 4148 38652
rect 3852 38598 3898 38650
rect 3898 38598 3908 38650
rect 3932 38598 3962 38650
rect 3962 38598 3974 38650
rect 3974 38598 3988 38650
rect 4012 38598 4026 38650
rect 4026 38598 4038 38650
rect 4038 38598 4068 38650
rect 4092 38598 4102 38650
rect 4102 38598 4148 38650
rect 3852 38596 3908 38598
rect 3932 38596 3988 38598
rect 4012 38596 4068 38598
rect 4092 38596 4148 38598
rect 3852 37562 3908 37564
rect 3932 37562 3988 37564
rect 4012 37562 4068 37564
rect 4092 37562 4148 37564
rect 3852 37510 3898 37562
rect 3898 37510 3908 37562
rect 3932 37510 3962 37562
rect 3962 37510 3974 37562
rect 3974 37510 3988 37562
rect 4012 37510 4026 37562
rect 4026 37510 4038 37562
rect 4038 37510 4068 37562
rect 4092 37510 4102 37562
rect 4102 37510 4148 37562
rect 3852 37508 3908 37510
rect 3932 37508 3988 37510
rect 4012 37508 4068 37510
rect 4092 37508 4148 37510
rect 3852 36474 3908 36476
rect 3932 36474 3988 36476
rect 4012 36474 4068 36476
rect 4092 36474 4148 36476
rect 3852 36422 3898 36474
rect 3898 36422 3908 36474
rect 3932 36422 3962 36474
rect 3962 36422 3974 36474
rect 3974 36422 3988 36474
rect 4012 36422 4026 36474
rect 4026 36422 4038 36474
rect 4038 36422 4068 36474
rect 4092 36422 4102 36474
rect 4102 36422 4148 36474
rect 3852 36420 3908 36422
rect 3932 36420 3988 36422
rect 4012 36420 4068 36422
rect 4092 36420 4148 36422
rect 3852 35386 3908 35388
rect 3932 35386 3988 35388
rect 4012 35386 4068 35388
rect 4092 35386 4148 35388
rect 3852 35334 3898 35386
rect 3898 35334 3908 35386
rect 3932 35334 3962 35386
rect 3962 35334 3974 35386
rect 3974 35334 3988 35386
rect 4012 35334 4026 35386
rect 4026 35334 4038 35386
rect 4038 35334 4068 35386
rect 4092 35334 4102 35386
rect 4102 35334 4148 35386
rect 3852 35332 3908 35334
rect 3932 35332 3988 35334
rect 4012 35332 4068 35334
rect 4092 35332 4148 35334
rect 3852 34298 3908 34300
rect 3932 34298 3988 34300
rect 4012 34298 4068 34300
rect 4092 34298 4148 34300
rect 3852 34246 3898 34298
rect 3898 34246 3908 34298
rect 3932 34246 3962 34298
rect 3962 34246 3974 34298
rect 3974 34246 3988 34298
rect 4012 34246 4026 34298
rect 4026 34246 4038 34298
rect 4038 34246 4068 34298
rect 4092 34246 4102 34298
rect 4102 34246 4148 34298
rect 3852 34244 3908 34246
rect 3932 34244 3988 34246
rect 4012 34244 4068 34246
rect 4092 34244 4148 34246
rect 3852 33210 3908 33212
rect 3932 33210 3988 33212
rect 4012 33210 4068 33212
rect 4092 33210 4148 33212
rect 3852 33158 3898 33210
rect 3898 33158 3908 33210
rect 3932 33158 3962 33210
rect 3962 33158 3974 33210
rect 3974 33158 3988 33210
rect 4012 33158 4026 33210
rect 4026 33158 4038 33210
rect 4038 33158 4068 33210
rect 4092 33158 4102 33210
rect 4102 33158 4148 33210
rect 3852 33156 3908 33158
rect 3932 33156 3988 33158
rect 4012 33156 4068 33158
rect 4092 33156 4148 33158
rect 3852 32122 3908 32124
rect 3932 32122 3988 32124
rect 4012 32122 4068 32124
rect 4092 32122 4148 32124
rect 3852 32070 3898 32122
rect 3898 32070 3908 32122
rect 3932 32070 3962 32122
rect 3962 32070 3974 32122
rect 3974 32070 3988 32122
rect 4012 32070 4026 32122
rect 4026 32070 4038 32122
rect 4038 32070 4068 32122
rect 4092 32070 4102 32122
rect 4102 32070 4148 32122
rect 3852 32068 3908 32070
rect 3932 32068 3988 32070
rect 4012 32068 4068 32070
rect 4092 32068 4148 32070
rect 3852 31034 3908 31036
rect 3932 31034 3988 31036
rect 4012 31034 4068 31036
rect 4092 31034 4148 31036
rect 3852 30982 3898 31034
rect 3898 30982 3908 31034
rect 3932 30982 3962 31034
rect 3962 30982 3974 31034
rect 3974 30982 3988 31034
rect 4012 30982 4026 31034
rect 4026 30982 4038 31034
rect 4038 30982 4068 31034
rect 4092 30982 4102 31034
rect 4102 30982 4148 31034
rect 3852 30980 3908 30982
rect 3932 30980 3988 30982
rect 4012 30980 4068 30982
rect 4092 30980 4148 30982
rect 3852 29946 3908 29948
rect 3932 29946 3988 29948
rect 4012 29946 4068 29948
rect 4092 29946 4148 29948
rect 3852 29894 3898 29946
rect 3898 29894 3908 29946
rect 3932 29894 3962 29946
rect 3962 29894 3974 29946
rect 3974 29894 3988 29946
rect 4012 29894 4026 29946
rect 4026 29894 4038 29946
rect 4038 29894 4068 29946
rect 4092 29894 4102 29946
rect 4102 29894 4148 29946
rect 3852 29892 3908 29894
rect 3932 29892 3988 29894
rect 4012 29892 4068 29894
rect 4092 29892 4148 29894
rect 3852 28858 3908 28860
rect 3932 28858 3988 28860
rect 4012 28858 4068 28860
rect 4092 28858 4148 28860
rect 3852 28806 3898 28858
rect 3898 28806 3908 28858
rect 3932 28806 3962 28858
rect 3962 28806 3974 28858
rect 3974 28806 3988 28858
rect 4012 28806 4026 28858
rect 4026 28806 4038 28858
rect 4038 28806 4068 28858
rect 4092 28806 4102 28858
rect 4102 28806 4148 28858
rect 3852 28804 3908 28806
rect 3932 28804 3988 28806
rect 4012 28804 4068 28806
rect 4092 28804 4148 28806
rect 2886 28314 2942 28316
rect 2966 28314 3022 28316
rect 3046 28314 3102 28316
rect 3126 28314 3182 28316
rect 2886 28262 2932 28314
rect 2932 28262 2942 28314
rect 2966 28262 2996 28314
rect 2996 28262 3008 28314
rect 3008 28262 3022 28314
rect 3046 28262 3060 28314
rect 3060 28262 3072 28314
rect 3072 28262 3102 28314
rect 3126 28262 3136 28314
rect 3136 28262 3182 28314
rect 2886 28260 2942 28262
rect 2966 28260 3022 28262
rect 3046 28260 3102 28262
rect 3126 28260 3182 28262
rect 3852 27770 3908 27772
rect 3932 27770 3988 27772
rect 4012 27770 4068 27772
rect 4092 27770 4148 27772
rect 3852 27718 3898 27770
rect 3898 27718 3908 27770
rect 3932 27718 3962 27770
rect 3962 27718 3974 27770
rect 3974 27718 3988 27770
rect 4012 27718 4026 27770
rect 4026 27718 4038 27770
rect 4038 27718 4068 27770
rect 4092 27718 4102 27770
rect 4102 27718 4148 27770
rect 3852 27716 3908 27718
rect 3932 27716 3988 27718
rect 4012 27716 4068 27718
rect 4092 27716 4148 27718
rect 2778 27512 2834 27568
rect 2886 27226 2942 27228
rect 2966 27226 3022 27228
rect 3046 27226 3102 27228
rect 3126 27226 3182 27228
rect 2886 27174 2932 27226
rect 2932 27174 2942 27226
rect 2966 27174 2996 27226
rect 2996 27174 3008 27226
rect 3008 27174 3022 27226
rect 3046 27174 3060 27226
rect 3060 27174 3072 27226
rect 3072 27174 3102 27226
rect 3126 27174 3136 27226
rect 3136 27174 3182 27226
rect 2886 27172 2942 27174
rect 2966 27172 3022 27174
rect 3046 27172 3102 27174
rect 3126 27172 3182 27174
rect 3852 26682 3908 26684
rect 3932 26682 3988 26684
rect 4012 26682 4068 26684
rect 4092 26682 4148 26684
rect 3852 26630 3898 26682
rect 3898 26630 3908 26682
rect 3932 26630 3962 26682
rect 3962 26630 3974 26682
rect 3974 26630 3988 26682
rect 4012 26630 4026 26682
rect 4026 26630 4038 26682
rect 4038 26630 4068 26682
rect 4092 26630 4102 26682
rect 4102 26630 4148 26682
rect 3852 26628 3908 26630
rect 3932 26628 3988 26630
rect 4012 26628 4068 26630
rect 4092 26628 4148 26630
rect 1582 25336 1638 25392
rect 1582 24520 1638 24576
rect 1582 23840 1638 23896
rect 1582 23060 1584 23080
rect 1584 23060 1636 23080
rect 1636 23060 1638 23080
rect 1582 23024 1638 23060
rect 1582 22208 1638 22264
rect 1582 21528 1638 21584
rect 1582 20712 1638 20768
rect 2886 26138 2942 26140
rect 2966 26138 3022 26140
rect 3046 26138 3102 26140
rect 3126 26138 3182 26140
rect 2886 26086 2932 26138
rect 2932 26086 2942 26138
rect 2966 26086 2996 26138
rect 2996 26086 3008 26138
rect 3008 26086 3022 26138
rect 3046 26086 3060 26138
rect 3060 26086 3072 26138
rect 3072 26086 3102 26138
rect 3126 26086 3136 26138
rect 3136 26086 3182 26138
rect 2886 26084 2942 26086
rect 2966 26084 3022 26086
rect 3046 26084 3102 26086
rect 3126 26084 3182 26086
rect 1921 25594 1977 25596
rect 2001 25594 2057 25596
rect 2081 25594 2137 25596
rect 2161 25594 2217 25596
rect 1921 25542 1967 25594
rect 1967 25542 1977 25594
rect 2001 25542 2031 25594
rect 2031 25542 2043 25594
rect 2043 25542 2057 25594
rect 2081 25542 2095 25594
rect 2095 25542 2107 25594
rect 2107 25542 2137 25594
rect 2161 25542 2171 25594
rect 2171 25542 2217 25594
rect 1921 25540 1977 25542
rect 2001 25540 2057 25542
rect 2081 25540 2137 25542
rect 2161 25540 2217 25542
rect 2886 25050 2942 25052
rect 2966 25050 3022 25052
rect 3046 25050 3102 25052
rect 3126 25050 3182 25052
rect 2886 24998 2932 25050
rect 2932 24998 2942 25050
rect 2966 24998 2996 25050
rect 2996 24998 3008 25050
rect 3008 24998 3022 25050
rect 3046 24998 3060 25050
rect 3060 24998 3072 25050
rect 3072 24998 3102 25050
rect 3126 24998 3136 25050
rect 3136 24998 3182 25050
rect 2886 24996 2942 24998
rect 2966 24996 3022 24998
rect 3046 24996 3102 24998
rect 3126 24996 3182 24998
rect 1921 24506 1977 24508
rect 2001 24506 2057 24508
rect 2081 24506 2137 24508
rect 2161 24506 2217 24508
rect 1921 24454 1967 24506
rect 1967 24454 1977 24506
rect 2001 24454 2031 24506
rect 2031 24454 2043 24506
rect 2043 24454 2057 24506
rect 2081 24454 2095 24506
rect 2095 24454 2107 24506
rect 2107 24454 2137 24506
rect 2161 24454 2171 24506
rect 2171 24454 2217 24506
rect 1921 24452 1977 24454
rect 2001 24452 2057 24454
rect 2081 24452 2137 24454
rect 2161 24452 2217 24454
rect 1921 23418 1977 23420
rect 2001 23418 2057 23420
rect 2081 23418 2137 23420
rect 2161 23418 2217 23420
rect 1921 23366 1967 23418
rect 1967 23366 1977 23418
rect 2001 23366 2031 23418
rect 2031 23366 2043 23418
rect 2043 23366 2057 23418
rect 2081 23366 2095 23418
rect 2095 23366 2107 23418
rect 2107 23366 2137 23418
rect 2161 23366 2171 23418
rect 2171 23366 2217 23418
rect 1921 23364 1977 23366
rect 2001 23364 2057 23366
rect 2081 23364 2137 23366
rect 2161 23364 2217 23366
rect 1921 22330 1977 22332
rect 2001 22330 2057 22332
rect 2081 22330 2137 22332
rect 2161 22330 2217 22332
rect 1921 22278 1967 22330
rect 1967 22278 1977 22330
rect 2001 22278 2031 22330
rect 2031 22278 2043 22330
rect 2043 22278 2057 22330
rect 2081 22278 2095 22330
rect 2095 22278 2107 22330
rect 2107 22278 2137 22330
rect 2161 22278 2171 22330
rect 2171 22278 2217 22330
rect 1921 22276 1977 22278
rect 2001 22276 2057 22278
rect 2081 22276 2137 22278
rect 2161 22276 2217 22278
rect 2886 23962 2942 23964
rect 2966 23962 3022 23964
rect 3046 23962 3102 23964
rect 3126 23962 3182 23964
rect 2886 23910 2932 23962
rect 2932 23910 2942 23962
rect 2966 23910 2996 23962
rect 2996 23910 3008 23962
rect 3008 23910 3022 23962
rect 3046 23910 3060 23962
rect 3060 23910 3072 23962
rect 3072 23910 3102 23962
rect 3126 23910 3136 23962
rect 3136 23910 3182 23962
rect 2886 23908 2942 23910
rect 2966 23908 3022 23910
rect 3046 23908 3102 23910
rect 3126 23908 3182 23910
rect 2886 22874 2942 22876
rect 2966 22874 3022 22876
rect 3046 22874 3102 22876
rect 3126 22874 3182 22876
rect 2886 22822 2932 22874
rect 2932 22822 2942 22874
rect 2966 22822 2996 22874
rect 2996 22822 3008 22874
rect 3008 22822 3022 22874
rect 3046 22822 3060 22874
rect 3060 22822 3072 22874
rect 3072 22822 3102 22874
rect 3126 22822 3136 22874
rect 3136 22822 3182 22874
rect 2886 22820 2942 22822
rect 2966 22820 3022 22822
rect 3046 22820 3102 22822
rect 3126 22820 3182 22822
rect 2886 21786 2942 21788
rect 2966 21786 3022 21788
rect 3046 21786 3102 21788
rect 3126 21786 3182 21788
rect 2886 21734 2932 21786
rect 2932 21734 2942 21786
rect 2966 21734 2996 21786
rect 2996 21734 3008 21786
rect 3008 21734 3022 21786
rect 3046 21734 3060 21786
rect 3060 21734 3072 21786
rect 3072 21734 3102 21786
rect 3126 21734 3136 21786
rect 3136 21734 3182 21786
rect 2886 21732 2942 21734
rect 2966 21732 3022 21734
rect 3046 21732 3102 21734
rect 3126 21732 3182 21734
rect 1921 21242 1977 21244
rect 2001 21242 2057 21244
rect 2081 21242 2137 21244
rect 2161 21242 2217 21244
rect 1921 21190 1967 21242
rect 1967 21190 1977 21242
rect 2001 21190 2031 21242
rect 2031 21190 2043 21242
rect 2043 21190 2057 21242
rect 2081 21190 2095 21242
rect 2095 21190 2107 21242
rect 2107 21190 2137 21242
rect 2161 21190 2171 21242
rect 2171 21190 2217 21242
rect 1921 21188 1977 21190
rect 2001 21188 2057 21190
rect 2081 21188 2137 21190
rect 2161 21188 2217 21190
rect 2886 20698 2942 20700
rect 2966 20698 3022 20700
rect 3046 20698 3102 20700
rect 3126 20698 3182 20700
rect 2886 20646 2932 20698
rect 2932 20646 2942 20698
rect 2966 20646 2996 20698
rect 2996 20646 3008 20698
rect 3008 20646 3022 20698
rect 3046 20646 3060 20698
rect 3060 20646 3072 20698
rect 3072 20646 3102 20698
rect 3126 20646 3136 20698
rect 3136 20646 3182 20698
rect 2886 20644 2942 20646
rect 2966 20644 3022 20646
rect 3046 20644 3102 20646
rect 3126 20644 3182 20646
rect 1921 20154 1977 20156
rect 2001 20154 2057 20156
rect 2081 20154 2137 20156
rect 2161 20154 2217 20156
rect 1921 20102 1967 20154
rect 1967 20102 1977 20154
rect 2001 20102 2031 20154
rect 2031 20102 2043 20154
rect 2043 20102 2057 20154
rect 2081 20102 2095 20154
rect 2095 20102 2107 20154
rect 2107 20102 2137 20154
rect 2161 20102 2171 20154
rect 2171 20102 2217 20154
rect 1921 20100 1977 20102
rect 2001 20100 2057 20102
rect 2081 20100 2137 20102
rect 2161 20100 2217 20102
rect 1582 20032 1638 20088
rect 2886 19610 2942 19612
rect 2966 19610 3022 19612
rect 3046 19610 3102 19612
rect 3126 19610 3182 19612
rect 2886 19558 2932 19610
rect 2932 19558 2942 19610
rect 2966 19558 2996 19610
rect 2996 19558 3008 19610
rect 3008 19558 3022 19610
rect 3046 19558 3060 19610
rect 3060 19558 3072 19610
rect 3072 19558 3102 19610
rect 3126 19558 3136 19610
rect 3136 19558 3182 19610
rect 2886 19556 2942 19558
rect 2966 19556 3022 19558
rect 3046 19556 3102 19558
rect 3126 19556 3182 19558
rect 1582 19216 1638 19272
rect 1921 19066 1977 19068
rect 2001 19066 2057 19068
rect 2081 19066 2137 19068
rect 2161 19066 2217 19068
rect 1921 19014 1967 19066
rect 1967 19014 1977 19066
rect 2001 19014 2031 19066
rect 2031 19014 2043 19066
rect 2043 19014 2057 19066
rect 2081 19014 2095 19066
rect 2095 19014 2107 19066
rect 2107 19014 2137 19066
rect 2161 19014 2171 19066
rect 2171 19014 2217 19066
rect 1921 19012 1977 19014
rect 2001 19012 2057 19014
rect 2081 19012 2137 19014
rect 2161 19012 2217 19014
rect 2886 18522 2942 18524
rect 2966 18522 3022 18524
rect 3046 18522 3102 18524
rect 3126 18522 3182 18524
rect 2886 18470 2932 18522
rect 2932 18470 2942 18522
rect 2966 18470 2996 18522
rect 2996 18470 3008 18522
rect 3008 18470 3022 18522
rect 3046 18470 3060 18522
rect 3060 18470 3072 18522
rect 3072 18470 3102 18522
rect 3126 18470 3136 18522
rect 3136 18470 3182 18522
rect 2886 18468 2942 18470
rect 2966 18468 3022 18470
rect 3046 18468 3102 18470
rect 3126 18468 3182 18470
rect 1582 18400 1638 18456
rect 3852 25594 3908 25596
rect 3932 25594 3988 25596
rect 4012 25594 4068 25596
rect 4092 25594 4148 25596
rect 3852 25542 3898 25594
rect 3898 25542 3908 25594
rect 3932 25542 3962 25594
rect 3962 25542 3974 25594
rect 3974 25542 3988 25594
rect 4012 25542 4026 25594
rect 4026 25542 4038 25594
rect 4038 25542 4068 25594
rect 4092 25542 4102 25594
rect 4102 25542 4148 25594
rect 3852 25540 3908 25542
rect 3932 25540 3988 25542
rect 4012 25540 4068 25542
rect 4092 25540 4148 25542
rect 3852 24506 3908 24508
rect 3932 24506 3988 24508
rect 4012 24506 4068 24508
rect 4092 24506 4148 24508
rect 3852 24454 3898 24506
rect 3898 24454 3908 24506
rect 3932 24454 3962 24506
rect 3962 24454 3974 24506
rect 3974 24454 3988 24506
rect 4012 24454 4026 24506
rect 4026 24454 4038 24506
rect 4038 24454 4068 24506
rect 4092 24454 4102 24506
rect 4102 24454 4148 24506
rect 3852 24452 3908 24454
rect 3932 24452 3988 24454
rect 4012 24452 4068 24454
rect 4092 24452 4148 24454
rect 3852 23418 3908 23420
rect 3932 23418 3988 23420
rect 4012 23418 4068 23420
rect 4092 23418 4148 23420
rect 3852 23366 3898 23418
rect 3898 23366 3908 23418
rect 3932 23366 3962 23418
rect 3962 23366 3974 23418
rect 3974 23366 3988 23418
rect 4012 23366 4026 23418
rect 4026 23366 4038 23418
rect 4038 23366 4068 23418
rect 4092 23366 4102 23418
rect 4102 23366 4148 23418
rect 3852 23364 3908 23366
rect 3932 23364 3988 23366
rect 4012 23364 4068 23366
rect 4092 23364 4148 23366
rect 3852 22330 3908 22332
rect 3932 22330 3988 22332
rect 4012 22330 4068 22332
rect 4092 22330 4148 22332
rect 3852 22278 3898 22330
rect 3898 22278 3908 22330
rect 3932 22278 3962 22330
rect 3962 22278 3974 22330
rect 3974 22278 3988 22330
rect 4012 22278 4026 22330
rect 4026 22278 4038 22330
rect 4038 22278 4068 22330
rect 4092 22278 4102 22330
rect 4102 22278 4148 22330
rect 3852 22276 3908 22278
rect 3932 22276 3988 22278
rect 4012 22276 4068 22278
rect 4092 22276 4148 22278
rect 3852 21242 3908 21244
rect 3932 21242 3988 21244
rect 4012 21242 4068 21244
rect 4092 21242 4148 21244
rect 3852 21190 3898 21242
rect 3898 21190 3908 21242
rect 3932 21190 3962 21242
rect 3962 21190 3974 21242
rect 3974 21190 3988 21242
rect 4012 21190 4026 21242
rect 4026 21190 4038 21242
rect 4038 21190 4068 21242
rect 4092 21190 4102 21242
rect 4102 21190 4148 21242
rect 3852 21188 3908 21190
rect 3932 21188 3988 21190
rect 4012 21188 4068 21190
rect 4092 21188 4148 21190
rect 3852 20154 3908 20156
rect 3932 20154 3988 20156
rect 4012 20154 4068 20156
rect 4092 20154 4148 20156
rect 3852 20102 3898 20154
rect 3898 20102 3908 20154
rect 3932 20102 3962 20154
rect 3962 20102 3974 20154
rect 3974 20102 3988 20154
rect 4012 20102 4026 20154
rect 4026 20102 4038 20154
rect 4038 20102 4068 20154
rect 4092 20102 4102 20154
rect 4102 20102 4148 20154
rect 3852 20100 3908 20102
rect 3932 20100 3988 20102
rect 4012 20100 4068 20102
rect 4092 20100 4148 20102
rect 3852 19066 3908 19068
rect 3932 19066 3988 19068
rect 4012 19066 4068 19068
rect 4092 19066 4148 19068
rect 3852 19014 3898 19066
rect 3898 19014 3908 19066
rect 3932 19014 3962 19066
rect 3962 19014 3974 19066
rect 3974 19014 3988 19066
rect 4012 19014 4026 19066
rect 4026 19014 4038 19066
rect 4038 19014 4068 19066
rect 4092 19014 4102 19066
rect 4102 19014 4148 19066
rect 3852 19012 3908 19014
rect 3932 19012 3988 19014
rect 4012 19012 4068 19014
rect 4092 19012 4148 19014
rect 1921 17978 1977 17980
rect 2001 17978 2057 17980
rect 2081 17978 2137 17980
rect 2161 17978 2217 17980
rect 1921 17926 1967 17978
rect 1967 17926 1977 17978
rect 2001 17926 2031 17978
rect 2031 17926 2043 17978
rect 2043 17926 2057 17978
rect 2081 17926 2095 17978
rect 2095 17926 2107 17978
rect 2107 17926 2137 17978
rect 2161 17926 2171 17978
rect 2171 17926 2217 17978
rect 1921 17924 1977 17926
rect 2001 17924 2057 17926
rect 2081 17924 2137 17926
rect 2161 17924 2217 17926
rect 3852 17978 3908 17980
rect 3932 17978 3988 17980
rect 4012 17978 4068 17980
rect 4092 17978 4148 17980
rect 3852 17926 3898 17978
rect 3898 17926 3908 17978
rect 3932 17926 3962 17978
rect 3962 17926 3974 17978
rect 3974 17926 3988 17978
rect 4012 17926 4026 17978
rect 4026 17926 4038 17978
rect 4038 17926 4068 17978
rect 4092 17926 4102 17978
rect 4102 17926 4148 17978
rect 3852 17924 3908 17926
rect 3932 17924 3988 17926
rect 4012 17924 4068 17926
rect 4092 17924 4148 17926
rect 1582 17720 1638 17776
rect 2886 17434 2942 17436
rect 2966 17434 3022 17436
rect 3046 17434 3102 17436
rect 3126 17434 3182 17436
rect 2886 17382 2932 17434
rect 2932 17382 2942 17434
rect 2966 17382 2996 17434
rect 2996 17382 3008 17434
rect 3008 17382 3022 17434
rect 3046 17382 3060 17434
rect 3060 17382 3072 17434
rect 3072 17382 3102 17434
rect 3126 17382 3136 17434
rect 3136 17382 3182 17434
rect 2886 17380 2942 17382
rect 2966 17380 3022 17382
rect 3046 17380 3102 17382
rect 3126 17380 3182 17382
rect 4434 41112 4490 41168
rect 4342 34448 4398 34504
rect 1582 16904 1638 16960
rect 1921 16890 1977 16892
rect 2001 16890 2057 16892
rect 2081 16890 2137 16892
rect 2161 16890 2217 16892
rect 1921 16838 1967 16890
rect 1967 16838 1977 16890
rect 2001 16838 2031 16890
rect 2031 16838 2043 16890
rect 2043 16838 2057 16890
rect 2081 16838 2095 16890
rect 2095 16838 2107 16890
rect 2107 16838 2137 16890
rect 2161 16838 2171 16890
rect 2171 16838 2217 16890
rect 1921 16836 1977 16838
rect 2001 16836 2057 16838
rect 2081 16836 2137 16838
rect 2161 16836 2217 16838
rect 3852 16890 3908 16892
rect 3932 16890 3988 16892
rect 4012 16890 4068 16892
rect 4092 16890 4148 16892
rect 3852 16838 3898 16890
rect 3898 16838 3908 16890
rect 3932 16838 3962 16890
rect 3962 16838 3974 16890
rect 3974 16838 3988 16890
rect 4012 16838 4026 16890
rect 4026 16838 4038 16890
rect 4038 16838 4068 16890
rect 4092 16838 4102 16890
rect 4102 16838 4148 16890
rect 3852 16836 3908 16838
rect 3932 16836 3988 16838
rect 4012 16836 4068 16838
rect 4092 16836 4148 16838
rect 4817 41370 4873 41372
rect 4897 41370 4953 41372
rect 4977 41370 5033 41372
rect 5057 41370 5113 41372
rect 4817 41318 4863 41370
rect 4863 41318 4873 41370
rect 4897 41318 4927 41370
rect 4927 41318 4939 41370
rect 4939 41318 4953 41370
rect 4977 41318 4991 41370
rect 4991 41318 5003 41370
rect 5003 41318 5033 41370
rect 5057 41318 5067 41370
rect 5067 41318 5113 41370
rect 4817 41316 4873 41318
rect 4897 41316 4953 41318
rect 4977 41316 5033 41318
rect 5057 41316 5113 41318
rect 5262 41556 5264 41576
rect 5264 41556 5316 41576
rect 5316 41556 5318 41576
rect 5262 41520 5318 41556
rect 4986 41012 4988 41032
rect 4988 41012 5040 41032
rect 5040 41012 5042 41032
rect 4986 40976 5042 41012
rect 4817 40282 4873 40284
rect 4897 40282 4953 40284
rect 4977 40282 5033 40284
rect 5057 40282 5113 40284
rect 4817 40230 4863 40282
rect 4863 40230 4873 40282
rect 4897 40230 4927 40282
rect 4927 40230 4939 40282
rect 4939 40230 4953 40282
rect 4977 40230 4991 40282
rect 4991 40230 5003 40282
rect 5003 40230 5033 40282
rect 5057 40230 5067 40282
rect 5067 40230 5113 40282
rect 4817 40228 4873 40230
rect 4897 40228 4953 40230
rect 4977 40228 5033 40230
rect 5057 40228 5113 40230
rect 4817 39194 4873 39196
rect 4897 39194 4953 39196
rect 4977 39194 5033 39196
rect 5057 39194 5113 39196
rect 4817 39142 4863 39194
rect 4863 39142 4873 39194
rect 4897 39142 4927 39194
rect 4927 39142 4939 39194
rect 4939 39142 4953 39194
rect 4977 39142 4991 39194
rect 4991 39142 5003 39194
rect 5003 39142 5033 39194
rect 5057 39142 5067 39194
rect 5067 39142 5113 39194
rect 4817 39140 4873 39142
rect 4897 39140 4953 39142
rect 4977 39140 5033 39142
rect 5057 39140 5113 39142
rect 5078 38936 5134 38992
rect 5078 38256 5134 38312
rect 4817 38106 4873 38108
rect 4897 38106 4953 38108
rect 4977 38106 5033 38108
rect 5057 38106 5113 38108
rect 4817 38054 4863 38106
rect 4863 38054 4873 38106
rect 4897 38054 4927 38106
rect 4927 38054 4939 38106
rect 4939 38054 4953 38106
rect 4977 38054 4991 38106
rect 4991 38054 5003 38106
rect 5003 38054 5033 38106
rect 5057 38054 5067 38106
rect 5067 38054 5113 38106
rect 4817 38052 4873 38054
rect 4897 38052 4953 38054
rect 4977 38052 5033 38054
rect 5057 38052 5113 38054
rect 4986 37748 4988 37768
rect 4988 37748 5040 37768
rect 5040 37748 5042 37768
rect 4986 37712 5042 37748
rect 4817 37018 4873 37020
rect 4897 37018 4953 37020
rect 4977 37018 5033 37020
rect 5057 37018 5113 37020
rect 4817 36966 4863 37018
rect 4863 36966 4873 37018
rect 4897 36966 4927 37018
rect 4927 36966 4939 37018
rect 4939 36966 4953 37018
rect 4977 36966 4991 37018
rect 4991 36966 5003 37018
rect 5003 36966 5033 37018
rect 5057 36966 5067 37018
rect 5067 36966 5113 37018
rect 4817 36964 4873 36966
rect 4897 36964 4953 36966
rect 4977 36964 5033 36966
rect 5057 36964 5113 36966
rect 4986 36660 4988 36680
rect 4988 36660 5040 36680
rect 5040 36660 5042 36680
rect 4986 36624 5042 36660
rect 4817 35930 4873 35932
rect 4897 35930 4953 35932
rect 4977 35930 5033 35932
rect 5057 35930 5113 35932
rect 4817 35878 4863 35930
rect 4863 35878 4873 35930
rect 4897 35878 4927 35930
rect 4927 35878 4939 35930
rect 4939 35878 4953 35930
rect 4977 35878 4991 35930
rect 4991 35878 5003 35930
rect 5003 35878 5033 35930
rect 5057 35878 5067 35930
rect 5067 35878 5113 35930
rect 4817 35876 4873 35878
rect 4897 35876 4953 35878
rect 4977 35876 5033 35878
rect 5057 35876 5113 35878
rect 5262 37032 5318 37088
rect 5262 35944 5318 36000
rect 4986 35572 4988 35592
rect 4988 35572 5040 35592
rect 5040 35572 5042 35592
rect 4986 35536 5042 35572
rect 4817 34842 4873 34844
rect 4897 34842 4953 34844
rect 4977 34842 5033 34844
rect 5057 34842 5113 34844
rect 4817 34790 4863 34842
rect 4863 34790 4873 34842
rect 4897 34790 4927 34842
rect 4927 34790 4939 34842
rect 4939 34790 4953 34842
rect 4977 34790 4991 34842
rect 4991 34790 5003 34842
rect 5003 34790 5033 34842
rect 5057 34790 5067 34842
rect 5067 34790 5113 34842
rect 4817 34788 4873 34790
rect 4897 34788 4953 34790
rect 4977 34788 5033 34790
rect 5057 34788 5113 34790
rect 4986 34484 4988 34504
rect 4988 34484 5040 34504
rect 5040 34484 5042 34504
rect 4986 34448 5042 34484
rect 4817 33754 4873 33756
rect 4897 33754 4953 33756
rect 4977 33754 5033 33756
rect 5057 33754 5113 33756
rect 4817 33702 4863 33754
rect 4863 33702 4873 33754
rect 4897 33702 4927 33754
rect 4927 33702 4939 33754
rect 4939 33702 4953 33754
rect 4977 33702 4991 33754
rect 4991 33702 5003 33754
rect 5003 33702 5033 33754
rect 5057 33702 5067 33754
rect 5067 33702 5113 33754
rect 4817 33700 4873 33702
rect 4897 33700 4953 33702
rect 4977 33700 5033 33702
rect 5057 33700 5113 33702
rect 4986 32952 5042 33008
rect 4817 32666 4873 32668
rect 4897 32666 4953 32668
rect 4977 32666 5033 32668
rect 5057 32666 5113 32668
rect 4817 32614 4863 32666
rect 4863 32614 4873 32666
rect 4897 32614 4927 32666
rect 4927 32614 4939 32666
rect 4939 32614 4953 32666
rect 4977 32614 4991 32666
rect 4991 32614 5003 32666
rect 5003 32614 5033 32666
rect 5057 32614 5067 32666
rect 5067 32614 5113 32666
rect 4817 32612 4873 32614
rect 4897 32612 4953 32614
rect 4977 32612 5033 32614
rect 5057 32612 5113 32614
rect 5262 34720 5318 34776
rect 5262 33632 5318 33688
rect 6366 50668 6368 50688
rect 6368 50668 6420 50688
rect 6420 50668 6422 50688
rect 6366 50632 6422 50668
rect 5782 50618 5838 50620
rect 5862 50618 5918 50620
rect 5942 50618 5998 50620
rect 6022 50618 6078 50620
rect 5782 50566 5828 50618
rect 5828 50566 5838 50618
rect 5862 50566 5892 50618
rect 5892 50566 5904 50618
rect 5904 50566 5918 50618
rect 5942 50566 5956 50618
rect 5956 50566 5968 50618
rect 5968 50566 5998 50618
rect 6022 50566 6032 50618
rect 6032 50566 6078 50618
rect 5782 50564 5838 50566
rect 5862 50564 5918 50566
rect 5942 50564 5998 50566
rect 6022 50564 6078 50566
rect 5998 50124 6000 50144
rect 6000 50124 6052 50144
rect 6052 50124 6054 50144
rect 5998 50088 6054 50124
rect 5782 49530 5838 49532
rect 5862 49530 5918 49532
rect 5942 49530 5998 49532
rect 6022 49530 6078 49532
rect 5782 49478 5828 49530
rect 5828 49478 5838 49530
rect 5862 49478 5892 49530
rect 5892 49478 5904 49530
rect 5904 49478 5918 49530
rect 5942 49478 5956 49530
rect 5956 49478 5968 49530
rect 5968 49478 5998 49530
rect 6022 49478 6032 49530
rect 6032 49478 6078 49530
rect 5782 49476 5838 49478
rect 5862 49476 5918 49478
rect 5942 49476 5998 49478
rect 6022 49476 6078 49478
rect 6182 49408 6238 49464
rect 5998 48864 6054 48920
rect 5782 48442 5838 48444
rect 5862 48442 5918 48444
rect 5942 48442 5998 48444
rect 6022 48442 6078 48444
rect 5782 48390 5828 48442
rect 5828 48390 5838 48442
rect 5862 48390 5892 48442
rect 5892 48390 5904 48442
rect 5904 48390 5918 48442
rect 5942 48390 5956 48442
rect 5956 48390 5968 48442
rect 5968 48390 5998 48442
rect 6022 48390 6032 48442
rect 6032 48390 6078 48442
rect 5782 48388 5838 48390
rect 5862 48388 5918 48390
rect 5942 48388 5998 48390
rect 6022 48388 6078 48390
rect 6182 48320 6238 48376
rect 5998 47776 6054 47832
rect 5782 47354 5838 47356
rect 5862 47354 5918 47356
rect 5942 47354 5998 47356
rect 6022 47354 6078 47356
rect 5782 47302 5828 47354
rect 5828 47302 5838 47354
rect 5862 47302 5892 47354
rect 5892 47302 5904 47354
rect 5904 47302 5918 47354
rect 5942 47302 5956 47354
rect 5956 47302 5968 47354
rect 5968 47302 5998 47354
rect 6022 47302 6032 47354
rect 6032 47302 6078 47354
rect 5782 47300 5838 47302
rect 5862 47300 5918 47302
rect 5942 47300 5998 47302
rect 6022 47300 6078 47302
rect 6182 47232 6238 47288
rect 5998 46688 6054 46744
rect 5782 46266 5838 46268
rect 5862 46266 5918 46268
rect 5942 46266 5998 46268
rect 6022 46266 6078 46268
rect 5782 46214 5828 46266
rect 5828 46214 5838 46266
rect 5862 46214 5892 46266
rect 5892 46214 5904 46266
rect 5904 46214 5918 46266
rect 5942 46214 5956 46266
rect 5956 46214 5968 46266
rect 5968 46214 5998 46266
rect 6022 46214 6032 46266
rect 6032 46214 6078 46266
rect 5782 46212 5838 46214
rect 5862 46212 5918 46214
rect 5942 46212 5998 46214
rect 6022 46212 6078 46214
rect 6182 46008 6238 46064
rect 5998 45464 6054 45520
rect 5814 45328 5870 45384
rect 5782 45178 5838 45180
rect 5862 45178 5918 45180
rect 5942 45178 5998 45180
rect 6022 45178 6078 45180
rect 5782 45126 5828 45178
rect 5828 45126 5838 45178
rect 5862 45126 5892 45178
rect 5892 45126 5904 45178
rect 5904 45126 5918 45178
rect 5942 45126 5956 45178
rect 5956 45126 5968 45178
rect 5968 45126 5998 45178
rect 6022 45126 6032 45178
rect 6032 45126 6078 45178
rect 5782 45124 5838 45126
rect 5862 45124 5918 45126
rect 5942 45124 5998 45126
rect 6022 45124 6078 45126
rect 6182 44920 6238 44976
rect 5998 44376 6054 44432
rect 5782 44090 5838 44092
rect 5862 44090 5918 44092
rect 5942 44090 5998 44092
rect 6022 44090 6078 44092
rect 5782 44038 5828 44090
rect 5828 44038 5838 44090
rect 5862 44038 5892 44090
rect 5892 44038 5904 44090
rect 5904 44038 5918 44090
rect 5942 44038 5956 44090
rect 5956 44038 5968 44090
rect 5968 44038 5998 44090
rect 6022 44038 6032 44090
rect 6032 44038 6078 44090
rect 5782 44036 5838 44038
rect 5862 44036 5918 44038
rect 5942 44036 5998 44038
rect 6022 44036 6078 44038
rect 5630 43832 5686 43888
rect 5998 43288 6054 43344
rect 5782 43002 5838 43004
rect 5862 43002 5918 43004
rect 5942 43002 5998 43004
rect 6022 43002 6078 43004
rect 5782 42950 5828 43002
rect 5828 42950 5838 43002
rect 5862 42950 5892 43002
rect 5892 42950 5904 43002
rect 5904 42950 5918 43002
rect 5942 42950 5956 43002
rect 5956 42950 5968 43002
rect 5968 42950 5998 43002
rect 6022 42950 6032 43002
rect 6032 42950 6078 43002
rect 5782 42948 5838 42950
rect 5862 42948 5918 42950
rect 5942 42948 5998 42950
rect 6022 42948 6078 42950
rect 5630 42744 5686 42800
rect 5262 32544 5318 32600
rect 4986 31864 5042 31920
rect 4817 31578 4873 31580
rect 4897 31578 4953 31580
rect 4977 31578 5033 31580
rect 5057 31578 5113 31580
rect 4817 31526 4863 31578
rect 4863 31526 4873 31578
rect 4897 31526 4927 31578
rect 4927 31526 4939 31578
rect 4939 31526 4953 31578
rect 4977 31526 4991 31578
rect 4991 31526 5003 31578
rect 5003 31526 5033 31578
rect 5057 31526 5067 31578
rect 5067 31526 5113 31578
rect 4817 31524 4873 31526
rect 4897 31524 4953 31526
rect 4977 31524 5033 31526
rect 5057 31524 5113 31526
rect 5722 42084 5778 42120
rect 5722 42064 5724 42084
rect 5724 42064 5776 42084
rect 5776 42064 5778 42084
rect 5782 41914 5838 41916
rect 5862 41914 5918 41916
rect 5942 41914 5998 41916
rect 6022 41914 6078 41916
rect 5782 41862 5828 41914
rect 5828 41862 5838 41914
rect 5862 41862 5892 41914
rect 5892 41862 5904 41914
rect 5904 41862 5918 41914
rect 5942 41862 5956 41914
rect 5956 41862 5968 41914
rect 5968 41862 5998 41914
rect 6022 41862 6032 41914
rect 6032 41862 6078 41914
rect 5782 41860 5838 41862
rect 5862 41860 5918 41862
rect 5942 41860 5998 41862
rect 6022 41860 6078 41862
rect 5782 40826 5838 40828
rect 5862 40826 5918 40828
rect 5942 40826 5998 40828
rect 6022 40826 6078 40828
rect 5782 40774 5828 40826
rect 5828 40774 5838 40826
rect 5862 40774 5892 40826
rect 5892 40774 5904 40826
rect 5904 40774 5918 40826
rect 5942 40774 5956 40826
rect 5956 40774 5968 40826
rect 5968 40774 5998 40826
rect 6022 40774 6032 40826
rect 6032 40774 6078 40826
rect 5782 40772 5838 40774
rect 5862 40772 5918 40774
rect 5942 40772 5998 40774
rect 6022 40772 6078 40774
rect 5722 40468 5724 40488
rect 5724 40468 5776 40488
rect 5776 40468 5778 40488
rect 5722 40432 5778 40468
rect 5814 39888 5870 39944
rect 5782 39738 5838 39740
rect 5862 39738 5918 39740
rect 5942 39738 5998 39740
rect 6022 39738 6078 39740
rect 5782 39686 5828 39738
rect 5828 39686 5838 39738
rect 5862 39686 5892 39738
rect 5892 39686 5904 39738
rect 5904 39686 5918 39738
rect 5942 39686 5956 39738
rect 5956 39686 5968 39738
rect 5968 39686 5998 39738
rect 6022 39686 6032 39738
rect 6032 39686 6078 39738
rect 5782 39684 5838 39686
rect 5862 39684 5918 39686
rect 5942 39684 5998 39686
rect 6022 39684 6078 39686
rect 6090 39380 6092 39400
rect 6092 39380 6144 39400
rect 6144 39380 6146 39400
rect 6090 39344 6146 39380
rect 6182 38664 6238 38720
rect 5782 38650 5838 38652
rect 5862 38650 5918 38652
rect 5942 38650 5998 38652
rect 6022 38650 6078 38652
rect 5782 38598 5828 38650
rect 5828 38598 5838 38650
rect 5862 38598 5892 38650
rect 5892 38598 5904 38650
rect 5904 38598 5918 38650
rect 5942 38598 5956 38650
rect 5956 38598 5968 38650
rect 5968 38598 5998 38650
rect 6022 38598 6032 38650
rect 6032 38598 6078 38650
rect 5782 38596 5838 38598
rect 5862 38596 5918 38598
rect 5942 38596 5998 38598
rect 6022 38596 6078 38598
rect 5630 38392 5686 38448
rect 5354 32272 5410 32328
rect 5354 31728 5410 31784
rect 4817 30490 4873 30492
rect 4897 30490 4953 30492
rect 4977 30490 5033 30492
rect 5057 30490 5113 30492
rect 4817 30438 4863 30490
rect 4863 30438 4873 30490
rect 4897 30438 4927 30490
rect 4927 30438 4939 30490
rect 4939 30438 4953 30490
rect 4977 30438 4991 30490
rect 4991 30438 5003 30490
rect 5003 30438 5033 30490
rect 5057 30438 5067 30490
rect 5067 30438 5113 30490
rect 4817 30436 4873 30438
rect 4897 30436 4953 30438
rect 4977 30436 5033 30438
rect 5057 30436 5113 30438
rect 4817 29402 4873 29404
rect 4897 29402 4953 29404
rect 4977 29402 5033 29404
rect 5057 29402 5113 29404
rect 4817 29350 4863 29402
rect 4863 29350 4873 29402
rect 4897 29350 4927 29402
rect 4927 29350 4939 29402
rect 4939 29350 4953 29402
rect 4977 29350 4991 29402
rect 4991 29350 5003 29402
rect 5003 29350 5033 29402
rect 5057 29350 5067 29402
rect 5067 29350 5113 29402
rect 4817 29348 4873 29350
rect 4897 29348 4953 29350
rect 4977 29348 5033 29350
rect 5057 29348 5113 29350
rect 6090 38120 6146 38176
rect 5782 37562 5838 37564
rect 5862 37562 5918 37564
rect 5942 37562 5998 37564
rect 6022 37562 6078 37564
rect 5782 37510 5828 37562
rect 5828 37510 5838 37562
rect 5862 37510 5892 37562
rect 5892 37510 5904 37562
rect 5904 37510 5918 37562
rect 5942 37510 5956 37562
rect 5956 37510 5968 37562
rect 5968 37510 5998 37562
rect 6022 37510 6032 37562
rect 6032 37510 6078 37562
rect 5782 37508 5838 37510
rect 5862 37508 5918 37510
rect 5942 37508 5998 37510
rect 6022 37508 6078 37510
rect 5782 36474 5838 36476
rect 5862 36474 5918 36476
rect 5942 36474 5998 36476
rect 6022 36474 6078 36476
rect 5782 36422 5828 36474
rect 5828 36422 5838 36474
rect 5862 36422 5892 36474
rect 5892 36422 5904 36474
rect 5904 36422 5918 36474
rect 5942 36422 5956 36474
rect 5956 36422 5968 36474
rect 5968 36422 5998 36474
rect 6022 36422 6032 36474
rect 6032 36422 6078 36474
rect 5782 36420 5838 36422
rect 5862 36420 5918 36422
rect 5942 36420 5998 36422
rect 6022 36420 6078 36422
rect 5782 35386 5838 35388
rect 5862 35386 5918 35388
rect 5942 35386 5998 35388
rect 6022 35386 6078 35388
rect 5782 35334 5828 35386
rect 5828 35334 5838 35386
rect 5862 35334 5892 35386
rect 5892 35334 5904 35386
rect 5904 35334 5918 35386
rect 5942 35334 5956 35386
rect 5956 35334 5968 35386
rect 5968 35334 5998 35386
rect 6022 35334 6032 35386
rect 6032 35334 6078 35386
rect 5782 35332 5838 35334
rect 5862 35332 5918 35334
rect 5942 35332 5998 35334
rect 6022 35332 6078 35334
rect 5782 34298 5838 34300
rect 5862 34298 5918 34300
rect 5942 34298 5998 34300
rect 6022 34298 6078 34300
rect 5782 34246 5828 34298
rect 5828 34246 5838 34298
rect 5862 34246 5892 34298
rect 5892 34246 5904 34298
rect 5904 34246 5918 34298
rect 5942 34246 5956 34298
rect 5956 34246 5968 34298
rect 5968 34246 5998 34298
rect 6022 34246 6032 34298
rect 6032 34246 6078 34298
rect 5782 34244 5838 34246
rect 5862 34244 5918 34246
rect 5942 34244 5998 34246
rect 6022 34244 6078 34246
rect 5782 33210 5838 33212
rect 5862 33210 5918 33212
rect 5942 33210 5998 33212
rect 6022 33210 6078 33212
rect 5782 33158 5828 33210
rect 5828 33158 5838 33210
rect 5862 33158 5892 33210
rect 5892 33158 5904 33210
rect 5904 33158 5918 33210
rect 5942 33158 5956 33210
rect 5956 33158 5968 33210
rect 5968 33158 5998 33210
rect 6022 33158 6032 33210
rect 6032 33158 6078 33210
rect 5782 33156 5838 33158
rect 5862 33156 5918 33158
rect 5942 33156 5998 33158
rect 6022 33156 6078 33158
rect 5782 32122 5838 32124
rect 5862 32122 5918 32124
rect 5942 32122 5998 32124
rect 6022 32122 6078 32124
rect 5782 32070 5828 32122
rect 5828 32070 5838 32122
rect 5862 32070 5892 32122
rect 5892 32070 5904 32122
rect 5904 32070 5918 32122
rect 5942 32070 5956 32122
rect 5956 32070 5968 32122
rect 5968 32070 5998 32122
rect 6022 32070 6032 32122
rect 6032 32070 6078 32122
rect 5782 32068 5838 32070
rect 5862 32068 5918 32070
rect 5942 32068 5998 32070
rect 6022 32068 6078 32070
rect 5782 31034 5838 31036
rect 5862 31034 5918 31036
rect 5942 31034 5998 31036
rect 6022 31034 6078 31036
rect 5782 30982 5828 31034
rect 5828 30982 5838 31034
rect 5862 30982 5892 31034
rect 5892 30982 5904 31034
rect 5904 30982 5918 31034
rect 5942 30982 5956 31034
rect 5956 30982 5968 31034
rect 5968 30982 5998 31034
rect 6022 30982 6032 31034
rect 6032 30982 6078 31034
rect 5782 30980 5838 30982
rect 5862 30980 5918 30982
rect 5942 30980 5998 30982
rect 6022 30980 6078 30982
rect 5446 30232 5502 30288
rect 5262 29144 5318 29200
rect 4986 28600 5042 28656
rect 4817 28314 4873 28316
rect 4897 28314 4953 28316
rect 4977 28314 5033 28316
rect 5057 28314 5113 28316
rect 4817 28262 4863 28314
rect 4863 28262 4873 28314
rect 4897 28262 4927 28314
rect 4927 28262 4939 28314
rect 4939 28262 4953 28314
rect 4977 28262 4991 28314
rect 4991 28262 5003 28314
rect 5003 28262 5033 28314
rect 5057 28262 5067 28314
rect 5067 28262 5113 28314
rect 4817 28260 4873 28262
rect 4897 28260 4953 28262
rect 4977 28260 5033 28262
rect 5057 28260 5113 28262
rect 4817 27226 4873 27228
rect 4897 27226 4953 27228
rect 4977 27226 5033 27228
rect 5057 27226 5113 27228
rect 4817 27174 4863 27226
rect 4863 27174 4873 27226
rect 4897 27174 4927 27226
rect 4927 27174 4939 27226
rect 4939 27174 4953 27226
rect 4977 27174 4991 27226
rect 4991 27174 5003 27226
rect 5003 27174 5033 27226
rect 5057 27174 5067 27226
rect 5067 27174 5113 27226
rect 4817 27172 4873 27174
rect 4897 27172 4953 27174
rect 4977 27172 5033 27174
rect 5057 27172 5113 27174
rect 5078 26832 5134 26888
rect 4817 26138 4873 26140
rect 4897 26138 4953 26140
rect 4977 26138 5033 26140
rect 5057 26138 5113 26140
rect 4817 26086 4863 26138
rect 4863 26086 4873 26138
rect 4897 26086 4927 26138
rect 4927 26086 4939 26138
rect 4939 26086 4953 26138
rect 4977 26086 4991 26138
rect 4991 26086 5003 26138
rect 5003 26086 5033 26138
rect 5057 26086 5067 26138
rect 5067 26086 5113 26138
rect 4817 26084 4873 26086
rect 4897 26084 4953 26086
rect 4977 26084 5033 26086
rect 5057 26084 5113 26086
rect 4817 25050 4873 25052
rect 4897 25050 4953 25052
rect 4977 25050 5033 25052
rect 5057 25050 5113 25052
rect 4817 24998 4863 25050
rect 4863 24998 4873 25050
rect 4897 24998 4927 25050
rect 4927 24998 4939 25050
rect 4939 24998 4953 25050
rect 4977 24998 4991 25050
rect 4991 24998 5003 25050
rect 5003 24998 5033 25050
rect 5057 24998 5067 25050
rect 5067 24998 5113 25050
rect 4817 24996 4873 24998
rect 4897 24996 4953 24998
rect 4977 24996 5033 24998
rect 5057 24996 5113 24998
rect 4817 23962 4873 23964
rect 4897 23962 4953 23964
rect 4977 23962 5033 23964
rect 5057 23962 5113 23964
rect 4817 23910 4863 23962
rect 4863 23910 4873 23962
rect 4897 23910 4927 23962
rect 4927 23910 4939 23962
rect 4939 23910 4953 23962
rect 4977 23910 4991 23962
rect 4991 23910 5003 23962
rect 5003 23910 5033 23962
rect 5057 23910 5067 23962
rect 5067 23910 5113 23962
rect 4817 23908 4873 23910
rect 4897 23908 4953 23910
rect 4977 23908 5033 23910
rect 5057 23908 5113 23910
rect 4817 22874 4873 22876
rect 4897 22874 4953 22876
rect 4977 22874 5033 22876
rect 5057 22874 5113 22876
rect 4817 22822 4863 22874
rect 4863 22822 4873 22874
rect 4897 22822 4927 22874
rect 4927 22822 4939 22874
rect 4939 22822 4953 22874
rect 4977 22822 4991 22874
rect 4991 22822 5003 22874
rect 5003 22822 5033 22874
rect 5057 22822 5067 22874
rect 5067 22822 5113 22874
rect 4817 22820 4873 22822
rect 4897 22820 4953 22822
rect 4977 22820 5033 22822
rect 5057 22820 5113 22822
rect 5262 22888 5318 22944
rect 5170 22480 5226 22536
rect 6182 30776 6238 30832
rect 5782 29946 5838 29948
rect 5862 29946 5918 29948
rect 5942 29946 5998 29948
rect 6022 29946 6078 29948
rect 5782 29894 5828 29946
rect 5828 29894 5838 29946
rect 5862 29894 5892 29946
rect 5892 29894 5904 29946
rect 5904 29894 5918 29946
rect 5942 29894 5956 29946
rect 5956 29894 5968 29946
rect 5968 29894 5998 29946
rect 6022 29894 6032 29946
rect 6032 29894 6078 29946
rect 5782 29892 5838 29894
rect 5862 29892 5918 29894
rect 5942 29892 5998 29894
rect 6022 29892 6078 29894
rect 6182 29688 6238 29744
rect 5782 28858 5838 28860
rect 5862 28858 5918 28860
rect 5942 28858 5998 28860
rect 6022 28858 6078 28860
rect 5782 28806 5828 28858
rect 5828 28806 5838 28858
rect 5862 28806 5892 28858
rect 5892 28806 5904 28858
rect 5904 28806 5918 28858
rect 5942 28806 5956 28858
rect 5956 28806 5968 28858
rect 5968 28806 5998 28858
rect 6022 28806 6032 28858
rect 6032 28806 6078 28858
rect 5782 28804 5838 28806
rect 5862 28804 5918 28806
rect 5942 28804 5998 28806
rect 6022 28804 6078 28806
rect 6090 27920 6146 27976
rect 5782 27770 5838 27772
rect 5862 27770 5918 27772
rect 5942 27770 5998 27772
rect 6022 27770 6078 27772
rect 5782 27718 5828 27770
rect 5828 27718 5838 27770
rect 5862 27718 5892 27770
rect 5892 27718 5904 27770
rect 5904 27718 5918 27770
rect 5942 27718 5956 27770
rect 5956 27718 5968 27770
rect 5968 27718 5998 27770
rect 6022 27718 6032 27770
rect 6032 27718 6078 27770
rect 5782 27716 5838 27718
rect 5862 27716 5918 27718
rect 5942 27716 5998 27718
rect 6022 27716 6078 27718
rect 5446 26324 5448 26344
rect 5448 26324 5500 26344
rect 5500 26324 5502 26344
rect 5446 26288 5502 26324
rect 5446 23976 5502 24032
rect 4817 21786 4873 21788
rect 4897 21786 4953 21788
rect 4977 21786 5033 21788
rect 5057 21786 5113 21788
rect 4817 21734 4863 21786
rect 4863 21734 4873 21786
rect 4897 21734 4927 21786
rect 4927 21734 4939 21786
rect 4939 21734 4953 21786
rect 4977 21734 4991 21786
rect 4991 21734 5003 21786
rect 5003 21734 5033 21786
rect 5057 21734 5067 21786
rect 5067 21734 5113 21786
rect 4817 21732 4873 21734
rect 4897 21732 4953 21734
rect 4977 21732 5033 21734
rect 5057 21732 5113 21734
rect 6182 27376 6238 27432
rect 5782 26682 5838 26684
rect 5862 26682 5918 26684
rect 5942 26682 5998 26684
rect 6022 26682 6078 26684
rect 5782 26630 5828 26682
rect 5828 26630 5838 26682
rect 5862 26630 5892 26682
rect 5892 26630 5904 26682
rect 5904 26630 5918 26682
rect 5942 26630 5956 26682
rect 5956 26630 5968 26682
rect 5968 26630 5998 26682
rect 6022 26630 6032 26682
rect 6032 26630 6078 26682
rect 5782 26628 5838 26630
rect 5862 26628 5918 26630
rect 5942 26628 5998 26630
rect 6022 26628 6078 26630
rect 5782 25594 5838 25596
rect 5862 25594 5918 25596
rect 5942 25594 5998 25596
rect 6022 25594 6078 25596
rect 5782 25542 5828 25594
rect 5828 25542 5838 25594
rect 5862 25542 5892 25594
rect 5892 25542 5904 25594
rect 5904 25542 5918 25594
rect 5942 25542 5956 25594
rect 5956 25542 5968 25594
rect 5968 25542 5998 25594
rect 6022 25542 6032 25594
rect 6032 25542 6078 25594
rect 5782 25540 5838 25542
rect 5862 25540 5918 25542
rect 5942 25540 5998 25542
rect 6022 25540 6078 25542
rect 6090 25236 6092 25256
rect 6092 25236 6144 25256
rect 6144 25236 6146 25256
rect 6090 25200 6146 25236
rect 6182 24520 6238 24576
rect 5782 24506 5838 24508
rect 5862 24506 5918 24508
rect 5942 24506 5998 24508
rect 6022 24506 6078 24508
rect 5782 24454 5828 24506
rect 5828 24454 5838 24506
rect 5862 24454 5892 24506
rect 5892 24454 5904 24506
rect 5904 24454 5918 24506
rect 5942 24454 5956 24506
rect 5956 24454 5968 24506
rect 5968 24454 5998 24506
rect 6022 24454 6032 24506
rect 6032 24454 6078 24506
rect 5782 24452 5838 24454
rect 5862 24452 5918 24454
rect 5942 24452 5998 24454
rect 6022 24452 6078 24454
rect 6182 23432 6238 23488
rect 5782 23418 5838 23420
rect 5862 23418 5918 23420
rect 5942 23418 5998 23420
rect 6022 23418 6078 23420
rect 5782 23366 5828 23418
rect 5828 23366 5838 23418
rect 5862 23366 5892 23418
rect 5892 23366 5904 23418
rect 5904 23366 5918 23418
rect 5942 23366 5956 23418
rect 5956 23366 5968 23418
rect 5968 23366 5998 23418
rect 6022 23366 6032 23418
rect 6032 23366 6078 23418
rect 5782 23364 5838 23366
rect 5862 23364 5918 23366
rect 5942 23364 5998 23366
rect 6022 23364 6078 23366
rect 5782 22330 5838 22332
rect 5862 22330 5918 22332
rect 5942 22330 5998 22332
rect 6022 22330 6078 22332
rect 5782 22278 5828 22330
rect 5828 22278 5838 22330
rect 5862 22278 5892 22330
rect 5892 22278 5904 22330
rect 5904 22278 5918 22330
rect 5942 22278 5956 22330
rect 5956 22278 5968 22330
rect 5968 22278 5998 22330
rect 6022 22278 6032 22330
rect 6032 22278 6078 22330
rect 5782 22276 5838 22278
rect 5862 22276 5918 22278
rect 5942 22276 5998 22278
rect 6022 22276 6078 22278
rect 4817 20698 4873 20700
rect 4897 20698 4953 20700
rect 4977 20698 5033 20700
rect 5057 20698 5113 20700
rect 4817 20646 4863 20698
rect 4863 20646 4873 20698
rect 4897 20646 4927 20698
rect 4927 20646 4939 20698
rect 4939 20646 4953 20698
rect 4977 20646 4991 20698
rect 4991 20646 5003 20698
rect 5003 20646 5033 20698
rect 5057 20646 5067 20698
rect 5067 20646 5113 20698
rect 4817 20644 4873 20646
rect 4897 20644 4953 20646
rect 4977 20644 5033 20646
rect 5057 20644 5113 20646
rect 4817 19610 4873 19612
rect 4897 19610 4953 19612
rect 4977 19610 5033 19612
rect 5057 19610 5113 19612
rect 4817 19558 4863 19610
rect 4863 19558 4873 19610
rect 4897 19558 4927 19610
rect 4927 19558 4939 19610
rect 4939 19558 4953 19610
rect 4977 19558 4991 19610
rect 4991 19558 5003 19610
rect 5003 19558 5033 19610
rect 5057 19558 5067 19610
rect 5067 19558 5113 19610
rect 4817 19556 4873 19558
rect 4897 19556 4953 19558
rect 4977 19556 5033 19558
rect 5057 19556 5113 19558
rect 4817 18522 4873 18524
rect 4897 18522 4953 18524
rect 4977 18522 5033 18524
rect 5057 18522 5113 18524
rect 4817 18470 4863 18522
rect 4863 18470 4873 18522
rect 4897 18470 4927 18522
rect 4927 18470 4939 18522
rect 4939 18470 4953 18522
rect 4977 18470 4991 18522
rect 4991 18470 5003 18522
rect 5003 18470 5033 18522
rect 5057 18470 5067 18522
rect 5067 18470 5113 18522
rect 4817 18468 4873 18470
rect 4897 18468 4953 18470
rect 4977 18468 5033 18470
rect 5057 18468 5113 18470
rect 2886 16346 2942 16348
rect 2966 16346 3022 16348
rect 3046 16346 3102 16348
rect 3126 16346 3182 16348
rect 2886 16294 2932 16346
rect 2932 16294 2942 16346
rect 2966 16294 2996 16346
rect 2996 16294 3008 16346
rect 3008 16294 3022 16346
rect 3046 16294 3060 16346
rect 3060 16294 3072 16346
rect 3072 16294 3102 16346
rect 3126 16294 3136 16346
rect 3136 16294 3182 16346
rect 2886 16292 2942 16294
rect 2966 16292 3022 16294
rect 3046 16292 3102 16294
rect 3126 16292 3182 16294
rect 1582 16224 1638 16280
rect 1921 15802 1977 15804
rect 2001 15802 2057 15804
rect 2081 15802 2137 15804
rect 2161 15802 2217 15804
rect 1921 15750 1967 15802
rect 1967 15750 1977 15802
rect 2001 15750 2031 15802
rect 2031 15750 2043 15802
rect 2043 15750 2057 15802
rect 2081 15750 2095 15802
rect 2095 15750 2107 15802
rect 2107 15750 2137 15802
rect 2161 15750 2171 15802
rect 2171 15750 2217 15802
rect 1921 15748 1977 15750
rect 2001 15748 2057 15750
rect 2081 15748 2137 15750
rect 2161 15748 2217 15750
rect 3852 15802 3908 15804
rect 3932 15802 3988 15804
rect 4012 15802 4068 15804
rect 4092 15802 4148 15804
rect 3852 15750 3898 15802
rect 3898 15750 3908 15802
rect 3932 15750 3962 15802
rect 3962 15750 3974 15802
rect 3974 15750 3988 15802
rect 4012 15750 4026 15802
rect 4026 15750 4038 15802
rect 4038 15750 4068 15802
rect 4092 15750 4102 15802
rect 4102 15750 4148 15802
rect 3852 15748 3908 15750
rect 3932 15748 3988 15750
rect 4012 15748 4068 15750
rect 4092 15748 4148 15750
rect 1582 15444 1584 15464
rect 1584 15444 1636 15464
rect 1636 15444 1638 15464
rect 1582 15408 1638 15444
rect 2886 15258 2942 15260
rect 2966 15258 3022 15260
rect 3046 15258 3102 15260
rect 3126 15258 3182 15260
rect 2886 15206 2932 15258
rect 2932 15206 2942 15258
rect 2966 15206 2996 15258
rect 2996 15206 3008 15258
rect 3008 15206 3022 15258
rect 3046 15206 3060 15258
rect 3060 15206 3072 15258
rect 3072 15206 3102 15258
rect 3126 15206 3136 15258
rect 3136 15206 3182 15258
rect 2886 15204 2942 15206
rect 2966 15204 3022 15206
rect 3046 15204 3102 15206
rect 3126 15204 3182 15206
rect 1582 14728 1638 14784
rect 1921 14714 1977 14716
rect 2001 14714 2057 14716
rect 2081 14714 2137 14716
rect 2161 14714 2217 14716
rect 1921 14662 1967 14714
rect 1967 14662 1977 14714
rect 2001 14662 2031 14714
rect 2031 14662 2043 14714
rect 2043 14662 2057 14714
rect 2081 14662 2095 14714
rect 2095 14662 2107 14714
rect 2107 14662 2137 14714
rect 2161 14662 2171 14714
rect 2171 14662 2217 14714
rect 1921 14660 1977 14662
rect 2001 14660 2057 14662
rect 2081 14660 2137 14662
rect 2161 14660 2217 14662
rect 3852 14714 3908 14716
rect 3932 14714 3988 14716
rect 4012 14714 4068 14716
rect 4092 14714 4148 14716
rect 3852 14662 3898 14714
rect 3898 14662 3908 14714
rect 3932 14662 3962 14714
rect 3962 14662 3974 14714
rect 3974 14662 3988 14714
rect 4012 14662 4026 14714
rect 4026 14662 4038 14714
rect 4038 14662 4068 14714
rect 4092 14662 4102 14714
rect 4102 14662 4148 14714
rect 3852 14660 3908 14662
rect 3932 14660 3988 14662
rect 4012 14660 4068 14662
rect 4092 14660 4148 14662
rect 4817 17434 4873 17436
rect 4897 17434 4953 17436
rect 4977 17434 5033 17436
rect 5057 17434 5113 17436
rect 4817 17382 4863 17434
rect 4863 17382 4873 17434
rect 4897 17382 4927 17434
rect 4927 17382 4939 17434
rect 4939 17382 4953 17434
rect 4977 17382 4991 17434
rect 4991 17382 5003 17434
rect 5003 17382 5033 17434
rect 5057 17382 5067 17434
rect 5067 17382 5113 17434
rect 4817 17380 4873 17382
rect 4897 17380 4953 17382
rect 4977 17380 5033 17382
rect 5057 17380 5113 17382
rect 4817 16346 4873 16348
rect 4897 16346 4953 16348
rect 4977 16346 5033 16348
rect 5057 16346 5113 16348
rect 4817 16294 4863 16346
rect 4863 16294 4873 16346
rect 4897 16294 4927 16346
rect 4927 16294 4939 16346
rect 4939 16294 4953 16346
rect 4977 16294 4991 16346
rect 4991 16294 5003 16346
rect 5003 16294 5033 16346
rect 5057 16294 5067 16346
rect 5067 16294 5113 16346
rect 4817 16292 4873 16294
rect 4897 16292 4953 16294
rect 4977 16292 5033 16294
rect 5057 16292 5113 16294
rect 4817 15258 4873 15260
rect 4897 15258 4953 15260
rect 4977 15258 5033 15260
rect 5057 15258 5113 15260
rect 4817 15206 4863 15258
rect 4863 15206 4873 15258
rect 4897 15206 4927 15258
rect 4927 15206 4939 15258
rect 4939 15206 4953 15258
rect 4977 15206 4991 15258
rect 4991 15206 5003 15258
rect 5003 15206 5033 15258
rect 5057 15206 5067 15258
rect 5067 15206 5113 15258
rect 4817 15204 4873 15206
rect 4897 15204 4953 15206
rect 4977 15204 5033 15206
rect 5057 15204 5113 15206
rect 2886 14170 2942 14172
rect 2966 14170 3022 14172
rect 3046 14170 3102 14172
rect 3126 14170 3182 14172
rect 2886 14118 2932 14170
rect 2932 14118 2942 14170
rect 2966 14118 2996 14170
rect 2996 14118 3008 14170
rect 3008 14118 3022 14170
rect 3046 14118 3060 14170
rect 3060 14118 3072 14170
rect 3072 14118 3102 14170
rect 3126 14118 3136 14170
rect 3136 14118 3182 14170
rect 2886 14116 2942 14118
rect 2966 14116 3022 14118
rect 3046 14116 3102 14118
rect 3126 14116 3182 14118
rect 4817 14170 4873 14172
rect 4897 14170 4953 14172
rect 4977 14170 5033 14172
rect 5057 14170 5113 14172
rect 4817 14118 4863 14170
rect 4863 14118 4873 14170
rect 4897 14118 4927 14170
rect 4927 14118 4939 14170
rect 4939 14118 4953 14170
rect 4977 14118 4991 14170
rect 4991 14118 5003 14170
rect 5003 14118 5033 14170
rect 5057 14118 5067 14170
rect 5067 14118 5113 14170
rect 4817 14116 4873 14118
rect 4897 14116 4953 14118
rect 4977 14116 5033 14118
rect 5057 14116 5113 14118
rect 1582 13912 1638 13968
rect 1921 13626 1977 13628
rect 2001 13626 2057 13628
rect 2081 13626 2137 13628
rect 2161 13626 2217 13628
rect 1921 13574 1967 13626
rect 1967 13574 1977 13626
rect 2001 13574 2031 13626
rect 2031 13574 2043 13626
rect 2043 13574 2057 13626
rect 2081 13574 2095 13626
rect 2095 13574 2107 13626
rect 2107 13574 2137 13626
rect 2161 13574 2171 13626
rect 2171 13574 2217 13626
rect 1921 13572 1977 13574
rect 2001 13572 2057 13574
rect 2081 13572 2137 13574
rect 2161 13572 2217 13574
rect 3852 13626 3908 13628
rect 3932 13626 3988 13628
rect 4012 13626 4068 13628
rect 4092 13626 4148 13628
rect 3852 13574 3898 13626
rect 3898 13574 3908 13626
rect 3932 13574 3962 13626
rect 3962 13574 3974 13626
rect 3974 13574 3988 13626
rect 4012 13574 4026 13626
rect 4026 13574 4038 13626
rect 4038 13574 4068 13626
rect 4092 13574 4102 13626
rect 4102 13574 4148 13626
rect 3852 13572 3908 13574
rect 3932 13572 3988 13574
rect 4012 13572 4068 13574
rect 4092 13572 4148 13574
rect 1582 13096 1638 13152
rect 2886 13082 2942 13084
rect 2966 13082 3022 13084
rect 3046 13082 3102 13084
rect 3126 13082 3182 13084
rect 2886 13030 2932 13082
rect 2932 13030 2942 13082
rect 2966 13030 2996 13082
rect 2996 13030 3008 13082
rect 3008 13030 3022 13082
rect 3046 13030 3060 13082
rect 3060 13030 3072 13082
rect 3072 13030 3102 13082
rect 3126 13030 3136 13082
rect 3136 13030 3182 13082
rect 2886 13028 2942 13030
rect 2966 13028 3022 13030
rect 3046 13028 3102 13030
rect 3126 13028 3182 13030
rect 4817 13082 4873 13084
rect 4897 13082 4953 13084
rect 4977 13082 5033 13084
rect 5057 13082 5113 13084
rect 4817 13030 4863 13082
rect 4863 13030 4873 13082
rect 4897 13030 4927 13082
rect 4927 13030 4939 13082
rect 4939 13030 4953 13082
rect 4977 13030 4991 13082
rect 4991 13030 5003 13082
rect 5003 13030 5033 13082
rect 5057 13030 5067 13082
rect 5067 13030 5113 13082
rect 4817 13028 4873 13030
rect 4897 13028 4953 13030
rect 4977 13028 5033 13030
rect 5057 13028 5113 13030
rect 6182 21800 6238 21856
rect 5782 21242 5838 21244
rect 5862 21242 5918 21244
rect 5942 21242 5998 21244
rect 6022 21242 6078 21244
rect 5782 21190 5828 21242
rect 5828 21190 5838 21242
rect 5862 21190 5892 21242
rect 5892 21190 5904 21242
rect 5904 21190 5918 21242
rect 5942 21190 5956 21242
rect 5956 21190 5968 21242
rect 5968 21190 5998 21242
rect 6022 21190 6032 21242
rect 6032 21190 6078 21242
rect 5782 21188 5838 21190
rect 5862 21188 5918 21190
rect 5942 21188 5998 21190
rect 6022 21188 6078 21190
rect 6182 21120 6238 21176
rect 6090 20576 6146 20632
rect 5782 20154 5838 20156
rect 5862 20154 5918 20156
rect 5942 20154 5998 20156
rect 6022 20154 6078 20156
rect 5782 20102 5828 20154
rect 5828 20102 5838 20154
rect 5862 20102 5892 20154
rect 5892 20102 5904 20154
rect 5904 20102 5918 20154
rect 5942 20102 5956 20154
rect 5956 20102 5968 20154
rect 5968 20102 5998 20154
rect 6022 20102 6032 20154
rect 6032 20102 6078 20154
rect 5782 20100 5838 20102
rect 5862 20100 5918 20102
rect 5942 20100 5998 20102
rect 6022 20100 6078 20102
rect 6182 20032 6238 20088
rect 6090 19488 6146 19544
rect 5782 19066 5838 19068
rect 5862 19066 5918 19068
rect 5942 19066 5998 19068
rect 6022 19066 6078 19068
rect 5782 19014 5828 19066
rect 5828 19014 5838 19066
rect 5862 19014 5892 19066
rect 5892 19014 5904 19066
rect 5904 19014 5918 19066
rect 5942 19014 5956 19066
rect 5956 19014 5968 19066
rect 5968 19014 5998 19066
rect 6022 19014 6032 19066
rect 6032 19014 6078 19066
rect 5782 19012 5838 19014
rect 5862 19012 5918 19014
rect 5942 19012 5998 19014
rect 6022 19012 6078 19014
rect 6458 18944 6514 19000
rect 6090 18400 6146 18456
rect 5446 17176 5502 17232
rect 5782 17978 5838 17980
rect 5862 17978 5918 17980
rect 5942 17978 5998 17980
rect 6022 17978 6078 17980
rect 5782 17926 5828 17978
rect 5828 17926 5838 17978
rect 5862 17926 5892 17978
rect 5892 17926 5904 17978
rect 5904 17926 5918 17978
rect 5942 17926 5956 17978
rect 5956 17926 5968 17978
rect 5968 17926 5998 17978
rect 6022 17926 6032 17978
rect 6032 17926 6078 17978
rect 5782 17924 5838 17926
rect 5862 17924 5918 17926
rect 5942 17924 5998 17926
rect 6022 17924 6078 17926
rect 6182 17720 6238 17776
rect 5782 16890 5838 16892
rect 5862 16890 5918 16892
rect 5942 16890 5998 16892
rect 6022 16890 6078 16892
rect 5782 16838 5828 16890
rect 5828 16838 5838 16890
rect 5862 16838 5892 16890
rect 5892 16838 5904 16890
rect 5904 16838 5918 16890
rect 5942 16838 5956 16890
rect 5956 16838 5968 16890
rect 5968 16838 5998 16890
rect 6022 16838 6032 16890
rect 6032 16838 6078 16890
rect 5782 16836 5838 16838
rect 5862 16836 5918 16838
rect 5942 16836 5998 16838
rect 6022 16836 6078 16838
rect 6182 16632 6238 16688
rect 5446 15000 5502 15056
rect 5782 15802 5838 15804
rect 5862 15802 5918 15804
rect 5942 15802 5998 15804
rect 6022 15802 6078 15804
rect 5782 15750 5828 15802
rect 5828 15750 5838 15802
rect 5862 15750 5892 15802
rect 5892 15750 5904 15802
rect 5904 15750 5918 15802
rect 5942 15750 5956 15802
rect 5956 15750 5968 15802
rect 5968 15750 5998 15802
rect 6022 15750 6032 15802
rect 6032 15750 6078 15802
rect 5782 15748 5838 15750
rect 5862 15748 5918 15750
rect 5942 15748 5998 15750
rect 6022 15748 6078 15750
rect 6182 15544 6238 15600
rect 5782 14714 5838 14716
rect 5862 14714 5918 14716
rect 5942 14714 5998 14716
rect 6022 14714 6078 14716
rect 5782 14662 5828 14714
rect 5828 14662 5838 14714
rect 5862 14662 5892 14714
rect 5892 14662 5904 14714
rect 5904 14662 5918 14714
rect 5942 14662 5956 14714
rect 5956 14662 5968 14714
rect 5968 14662 5998 14714
rect 6022 14662 6032 14714
rect 6032 14662 6078 14714
rect 5782 14660 5838 14662
rect 5862 14660 5918 14662
rect 5942 14660 5998 14662
rect 6022 14660 6078 14662
rect 6366 16088 6422 16144
rect 6182 14456 6238 14512
rect 1921 12538 1977 12540
rect 2001 12538 2057 12540
rect 2081 12538 2137 12540
rect 2161 12538 2217 12540
rect 1921 12486 1967 12538
rect 1967 12486 1977 12538
rect 2001 12486 2031 12538
rect 2031 12486 2043 12538
rect 2043 12486 2057 12538
rect 2081 12486 2095 12538
rect 2095 12486 2107 12538
rect 2107 12486 2137 12538
rect 2161 12486 2171 12538
rect 2171 12486 2217 12538
rect 1921 12484 1977 12486
rect 2001 12484 2057 12486
rect 2081 12484 2137 12486
rect 2161 12484 2217 12486
rect 1582 12416 1638 12472
rect 3852 12538 3908 12540
rect 3932 12538 3988 12540
rect 4012 12538 4068 12540
rect 4092 12538 4148 12540
rect 3852 12486 3898 12538
rect 3898 12486 3908 12538
rect 3932 12486 3962 12538
rect 3962 12486 3974 12538
rect 3974 12486 3988 12538
rect 4012 12486 4026 12538
rect 4026 12486 4038 12538
rect 4038 12486 4068 12538
rect 4092 12486 4102 12538
rect 4102 12486 4148 12538
rect 3852 12484 3908 12486
rect 3932 12484 3988 12486
rect 4012 12484 4068 12486
rect 4092 12484 4148 12486
rect 2886 11994 2942 11996
rect 2966 11994 3022 11996
rect 3046 11994 3102 11996
rect 3126 11994 3182 11996
rect 2886 11942 2932 11994
rect 2932 11942 2942 11994
rect 2966 11942 2996 11994
rect 2996 11942 3008 11994
rect 3008 11942 3022 11994
rect 3046 11942 3060 11994
rect 3060 11942 3072 11994
rect 3072 11942 3102 11994
rect 3126 11942 3136 11994
rect 3136 11942 3182 11994
rect 2886 11940 2942 11942
rect 2966 11940 3022 11942
rect 3046 11940 3102 11942
rect 3126 11940 3182 11942
rect 4817 11994 4873 11996
rect 4897 11994 4953 11996
rect 4977 11994 5033 11996
rect 5057 11994 5113 11996
rect 4817 11942 4863 11994
rect 4863 11942 4873 11994
rect 4897 11942 4927 11994
rect 4927 11942 4939 11994
rect 4939 11942 4953 11994
rect 4977 11942 4991 11994
rect 4991 11942 5003 11994
rect 5003 11942 5033 11994
rect 5057 11942 5067 11994
rect 5067 11942 5113 11994
rect 4817 11940 4873 11942
rect 4897 11940 4953 11942
rect 4977 11940 5033 11942
rect 5057 11940 5113 11942
rect 5814 13776 5870 13832
rect 5782 13626 5838 13628
rect 5862 13626 5918 13628
rect 5942 13626 5998 13628
rect 6022 13626 6078 13628
rect 5782 13574 5828 13626
rect 5828 13574 5838 13626
rect 5862 13574 5892 13626
rect 5892 13574 5904 13626
rect 5904 13574 5918 13626
rect 5942 13574 5956 13626
rect 5956 13574 5968 13626
rect 5968 13574 5998 13626
rect 6022 13574 6032 13626
rect 6032 13574 6078 13626
rect 5782 13572 5838 13574
rect 5862 13572 5918 13574
rect 5942 13572 5998 13574
rect 6022 13572 6078 13574
rect 6826 31320 6882 31376
rect 6826 25744 6882 25800
rect 6090 13268 6092 13288
rect 6092 13268 6144 13288
rect 6144 13268 6146 13288
rect 6090 13232 6146 13268
rect 5814 12688 5870 12744
rect 5782 12538 5838 12540
rect 5862 12538 5918 12540
rect 5942 12538 5998 12540
rect 6022 12538 6078 12540
rect 5782 12486 5828 12538
rect 5828 12486 5838 12538
rect 5862 12486 5892 12538
rect 5892 12486 5904 12538
rect 5904 12486 5918 12538
rect 5942 12486 5956 12538
rect 5956 12486 5968 12538
rect 5968 12486 5998 12538
rect 6022 12486 6032 12538
rect 6032 12486 6078 12538
rect 5782 12484 5838 12486
rect 5862 12484 5918 12486
rect 5942 12484 5998 12486
rect 6022 12484 6078 12486
rect 6090 12180 6092 12200
rect 6092 12180 6144 12200
rect 6144 12180 6146 12200
rect 6090 12144 6146 12180
rect 1582 11600 1638 11656
rect 1921 11450 1977 11452
rect 2001 11450 2057 11452
rect 2081 11450 2137 11452
rect 2161 11450 2217 11452
rect 1921 11398 1967 11450
rect 1967 11398 1977 11450
rect 2001 11398 2031 11450
rect 2031 11398 2043 11450
rect 2043 11398 2057 11450
rect 2081 11398 2095 11450
rect 2095 11398 2107 11450
rect 2107 11398 2137 11450
rect 2161 11398 2171 11450
rect 2171 11398 2217 11450
rect 1921 11396 1977 11398
rect 2001 11396 2057 11398
rect 2081 11396 2137 11398
rect 2161 11396 2217 11398
rect 3852 11450 3908 11452
rect 3932 11450 3988 11452
rect 4012 11450 4068 11452
rect 4092 11450 4148 11452
rect 3852 11398 3898 11450
rect 3898 11398 3908 11450
rect 3932 11398 3962 11450
rect 3962 11398 3974 11450
rect 3974 11398 3988 11450
rect 4012 11398 4026 11450
rect 4026 11398 4038 11450
rect 4038 11398 4068 11450
rect 4092 11398 4102 11450
rect 4102 11398 4148 11450
rect 3852 11396 3908 11398
rect 3932 11396 3988 11398
rect 4012 11396 4068 11398
rect 4092 11396 4148 11398
rect 6182 11600 6238 11656
rect 5782 11450 5838 11452
rect 5862 11450 5918 11452
rect 5942 11450 5998 11452
rect 6022 11450 6078 11452
rect 5782 11398 5828 11450
rect 5828 11398 5838 11450
rect 5862 11398 5892 11450
rect 5892 11398 5904 11450
rect 5904 11398 5918 11450
rect 5942 11398 5956 11450
rect 5956 11398 5968 11450
rect 5968 11398 5998 11450
rect 6022 11398 6032 11450
rect 6032 11398 6078 11450
rect 5782 11396 5838 11398
rect 5862 11396 5918 11398
rect 5942 11396 5998 11398
rect 6022 11396 6078 11398
rect 4802 11092 4804 11112
rect 4804 11092 4856 11112
rect 4856 11092 4858 11112
rect 1582 10956 1584 10976
rect 1584 10956 1636 10976
rect 1636 10956 1638 10976
rect 1582 10920 1638 10956
rect 2886 10906 2942 10908
rect 2966 10906 3022 10908
rect 3046 10906 3102 10908
rect 3126 10906 3182 10908
rect 2886 10854 2932 10906
rect 2932 10854 2942 10906
rect 2966 10854 2996 10906
rect 2996 10854 3008 10906
rect 3008 10854 3022 10906
rect 3046 10854 3060 10906
rect 3060 10854 3072 10906
rect 3072 10854 3102 10906
rect 3126 10854 3136 10906
rect 3136 10854 3182 10906
rect 2886 10852 2942 10854
rect 2966 10852 3022 10854
rect 3046 10852 3102 10854
rect 3126 10852 3182 10854
rect 4802 11056 4858 11092
rect 4817 10906 4873 10908
rect 4897 10906 4953 10908
rect 4977 10906 5033 10908
rect 5057 10906 5113 10908
rect 4817 10854 4863 10906
rect 4863 10854 4873 10906
rect 4897 10854 4927 10906
rect 4927 10854 4939 10906
rect 4939 10854 4953 10906
rect 4977 10854 4991 10906
rect 4991 10854 5003 10906
rect 5003 10854 5033 10906
rect 5057 10854 5067 10906
rect 5067 10854 5113 10906
rect 4817 10852 4873 10854
rect 4897 10852 4953 10854
rect 4977 10852 5033 10854
rect 5057 10852 5113 10854
rect 5354 10512 5410 10568
rect 1921 10362 1977 10364
rect 2001 10362 2057 10364
rect 2081 10362 2137 10364
rect 2161 10362 2217 10364
rect 1921 10310 1967 10362
rect 1967 10310 1977 10362
rect 2001 10310 2031 10362
rect 2031 10310 2043 10362
rect 2043 10310 2057 10362
rect 2081 10310 2095 10362
rect 2095 10310 2107 10362
rect 2107 10310 2137 10362
rect 2161 10310 2171 10362
rect 2171 10310 2217 10362
rect 1921 10308 1977 10310
rect 2001 10308 2057 10310
rect 2081 10308 2137 10310
rect 2161 10308 2217 10310
rect 3852 10362 3908 10364
rect 3932 10362 3988 10364
rect 4012 10362 4068 10364
rect 4092 10362 4148 10364
rect 3852 10310 3898 10362
rect 3898 10310 3908 10362
rect 3932 10310 3962 10362
rect 3962 10310 3974 10362
rect 3974 10310 3988 10362
rect 4012 10310 4026 10362
rect 4026 10310 4038 10362
rect 4038 10310 4068 10362
rect 4092 10310 4102 10362
rect 4102 10310 4148 10362
rect 3852 10308 3908 10310
rect 3932 10308 3988 10310
rect 4012 10308 4068 10310
rect 4092 10308 4148 10310
rect 1582 10104 1638 10160
rect 2886 9818 2942 9820
rect 2966 9818 3022 9820
rect 3046 9818 3102 9820
rect 3126 9818 3182 9820
rect 2886 9766 2932 9818
rect 2932 9766 2942 9818
rect 2966 9766 2996 9818
rect 2996 9766 3008 9818
rect 3008 9766 3022 9818
rect 3046 9766 3060 9818
rect 3060 9766 3072 9818
rect 3072 9766 3102 9818
rect 3126 9766 3136 9818
rect 3136 9766 3182 9818
rect 2886 9764 2942 9766
rect 2966 9764 3022 9766
rect 3046 9764 3102 9766
rect 3126 9764 3182 9766
rect 4817 9818 4873 9820
rect 4897 9818 4953 9820
rect 4977 9818 5033 9820
rect 5057 9818 5113 9820
rect 4817 9766 4863 9818
rect 4863 9766 4873 9818
rect 4897 9766 4927 9818
rect 4927 9766 4939 9818
rect 4939 9766 4953 9818
rect 4977 9766 4991 9818
rect 4991 9766 5003 9818
rect 5003 9766 5033 9818
rect 5057 9766 5067 9818
rect 5067 9766 5113 9818
rect 4817 9764 4873 9766
rect 4897 9764 4953 9766
rect 4977 9764 5033 9766
rect 5057 9764 5113 9766
rect 5782 10362 5838 10364
rect 5862 10362 5918 10364
rect 5942 10362 5998 10364
rect 6022 10362 6078 10364
rect 5782 10310 5828 10362
rect 5828 10310 5838 10362
rect 5862 10310 5892 10362
rect 5892 10310 5904 10362
rect 5904 10310 5918 10362
rect 5942 10310 5956 10362
rect 5956 10310 5968 10362
rect 5968 10310 5998 10362
rect 6022 10310 6032 10362
rect 6032 10310 6078 10362
rect 5782 10308 5838 10310
rect 5862 10308 5918 10310
rect 5942 10308 5998 10310
rect 6022 10308 6078 10310
rect 5446 9832 5502 9888
rect 5170 9424 5226 9480
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 1921 9274 1977 9276
rect 2001 9274 2057 9276
rect 2081 9274 2137 9276
rect 2161 9274 2217 9276
rect 1921 9222 1967 9274
rect 1967 9222 1977 9274
rect 2001 9222 2031 9274
rect 2031 9222 2043 9274
rect 2043 9222 2057 9274
rect 2081 9222 2095 9274
rect 2095 9222 2107 9274
rect 2107 9222 2137 9274
rect 2161 9222 2171 9274
rect 2171 9222 2217 9274
rect 1921 9220 1977 9222
rect 2001 9220 2057 9222
rect 2081 9220 2137 9222
rect 2161 9220 2217 9222
rect 3852 9274 3908 9276
rect 3932 9274 3988 9276
rect 4012 9274 4068 9276
rect 4092 9274 4148 9276
rect 3852 9222 3898 9274
rect 3898 9222 3908 9274
rect 3932 9222 3962 9274
rect 3962 9222 3974 9274
rect 3974 9222 3988 9274
rect 4012 9222 4026 9274
rect 4026 9222 4038 9274
rect 4038 9222 4068 9274
rect 4092 9222 4102 9274
rect 4102 9222 4148 9274
rect 3852 9220 3908 9222
rect 3932 9220 3988 9222
rect 4012 9220 4068 9222
rect 4092 9220 4148 9222
rect 2886 8730 2942 8732
rect 2966 8730 3022 8732
rect 3046 8730 3102 8732
rect 3126 8730 3182 8732
rect 2886 8678 2932 8730
rect 2932 8678 2942 8730
rect 2966 8678 2996 8730
rect 2996 8678 3008 8730
rect 3008 8678 3022 8730
rect 3046 8678 3060 8730
rect 3060 8678 3072 8730
rect 3072 8678 3102 8730
rect 3126 8678 3136 8730
rect 3136 8678 3182 8730
rect 2886 8676 2942 8678
rect 2966 8676 3022 8678
rect 3046 8676 3102 8678
rect 3126 8676 3182 8678
rect 1582 8608 1638 8664
rect 1921 8186 1977 8188
rect 2001 8186 2057 8188
rect 2081 8186 2137 8188
rect 2161 8186 2217 8188
rect 1921 8134 1967 8186
rect 1967 8134 1977 8186
rect 2001 8134 2031 8186
rect 2031 8134 2043 8186
rect 2043 8134 2057 8186
rect 2081 8134 2095 8186
rect 2095 8134 2107 8186
rect 2107 8134 2137 8186
rect 2161 8134 2171 8186
rect 2171 8134 2217 8186
rect 1921 8132 1977 8134
rect 2001 8132 2057 8134
rect 2081 8132 2137 8134
rect 2161 8132 2217 8134
rect 3852 8186 3908 8188
rect 3932 8186 3988 8188
rect 4012 8186 4068 8188
rect 4092 8186 4148 8188
rect 3852 8134 3898 8186
rect 3898 8134 3908 8186
rect 3932 8134 3962 8186
rect 3962 8134 3974 8186
rect 3974 8134 3988 8186
rect 4012 8134 4026 8186
rect 4026 8134 4038 8186
rect 4038 8134 4068 8186
rect 4092 8134 4102 8186
rect 4102 8134 4148 8186
rect 3852 8132 3908 8134
rect 3932 8132 3988 8134
rect 4012 8132 4068 8134
rect 4092 8132 4148 8134
rect 1582 7792 1638 7848
rect 2886 7642 2942 7644
rect 2966 7642 3022 7644
rect 3046 7642 3102 7644
rect 3126 7642 3182 7644
rect 2886 7590 2932 7642
rect 2932 7590 2942 7642
rect 2966 7590 2996 7642
rect 2996 7590 3008 7642
rect 3008 7590 3022 7642
rect 3046 7590 3060 7642
rect 3060 7590 3072 7642
rect 3072 7590 3102 7642
rect 3126 7590 3136 7642
rect 3136 7590 3182 7642
rect 2886 7588 2942 7590
rect 2966 7588 3022 7590
rect 3046 7588 3102 7590
rect 3126 7588 3182 7590
rect 1582 7148 1584 7168
rect 1584 7148 1636 7168
rect 1636 7148 1638 7168
rect 1582 7112 1638 7148
rect 1921 7098 1977 7100
rect 2001 7098 2057 7100
rect 2081 7098 2137 7100
rect 2161 7098 2217 7100
rect 1921 7046 1967 7098
rect 1967 7046 1977 7098
rect 2001 7046 2031 7098
rect 2031 7046 2043 7098
rect 2043 7046 2057 7098
rect 2081 7046 2095 7098
rect 2095 7046 2107 7098
rect 2107 7046 2137 7098
rect 2161 7046 2171 7098
rect 2171 7046 2217 7098
rect 1921 7044 1977 7046
rect 2001 7044 2057 7046
rect 2081 7044 2137 7046
rect 2161 7044 2217 7046
rect 2886 6554 2942 6556
rect 2966 6554 3022 6556
rect 3046 6554 3102 6556
rect 3126 6554 3182 6556
rect 2886 6502 2932 6554
rect 2932 6502 2942 6554
rect 2966 6502 2996 6554
rect 2996 6502 3008 6554
rect 3008 6502 3022 6554
rect 3046 6502 3060 6554
rect 3060 6502 3072 6554
rect 3072 6502 3102 6554
rect 3126 6502 3136 6554
rect 3136 6502 3182 6554
rect 2886 6500 2942 6502
rect 2966 6500 3022 6502
rect 3046 6500 3102 6502
rect 3126 6500 3182 6502
rect 1582 6296 1638 6352
rect 3852 7098 3908 7100
rect 3932 7098 3988 7100
rect 4012 7098 4068 7100
rect 4092 7098 4148 7100
rect 3852 7046 3898 7098
rect 3898 7046 3908 7098
rect 3932 7046 3962 7098
rect 3962 7046 3974 7098
rect 3974 7046 3988 7098
rect 4012 7046 4026 7098
rect 4026 7046 4038 7098
rect 4038 7046 4068 7098
rect 4092 7046 4102 7098
rect 4102 7046 4148 7098
rect 3852 7044 3908 7046
rect 3932 7044 3988 7046
rect 4012 7044 4068 7046
rect 4092 7044 4148 7046
rect 4817 8730 4873 8732
rect 4897 8730 4953 8732
rect 4977 8730 5033 8732
rect 5057 8730 5113 8732
rect 4817 8678 4863 8730
rect 4863 8678 4873 8730
rect 4897 8678 4927 8730
rect 4927 8678 4939 8730
rect 4939 8678 4953 8730
rect 4977 8678 4991 8730
rect 4991 8678 5003 8730
rect 5003 8678 5033 8730
rect 5057 8678 5067 8730
rect 5067 8678 5113 8730
rect 4817 8676 4873 8678
rect 4897 8676 4953 8678
rect 4977 8676 5033 8678
rect 5057 8676 5113 8678
rect 4817 7642 4873 7644
rect 4897 7642 4953 7644
rect 4977 7642 5033 7644
rect 5057 7642 5113 7644
rect 4817 7590 4863 7642
rect 4863 7590 4873 7642
rect 4897 7590 4927 7642
rect 4927 7590 4939 7642
rect 4939 7590 4953 7642
rect 4977 7590 4991 7642
rect 4991 7590 5003 7642
rect 5003 7590 5033 7642
rect 5057 7590 5067 7642
rect 5067 7590 5113 7642
rect 4817 7588 4873 7590
rect 4897 7588 4953 7590
rect 4977 7588 5033 7590
rect 5057 7588 5113 7590
rect 5782 9274 5838 9276
rect 5862 9274 5918 9276
rect 5942 9274 5998 9276
rect 6022 9274 6078 9276
rect 5782 9222 5828 9274
rect 5828 9222 5838 9274
rect 5862 9222 5892 9274
rect 5892 9222 5904 9274
rect 5904 9222 5918 9274
rect 5942 9222 5956 9274
rect 5956 9222 5968 9274
rect 5968 9222 5998 9274
rect 6022 9222 6032 9274
rect 6032 9222 6078 9274
rect 5782 9220 5838 9222
rect 5862 9220 5918 9222
rect 5942 9220 5998 9222
rect 6022 9220 6078 9222
rect 6918 8780 6920 8800
rect 6920 8780 6972 8800
rect 6972 8780 6974 8800
rect 5446 8336 5502 8392
rect 5782 8186 5838 8188
rect 5862 8186 5918 8188
rect 5942 8186 5998 8188
rect 6022 8186 6078 8188
rect 5782 8134 5828 8186
rect 5828 8134 5838 8186
rect 5862 8134 5892 8186
rect 5892 8134 5904 8186
rect 5904 8134 5918 8186
rect 5942 8134 5956 8186
rect 5956 8134 5968 8186
rect 5968 8134 5998 8186
rect 6022 8134 6032 8186
rect 6032 8134 6078 8186
rect 5782 8132 5838 8134
rect 5862 8132 5918 8134
rect 5942 8132 5998 8134
rect 6022 8132 6078 8134
rect 5354 7656 5410 7712
rect 1921 6010 1977 6012
rect 2001 6010 2057 6012
rect 2081 6010 2137 6012
rect 2161 6010 2217 6012
rect 1921 5958 1967 6010
rect 1967 5958 1977 6010
rect 2001 5958 2031 6010
rect 2031 5958 2043 6010
rect 2043 5958 2057 6010
rect 2081 5958 2095 6010
rect 2095 5958 2107 6010
rect 2107 5958 2137 6010
rect 2161 5958 2171 6010
rect 2171 5958 2217 6010
rect 1921 5956 1977 5958
rect 2001 5956 2057 5958
rect 2081 5956 2137 5958
rect 2161 5956 2217 5958
rect 3852 6010 3908 6012
rect 3932 6010 3988 6012
rect 4012 6010 4068 6012
rect 4092 6010 4148 6012
rect 3852 5958 3898 6010
rect 3898 5958 3908 6010
rect 3932 5958 3962 6010
rect 3962 5958 3974 6010
rect 3974 5958 3988 6010
rect 4012 5958 4026 6010
rect 4026 5958 4038 6010
rect 4038 5958 4068 6010
rect 4092 5958 4102 6010
rect 4102 5958 4148 6010
rect 3852 5956 3908 5958
rect 3932 5956 3988 5958
rect 4012 5956 4068 5958
rect 4092 5956 4148 5958
rect 1582 5616 1638 5672
rect 2886 5466 2942 5468
rect 2966 5466 3022 5468
rect 3046 5466 3102 5468
rect 3126 5466 3182 5468
rect 2886 5414 2932 5466
rect 2932 5414 2942 5466
rect 2966 5414 2996 5466
rect 2996 5414 3008 5466
rect 3008 5414 3022 5466
rect 3046 5414 3060 5466
rect 3060 5414 3072 5466
rect 3072 5414 3102 5466
rect 3126 5414 3136 5466
rect 3136 5414 3182 5466
rect 2886 5412 2942 5414
rect 2966 5412 3022 5414
rect 3046 5412 3102 5414
rect 3126 5412 3182 5414
rect 3606 5228 3662 5264
rect 3606 5208 3608 5228
rect 3608 5208 3660 5228
rect 3660 5208 3662 5228
rect 1921 4922 1977 4924
rect 2001 4922 2057 4924
rect 2081 4922 2137 4924
rect 2161 4922 2217 4924
rect 1921 4870 1967 4922
rect 1967 4870 1977 4922
rect 2001 4870 2031 4922
rect 2031 4870 2043 4922
rect 2043 4870 2057 4922
rect 2081 4870 2095 4922
rect 2095 4870 2107 4922
rect 2107 4870 2137 4922
rect 2161 4870 2171 4922
rect 2171 4870 2217 4922
rect 1921 4868 1977 4870
rect 2001 4868 2057 4870
rect 2081 4868 2137 4870
rect 2161 4868 2217 4870
rect 1582 4800 1638 4856
rect 3852 4922 3908 4924
rect 3932 4922 3988 4924
rect 4012 4922 4068 4924
rect 4092 4922 4148 4924
rect 3852 4870 3898 4922
rect 3898 4870 3908 4922
rect 3932 4870 3962 4922
rect 3962 4870 3974 4922
rect 3974 4870 3988 4922
rect 4012 4870 4026 4922
rect 4026 4870 4038 4922
rect 4038 4870 4068 4922
rect 4092 4870 4102 4922
rect 4102 4870 4148 4922
rect 3852 4868 3908 4870
rect 3932 4868 3988 4870
rect 4012 4868 4068 4870
rect 4092 4868 4148 4870
rect 1398 4004 1454 4040
rect 1398 3984 1400 4004
rect 1400 3984 1452 4004
rect 1452 3984 1454 4004
rect 1921 3834 1977 3836
rect 2001 3834 2057 3836
rect 2081 3834 2137 3836
rect 2161 3834 2217 3836
rect 1921 3782 1967 3834
rect 1967 3782 1977 3834
rect 2001 3782 2031 3834
rect 2031 3782 2043 3834
rect 2043 3782 2057 3834
rect 2081 3782 2095 3834
rect 2095 3782 2107 3834
rect 2107 3782 2137 3834
rect 2161 3782 2171 3834
rect 2171 3782 2217 3834
rect 1921 3780 1977 3782
rect 2001 3780 2057 3782
rect 2081 3780 2137 3782
rect 2161 3780 2217 3782
rect 1582 3304 1638 3360
rect 1398 2488 1454 2544
rect 1921 2746 1977 2748
rect 2001 2746 2057 2748
rect 2081 2746 2137 2748
rect 2161 2746 2217 2748
rect 1921 2694 1967 2746
rect 1967 2694 1977 2746
rect 2001 2694 2031 2746
rect 2031 2694 2043 2746
rect 2043 2694 2057 2746
rect 2081 2694 2095 2746
rect 2095 2694 2107 2746
rect 2107 2694 2137 2746
rect 2161 2694 2171 2746
rect 2171 2694 2217 2746
rect 1921 2692 1977 2694
rect 2001 2692 2057 2694
rect 2081 2692 2137 2694
rect 2161 2692 2217 2694
rect 2886 4378 2942 4380
rect 2966 4378 3022 4380
rect 3046 4378 3102 4380
rect 3126 4378 3182 4380
rect 2886 4326 2932 4378
rect 2932 4326 2942 4378
rect 2966 4326 2996 4378
rect 2996 4326 3008 4378
rect 3008 4326 3022 4378
rect 3046 4326 3060 4378
rect 3060 4326 3072 4378
rect 3072 4326 3102 4378
rect 3126 4326 3136 4378
rect 3136 4326 3182 4378
rect 2886 4324 2942 4326
rect 2966 4324 3022 4326
rect 3046 4324 3102 4326
rect 3126 4324 3182 4326
rect 3852 3834 3908 3836
rect 3932 3834 3988 3836
rect 4012 3834 4068 3836
rect 4092 3834 4148 3836
rect 3852 3782 3898 3834
rect 3898 3782 3908 3834
rect 3932 3782 3962 3834
rect 3962 3782 3974 3834
rect 3974 3782 3988 3834
rect 4012 3782 4026 3834
rect 4026 3782 4038 3834
rect 4038 3782 4068 3834
rect 4092 3782 4102 3834
rect 4102 3782 4148 3834
rect 3852 3780 3908 3782
rect 3932 3780 3988 3782
rect 4012 3780 4068 3782
rect 4092 3780 4148 3782
rect 2886 3290 2942 3292
rect 2966 3290 3022 3292
rect 3046 3290 3102 3292
rect 3126 3290 3182 3292
rect 2886 3238 2932 3290
rect 2932 3238 2942 3290
rect 2966 3238 2996 3290
rect 2996 3238 3008 3290
rect 3008 3238 3022 3290
rect 3046 3238 3060 3290
rect 3060 3238 3072 3290
rect 3072 3238 3102 3290
rect 3126 3238 3136 3290
rect 3136 3238 3182 3290
rect 2886 3236 2942 3238
rect 2966 3236 3022 3238
rect 3046 3236 3102 3238
rect 3126 3236 3182 3238
rect 3852 2746 3908 2748
rect 3932 2746 3988 2748
rect 4012 2746 4068 2748
rect 4092 2746 4148 2748
rect 3852 2694 3898 2746
rect 3898 2694 3908 2746
rect 3932 2694 3962 2746
rect 3962 2694 3974 2746
rect 3974 2694 3988 2746
rect 4012 2694 4026 2746
rect 4026 2694 4038 2746
rect 4038 2694 4068 2746
rect 4092 2694 4102 2746
rect 4102 2694 4148 2746
rect 3852 2692 3908 2694
rect 3932 2692 3988 2694
rect 4012 2692 4068 2694
rect 4092 2692 4148 2694
rect 1490 1808 1546 1864
rect 1582 992 1638 1048
rect 2886 2202 2942 2204
rect 2966 2202 3022 2204
rect 3046 2202 3102 2204
rect 3126 2202 3182 2204
rect 2886 2150 2932 2202
rect 2932 2150 2942 2202
rect 2966 2150 2996 2202
rect 2996 2150 3008 2202
rect 3008 2150 3022 2202
rect 3046 2150 3060 2202
rect 3060 2150 3072 2202
rect 3072 2150 3102 2202
rect 3126 2150 3136 2202
rect 3136 2150 3182 2202
rect 2886 2148 2942 2150
rect 2966 2148 3022 2150
rect 3046 2148 3102 2150
rect 3126 2148 3182 2150
rect 4817 6554 4873 6556
rect 4897 6554 4953 6556
rect 4977 6554 5033 6556
rect 5057 6554 5113 6556
rect 4817 6502 4863 6554
rect 4863 6502 4873 6554
rect 4897 6502 4927 6554
rect 4927 6502 4939 6554
rect 4939 6502 4953 6554
rect 4977 6502 4991 6554
rect 4991 6502 5003 6554
rect 5003 6502 5033 6554
rect 5057 6502 5067 6554
rect 5067 6502 5113 6554
rect 4817 6500 4873 6502
rect 4897 6500 4953 6502
rect 4977 6500 5033 6502
rect 5057 6500 5113 6502
rect 5262 6432 5318 6488
rect 4526 3576 4582 3632
rect 4817 5466 4873 5468
rect 4897 5466 4953 5468
rect 4977 5466 5033 5468
rect 5057 5466 5113 5468
rect 4817 5414 4863 5466
rect 4863 5414 4873 5466
rect 4897 5414 4927 5466
rect 4927 5414 4939 5466
rect 4939 5414 4953 5466
rect 4977 5414 4991 5466
rect 4991 5414 5003 5466
rect 5003 5414 5033 5466
rect 5057 5414 5067 5466
rect 5067 5414 5113 5466
rect 4817 5412 4873 5414
rect 4897 5412 4953 5414
rect 4977 5412 5033 5414
rect 5057 5412 5113 5414
rect 5782 7098 5838 7100
rect 5862 7098 5918 7100
rect 5942 7098 5998 7100
rect 6022 7098 6078 7100
rect 5782 7046 5828 7098
rect 5828 7046 5838 7098
rect 5862 7046 5892 7098
rect 5892 7046 5904 7098
rect 5904 7046 5918 7098
rect 5942 7046 5956 7098
rect 5956 7046 5968 7098
rect 5968 7046 5998 7098
rect 6022 7046 6032 7098
rect 6032 7046 6078 7098
rect 5782 7044 5838 7046
rect 5862 7044 5918 7046
rect 5942 7044 5998 7046
rect 6022 7044 6078 7046
rect 6918 8744 6974 8780
rect 5782 6010 5838 6012
rect 5862 6010 5918 6012
rect 5942 6010 5998 6012
rect 6022 6010 6078 6012
rect 5782 5958 5828 6010
rect 5828 5958 5838 6010
rect 5862 5958 5892 6010
rect 5892 5958 5904 6010
rect 5904 5958 5918 6010
rect 5942 5958 5956 6010
rect 5956 5958 5968 6010
rect 5968 5958 5998 6010
rect 6022 5958 6032 6010
rect 6032 5958 6078 6010
rect 5782 5956 5838 5958
rect 5862 5956 5918 5958
rect 5942 5956 5998 5958
rect 6022 5956 6078 5958
rect 7010 7012 7012 7032
rect 7012 7012 7064 7032
rect 7064 7012 7066 7032
rect 7010 6976 7066 7012
rect 7010 5924 7012 5944
rect 7012 5924 7064 5944
rect 7064 5924 7066 5944
rect 7010 5888 7066 5924
rect 5446 5072 5502 5128
rect 5782 4922 5838 4924
rect 5862 4922 5918 4924
rect 5942 4922 5998 4924
rect 6022 4922 6078 4924
rect 5782 4870 5828 4922
rect 5828 4870 5838 4922
rect 5862 4870 5892 4922
rect 5892 4870 5904 4922
rect 5904 4870 5918 4922
rect 5942 4870 5956 4922
rect 5956 4870 5968 4922
rect 5968 4870 5998 4922
rect 6022 4870 6032 4922
rect 6032 4870 6078 4922
rect 5782 4868 5838 4870
rect 5862 4868 5918 4870
rect 5942 4868 5998 4870
rect 6022 4868 6078 4870
rect 4817 4378 4873 4380
rect 4897 4378 4953 4380
rect 4977 4378 5033 4380
rect 5057 4378 5113 4380
rect 4817 4326 4863 4378
rect 4863 4326 4873 4378
rect 4897 4326 4927 4378
rect 4927 4326 4939 4378
rect 4939 4326 4953 4378
rect 4977 4326 4991 4378
rect 4991 4326 5003 4378
rect 5003 4326 5033 4378
rect 5057 4326 5067 4378
rect 5067 4326 5113 4378
rect 4817 4324 4873 4326
rect 4897 4324 4953 4326
rect 4977 4324 5033 4326
rect 5057 4324 5113 4326
rect 5262 4256 5318 4312
rect 4817 3290 4873 3292
rect 4897 3290 4953 3292
rect 4977 3290 5033 3292
rect 5057 3290 5113 3292
rect 4817 3238 4863 3290
rect 4863 3238 4873 3290
rect 4897 3238 4927 3290
rect 4927 3238 4939 3290
rect 4939 3238 4953 3290
rect 4977 3238 4991 3290
rect 4991 3238 5003 3290
rect 5003 3238 5033 3290
rect 5057 3238 5067 3290
rect 5067 3238 5113 3290
rect 4817 3236 4873 3238
rect 4897 3236 4953 3238
rect 4977 3236 5033 3238
rect 5057 3236 5113 3238
rect 5170 2488 5226 2544
rect 5782 3834 5838 3836
rect 5862 3834 5918 3836
rect 5942 3834 5998 3836
rect 6022 3834 6078 3836
rect 5782 3782 5828 3834
rect 5828 3782 5838 3834
rect 5862 3782 5892 3834
rect 5892 3782 5904 3834
rect 5904 3782 5918 3834
rect 5942 3782 5956 3834
rect 5956 3782 5968 3834
rect 5968 3782 5998 3834
rect 6022 3782 6032 3834
rect 6032 3782 6078 3834
rect 5782 3780 5838 3782
rect 5862 3780 5918 3782
rect 5942 3780 5998 3782
rect 6022 3780 6078 3782
rect 5998 3032 6054 3088
rect 5782 2746 5838 2748
rect 5862 2746 5918 2748
rect 5942 2746 5998 2748
rect 6022 2746 6078 2748
rect 5782 2694 5828 2746
rect 5828 2694 5838 2746
rect 5862 2694 5892 2746
rect 5892 2694 5904 2746
rect 5904 2694 5918 2746
rect 5942 2694 5956 2746
rect 5956 2694 5968 2746
rect 5968 2694 5998 2746
rect 6022 2694 6032 2746
rect 6032 2694 6078 2746
rect 5782 2692 5838 2694
rect 5862 2692 5918 2694
rect 5942 2692 5998 2694
rect 6022 2692 6078 2694
rect 4817 2202 4873 2204
rect 4897 2202 4953 2204
rect 4977 2202 5033 2204
rect 5057 2202 5113 2204
rect 4817 2150 4863 2202
rect 4863 2150 4873 2202
rect 4897 2150 4927 2202
rect 4927 2150 4939 2202
rect 4939 2150 4953 2202
rect 4977 2150 4991 2202
rect 4991 2150 5003 2202
rect 5003 2150 5033 2202
rect 5057 2150 5067 2202
rect 5067 2150 5113 2202
rect 4817 2148 4873 2150
rect 4897 2148 4953 2150
rect 4977 2148 5033 2150
rect 5057 2148 5113 2150
rect 5170 1400 5226 1456
rect 6182 1944 6238 2000
rect 5814 856 5870 912
rect 2778 312 2834 368
rect 4250 312 4306 368
<< metal3 >>
rect 4521 59666 4587 59669
rect 7200 59666 8000 59696
rect 4521 59664 8000 59666
rect 4521 59608 4526 59664
rect 4582 59608 8000 59664
rect 4521 59606 8000 59608
rect 4521 59603 4587 59606
rect 7200 59576 8000 59606
rect 0 59530 800 59560
rect 3325 59530 3391 59533
rect 0 59528 3391 59530
rect 0 59472 3330 59528
rect 3386 59472 3391 59528
rect 0 59470 3391 59472
rect 0 59440 800 59470
rect 3325 59467 3391 59470
rect 4245 59122 4311 59125
rect 7200 59122 8000 59152
rect 4245 59120 8000 59122
rect 4245 59064 4250 59120
rect 4306 59064 8000 59120
rect 4245 59062 8000 59064
rect 4245 59059 4311 59062
rect 7200 59032 8000 59062
rect 0 58714 800 58744
rect 3233 58714 3299 58717
rect 0 58712 3299 58714
rect 0 58656 3238 58712
rect 3294 58656 3299 58712
rect 0 58654 3299 58656
rect 0 58624 800 58654
rect 3233 58651 3299 58654
rect 5257 58578 5323 58581
rect 7200 58578 8000 58608
rect 5257 58576 8000 58578
rect 5257 58520 5262 58576
rect 5318 58520 8000 58576
rect 5257 58518 8000 58520
rect 5257 58515 5323 58518
rect 7200 58488 8000 58518
rect 0 58034 800 58064
rect 2773 58034 2839 58037
rect 0 58032 2839 58034
rect 0 57976 2778 58032
rect 2834 57976 2839 58032
rect 0 57974 2839 57976
rect 0 57944 800 57974
rect 2773 57971 2839 57974
rect 5441 58034 5507 58037
rect 7200 58034 8000 58064
rect 5441 58032 8000 58034
rect 5441 57976 5446 58032
rect 5502 57976 8000 58032
rect 5441 57974 8000 57976
rect 5441 57971 5507 57974
rect 7200 57944 8000 57974
rect 2874 57696 3194 57697
rect 2874 57632 2882 57696
rect 2946 57632 2962 57696
rect 3026 57632 3042 57696
rect 3106 57632 3122 57696
rect 3186 57632 3194 57696
rect 2874 57631 3194 57632
rect 4805 57696 5125 57697
rect 4805 57632 4813 57696
rect 4877 57632 4893 57696
rect 4957 57632 4973 57696
rect 5037 57632 5053 57696
rect 5117 57632 5125 57696
rect 4805 57631 5125 57632
rect 6269 57490 6335 57493
rect 7200 57490 8000 57520
rect 6269 57488 8000 57490
rect 6269 57432 6274 57488
rect 6330 57432 8000 57488
rect 6269 57430 8000 57432
rect 6269 57427 6335 57430
rect 7200 57400 8000 57430
rect 0 57218 800 57248
rect 1577 57218 1643 57221
rect 0 57216 1643 57218
rect 0 57160 1582 57216
rect 1638 57160 1643 57216
rect 0 57158 1643 57160
rect 0 57128 800 57158
rect 1577 57155 1643 57158
rect 1909 57152 2229 57153
rect 1909 57088 1917 57152
rect 1981 57088 1997 57152
rect 2061 57088 2077 57152
rect 2141 57088 2157 57152
rect 2221 57088 2229 57152
rect 1909 57087 2229 57088
rect 3840 57152 4160 57153
rect 3840 57088 3848 57152
rect 3912 57088 3928 57152
rect 3992 57088 4008 57152
rect 4072 57088 4088 57152
rect 4152 57088 4160 57152
rect 3840 57087 4160 57088
rect 5770 57152 6090 57153
rect 5770 57088 5778 57152
rect 5842 57088 5858 57152
rect 5922 57088 5938 57152
rect 6002 57088 6018 57152
rect 6082 57088 6090 57152
rect 5770 57087 6090 57088
rect 6177 56946 6243 56949
rect 7200 56946 8000 56976
rect 6177 56944 8000 56946
rect 6177 56888 6182 56944
rect 6238 56888 8000 56944
rect 6177 56886 8000 56888
rect 6177 56883 6243 56886
rect 7200 56856 8000 56886
rect 2874 56608 3194 56609
rect 0 56538 800 56568
rect 2874 56544 2882 56608
rect 2946 56544 2962 56608
rect 3026 56544 3042 56608
rect 3106 56544 3122 56608
rect 3186 56544 3194 56608
rect 2874 56543 3194 56544
rect 4805 56608 5125 56609
rect 4805 56544 4813 56608
rect 4877 56544 4893 56608
rect 4957 56544 4973 56608
rect 5037 56544 5053 56608
rect 5117 56544 5125 56608
rect 4805 56543 5125 56544
rect 1577 56538 1643 56541
rect 0 56536 1643 56538
rect 0 56480 1582 56536
rect 1638 56480 1643 56536
rect 0 56478 1643 56480
rect 0 56448 800 56478
rect 1577 56475 1643 56478
rect 5717 56266 5783 56269
rect 7200 56266 8000 56296
rect 5717 56264 8000 56266
rect 5717 56208 5722 56264
rect 5778 56208 8000 56264
rect 5717 56206 8000 56208
rect 5717 56203 5783 56206
rect 7200 56176 8000 56206
rect 1909 56064 2229 56065
rect 1909 56000 1917 56064
rect 1981 56000 1997 56064
rect 2061 56000 2077 56064
rect 2141 56000 2157 56064
rect 2221 56000 2229 56064
rect 1909 55999 2229 56000
rect 3840 56064 4160 56065
rect 3840 56000 3848 56064
rect 3912 56000 3928 56064
rect 3992 56000 4008 56064
rect 4072 56000 4088 56064
rect 4152 56000 4160 56064
rect 3840 55999 4160 56000
rect 5770 56064 6090 56065
rect 5770 56000 5778 56064
rect 5842 56000 5858 56064
rect 5922 56000 5938 56064
rect 6002 56000 6018 56064
rect 6082 56000 6090 56064
rect 5770 55999 6090 56000
rect 0 55722 800 55752
rect 1577 55722 1643 55725
rect 0 55720 1643 55722
rect 0 55664 1582 55720
rect 1638 55664 1643 55720
rect 0 55662 1643 55664
rect 0 55632 800 55662
rect 1577 55659 1643 55662
rect 5993 55722 6059 55725
rect 7200 55722 8000 55752
rect 5993 55720 8000 55722
rect 5993 55664 5998 55720
rect 6054 55664 8000 55720
rect 5993 55662 8000 55664
rect 5993 55659 6059 55662
rect 7200 55632 8000 55662
rect 2874 55520 3194 55521
rect 2874 55456 2882 55520
rect 2946 55456 2962 55520
rect 3026 55456 3042 55520
rect 3106 55456 3122 55520
rect 3186 55456 3194 55520
rect 2874 55455 3194 55456
rect 4805 55520 5125 55521
rect 4805 55456 4813 55520
rect 4877 55456 4893 55520
rect 4957 55456 4973 55520
rect 5037 55456 5053 55520
rect 5117 55456 5125 55520
rect 4805 55455 5125 55456
rect 4245 55316 4311 55317
rect 4245 55312 4292 55316
rect 4356 55314 4362 55316
rect 4245 55256 4250 55312
rect 4245 55252 4292 55256
rect 4356 55254 4402 55314
rect 4356 55252 4362 55254
rect 4245 55251 4311 55252
rect 5717 55178 5783 55181
rect 7200 55178 8000 55208
rect 5717 55176 8000 55178
rect 5717 55120 5722 55176
rect 5778 55120 8000 55176
rect 5717 55118 8000 55120
rect 5717 55115 5783 55118
rect 7200 55088 8000 55118
rect 1909 54976 2229 54977
rect 0 54906 800 54936
rect 1909 54912 1917 54976
rect 1981 54912 1997 54976
rect 2061 54912 2077 54976
rect 2141 54912 2157 54976
rect 2221 54912 2229 54976
rect 1909 54911 2229 54912
rect 3840 54976 4160 54977
rect 3840 54912 3848 54976
rect 3912 54912 3928 54976
rect 3992 54912 4008 54976
rect 4072 54912 4088 54976
rect 4152 54912 4160 54976
rect 3840 54911 4160 54912
rect 5770 54976 6090 54977
rect 5770 54912 5778 54976
rect 5842 54912 5858 54976
rect 5922 54912 5938 54976
rect 6002 54912 6018 54976
rect 6082 54912 6090 54976
rect 5770 54911 6090 54912
rect 1577 54906 1643 54909
rect 0 54904 1643 54906
rect 0 54848 1582 54904
rect 1638 54848 1643 54904
rect 0 54846 1643 54848
rect 0 54816 800 54846
rect 1577 54843 1643 54846
rect 5993 54634 6059 54637
rect 7200 54634 8000 54664
rect 5993 54632 8000 54634
rect 5993 54576 5998 54632
rect 6054 54576 8000 54632
rect 5993 54574 8000 54576
rect 5993 54571 6059 54574
rect 7200 54544 8000 54574
rect 2874 54432 3194 54433
rect 2874 54368 2882 54432
rect 2946 54368 2962 54432
rect 3026 54368 3042 54432
rect 3106 54368 3122 54432
rect 3186 54368 3194 54432
rect 2874 54367 3194 54368
rect 4805 54432 5125 54433
rect 4805 54368 4813 54432
rect 4877 54368 4893 54432
rect 4957 54368 4973 54432
rect 5037 54368 5053 54432
rect 5117 54368 5125 54432
rect 4805 54367 5125 54368
rect 0 54226 800 54256
rect 1577 54226 1643 54229
rect 0 54224 1643 54226
rect 0 54168 1582 54224
rect 1638 54168 1643 54224
rect 0 54166 1643 54168
rect 0 54136 800 54166
rect 1577 54163 1643 54166
rect 5717 54090 5783 54093
rect 7200 54090 8000 54120
rect 5717 54088 8000 54090
rect 5717 54032 5722 54088
rect 5778 54032 8000 54088
rect 5717 54030 8000 54032
rect 5717 54027 5783 54030
rect 7200 54000 8000 54030
rect 1909 53888 2229 53889
rect 1909 53824 1917 53888
rect 1981 53824 1997 53888
rect 2061 53824 2077 53888
rect 2141 53824 2157 53888
rect 2221 53824 2229 53888
rect 1909 53823 2229 53824
rect 3840 53888 4160 53889
rect 3840 53824 3848 53888
rect 3912 53824 3928 53888
rect 3992 53824 4008 53888
rect 4072 53824 4088 53888
rect 4152 53824 4160 53888
rect 3840 53823 4160 53824
rect 5770 53888 6090 53889
rect 5770 53824 5778 53888
rect 5842 53824 5858 53888
rect 5922 53824 5938 53888
rect 6002 53824 6018 53888
rect 6082 53824 6090 53888
rect 5770 53823 6090 53824
rect 5993 53546 6059 53549
rect 7200 53546 8000 53576
rect 5993 53544 8000 53546
rect 5993 53488 5998 53544
rect 6054 53488 8000 53544
rect 5993 53486 8000 53488
rect 5993 53483 6059 53486
rect 7200 53456 8000 53486
rect 0 53410 800 53440
rect 1577 53410 1643 53413
rect 0 53408 1643 53410
rect 0 53352 1582 53408
rect 1638 53352 1643 53408
rect 0 53350 1643 53352
rect 0 53320 800 53350
rect 1577 53347 1643 53350
rect 2874 53344 3194 53345
rect 2874 53280 2882 53344
rect 2946 53280 2962 53344
rect 3026 53280 3042 53344
rect 3106 53280 3122 53344
rect 3186 53280 3194 53344
rect 2874 53279 3194 53280
rect 4805 53344 5125 53345
rect 4805 53280 4813 53344
rect 4877 53280 4893 53344
rect 4957 53280 4973 53344
rect 5037 53280 5053 53344
rect 5117 53280 5125 53344
rect 4805 53279 5125 53280
rect 6177 52866 6243 52869
rect 7200 52866 8000 52896
rect 6177 52864 8000 52866
rect 6177 52808 6182 52864
rect 6238 52808 8000 52864
rect 6177 52806 8000 52808
rect 6177 52803 6243 52806
rect 1909 52800 2229 52801
rect 0 52730 800 52760
rect 1909 52736 1917 52800
rect 1981 52736 1997 52800
rect 2061 52736 2077 52800
rect 2141 52736 2157 52800
rect 2221 52736 2229 52800
rect 1909 52735 2229 52736
rect 3840 52800 4160 52801
rect 3840 52736 3848 52800
rect 3912 52736 3928 52800
rect 3992 52736 4008 52800
rect 4072 52736 4088 52800
rect 4152 52736 4160 52800
rect 3840 52735 4160 52736
rect 5770 52800 6090 52801
rect 5770 52736 5778 52800
rect 5842 52736 5858 52800
rect 5922 52736 5938 52800
rect 6002 52736 6018 52800
rect 6082 52736 6090 52800
rect 7200 52776 8000 52806
rect 5770 52735 6090 52736
rect 1577 52730 1643 52733
rect 0 52728 1643 52730
rect 0 52672 1582 52728
rect 1638 52672 1643 52728
rect 0 52670 1643 52672
rect 0 52640 800 52670
rect 1577 52667 1643 52670
rect 5993 52322 6059 52325
rect 7200 52322 8000 52352
rect 5993 52320 8000 52322
rect 5993 52264 5998 52320
rect 6054 52264 8000 52320
rect 5993 52262 8000 52264
rect 5993 52259 6059 52262
rect 2874 52256 3194 52257
rect 2874 52192 2882 52256
rect 2946 52192 2962 52256
rect 3026 52192 3042 52256
rect 3106 52192 3122 52256
rect 3186 52192 3194 52256
rect 2874 52191 3194 52192
rect 4805 52256 5125 52257
rect 4805 52192 4813 52256
rect 4877 52192 4893 52256
rect 4957 52192 4973 52256
rect 5037 52192 5053 52256
rect 5117 52192 5125 52256
rect 7200 52232 8000 52262
rect 4805 52191 5125 52192
rect 0 51914 800 51944
rect 1577 51914 1643 51917
rect 0 51912 1643 51914
rect 0 51856 1582 51912
rect 1638 51856 1643 51912
rect 0 51854 1643 51856
rect 0 51824 800 51854
rect 1577 51851 1643 51854
rect 6177 51778 6243 51781
rect 7200 51778 8000 51808
rect 6177 51776 8000 51778
rect 6177 51720 6182 51776
rect 6238 51720 8000 51776
rect 6177 51718 8000 51720
rect 6177 51715 6243 51718
rect 1909 51712 2229 51713
rect 1909 51648 1917 51712
rect 1981 51648 1997 51712
rect 2061 51648 2077 51712
rect 2141 51648 2157 51712
rect 2221 51648 2229 51712
rect 1909 51647 2229 51648
rect 3840 51712 4160 51713
rect 3840 51648 3848 51712
rect 3912 51648 3928 51712
rect 3992 51648 4008 51712
rect 4072 51648 4088 51712
rect 4152 51648 4160 51712
rect 3840 51647 4160 51648
rect 5770 51712 6090 51713
rect 5770 51648 5778 51712
rect 5842 51648 5858 51712
rect 5922 51648 5938 51712
rect 6002 51648 6018 51712
rect 6082 51648 6090 51712
rect 7200 51688 8000 51718
rect 5770 51647 6090 51648
rect 0 51234 800 51264
rect 1577 51234 1643 51237
rect 0 51232 1643 51234
rect 0 51176 1582 51232
rect 1638 51176 1643 51232
rect 0 51174 1643 51176
rect 0 51144 800 51174
rect 1577 51171 1643 51174
rect 5993 51234 6059 51237
rect 7200 51234 8000 51264
rect 5993 51232 8000 51234
rect 5993 51176 5998 51232
rect 6054 51176 8000 51232
rect 5993 51174 8000 51176
rect 5993 51171 6059 51174
rect 2874 51168 3194 51169
rect 2874 51104 2882 51168
rect 2946 51104 2962 51168
rect 3026 51104 3042 51168
rect 3106 51104 3122 51168
rect 3186 51104 3194 51168
rect 2874 51103 3194 51104
rect 4805 51168 5125 51169
rect 4805 51104 4813 51168
rect 4877 51104 4893 51168
rect 4957 51104 4973 51168
rect 5037 51104 5053 51168
rect 5117 51104 5125 51168
rect 7200 51144 8000 51174
rect 4805 51103 5125 51104
rect 6361 50690 6427 50693
rect 7200 50690 8000 50720
rect 6361 50688 8000 50690
rect 6361 50632 6366 50688
rect 6422 50632 8000 50688
rect 6361 50630 8000 50632
rect 6361 50627 6427 50630
rect 1909 50624 2229 50625
rect 1909 50560 1917 50624
rect 1981 50560 1997 50624
rect 2061 50560 2077 50624
rect 2141 50560 2157 50624
rect 2221 50560 2229 50624
rect 1909 50559 2229 50560
rect 3840 50624 4160 50625
rect 3840 50560 3848 50624
rect 3912 50560 3928 50624
rect 3992 50560 4008 50624
rect 4072 50560 4088 50624
rect 4152 50560 4160 50624
rect 3840 50559 4160 50560
rect 5770 50624 6090 50625
rect 5770 50560 5778 50624
rect 5842 50560 5858 50624
rect 5922 50560 5938 50624
rect 6002 50560 6018 50624
rect 6082 50560 6090 50624
rect 7200 50600 8000 50630
rect 5770 50559 6090 50560
rect 0 50418 800 50448
rect 1577 50418 1643 50421
rect 0 50416 1643 50418
rect 0 50360 1582 50416
rect 1638 50360 1643 50416
rect 0 50358 1643 50360
rect 0 50328 800 50358
rect 1577 50355 1643 50358
rect 5993 50146 6059 50149
rect 7200 50146 8000 50176
rect 5993 50144 8000 50146
rect 5993 50088 5998 50144
rect 6054 50088 8000 50144
rect 5993 50086 8000 50088
rect 5993 50083 6059 50086
rect 2874 50080 3194 50081
rect 2874 50016 2882 50080
rect 2946 50016 2962 50080
rect 3026 50016 3042 50080
rect 3106 50016 3122 50080
rect 3186 50016 3194 50080
rect 2874 50015 3194 50016
rect 4805 50080 5125 50081
rect 4805 50016 4813 50080
rect 4877 50016 4893 50080
rect 4957 50016 4973 50080
rect 5037 50016 5053 50080
rect 5117 50016 5125 50080
rect 7200 50056 8000 50086
rect 4805 50015 5125 50016
rect 0 49602 800 49632
rect 1577 49602 1643 49605
rect 0 49600 1643 49602
rect 0 49544 1582 49600
rect 1638 49544 1643 49600
rect 0 49542 1643 49544
rect 0 49512 800 49542
rect 1577 49539 1643 49542
rect 1909 49536 2229 49537
rect 1909 49472 1917 49536
rect 1981 49472 1997 49536
rect 2061 49472 2077 49536
rect 2141 49472 2157 49536
rect 2221 49472 2229 49536
rect 1909 49471 2229 49472
rect 3840 49536 4160 49537
rect 3840 49472 3848 49536
rect 3912 49472 3928 49536
rect 3992 49472 4008 49536
rect 4072 49472 4088 49536
rect 4152 49472 4160 49536
rect 3840 49471 4160 49472
rect 5770 49536 6090 49537
rect 5770 49472 5778 49536
rect 5842 49472 5858 49536
rect 5922 49472 5938 49536
rect 6002 49472 6018 49536
rect 6082 49472 6090 49536
rect 5770 49471 6090 49472
rect 6177 49466 6243 49469
rect 7200 49466 8000 49496
rect 6177 49464 8000 49466
rect 6177 49408 6182 49464
rect 6238 49408 8000 49464
rect 6177 49406 8000 49408
rect 6177 49403 6243 49406
rect 7200 49376 8000 49406
rect 2874 48992 3194 48993
rect 0 48922 800 48952
rect 2874 48928 2882 48992
rect 2946 48928 2962 48992
rect 3026 48928 3042 48992
rect 3106 48928 3122 48992
rect 3186 48928 3194 48992
rect 2874 48927 3194 48928
rect 4805 48992 5125 48993
rect 4805 48928 4813 48992
rect 4877 48928 4893 48992
rect 4957 48928 4973 48992
rect 5037 48928 5053 48992
rect 5117 48928 5125 48992
rect 4805 48927 5125 48928
rect 1577 48922 1643 48925
rect 0 48920 1643 48922
rect 0 48864 1582 48920
rect 1638 48864 1643 48920
rect 0 48862 1643 48864
rect 0 48832 800 48862
rect 1577 48859 1643 48862
rect 5993 48922 6059 48925
rect 7200 48922 8000 48952
rect 5993 48920 8000 48922
rect 5993 48864 5998 48920
rect 6054 48864 8000 48920
rect 5993 48862 8000 48864
rect 5993 48859 6059 48862
rect 7200 48832 8000 48862
rect 1909 48448 2229 48449
rect 1909 48384 1917 48448
rect 1981 48384 1997 48448
rect 2061 48384 2077 48448
rect 2141 48384 2157 48448
rect 2221 48384 2229 48448
rect 1909 48383 2229 48384
rect 3840 48448 4160 48449
rect 3840 48384 3848 48448
rect 3912 48384 3928 48448
rect 3992 48384 4008 48448
rect 4072 48384 4088 48448
rect 4152 48384 4160 48448
rect 3840 48383 4160 48384
rect 5770 48448 6090 48449
rect 5770 48384 5778 48448
rect 5842 48384 5858 48448
rect 5922 48384 5938 48448
rect 6002 48384 6018 48448
rect 6082 48384 6090 48448
rect 5770 48383 6090 48384
rect 6177 48378 6243 48381
rect 7200 48378 8000 48408
rect 6177 48376 8000 48378
rect 6177 48320 6182 48376
rect 6238 48320 8000 48376
rect 6177 48318 8000 48320
rect 6177 48315 6243 48318
rect 7200 48288 8000 48318
rect 0 48106 800 48136
rect 1577 48106 1643 48109
rect 0 48104 1643 48106
rect 0 48048 1582 48104
rect 1638 48048 1643 48104
rect 0 48046 1643 48048
rect 0 48016 800 48046
rect 1577 48043 1643 48046
rect 2630 48044 2636 48108
rect 2700 48106 2706 48108
rect 2865 48106 2931 48109
rect 2700 48104 2931 48106
rect 2700 48048 2870 48104
rect 2926 48048 2931 48104
rect 2700 48046 2931 48048
rect 2700 48044 2706 48046
rect 2865 48043 2931 48046
rect 4797 48106 4863 48109
rect 5390 48106 5396 48108
rect 4797 48104 5396 48106
rect 4797 48048 4802 48104
rect 4858 48048 5396 48104
rect 4797 48046 5396 48048
rect 4797 48043 4863 48046
rect 5390 48044 5396 48046
rect 5460 48044 5466 48108
rect 2874 47904 3194 47905
rect 2874 47840 2882 47904
rect 2946 47840 2962 47904
rect 3026 47840 3042 47904
rect 3106 47840 3122 47904
rect 3186 47840 3194 47904
rect 2874 47839 3194 47840
rect 4805 47904 5125 47905
rect 4805 47840 4813 47904
rect 4877 47840 4893 47904
rect 4957 47840 4973 47904
rect 5037 47840 5053 47904
rect 5117 47840 5125 47904
rect 4805 47839 5125 47840
rect 4337 47834 4403 47837
rect 4654 47834 4660 47836
rect 4337 47832 4660 47834
rect 4337 47776 4342 47832
rect 4398 47776 4660 47832
rect 4337 47774 4660 47776
rect 4337 47771 4403 47774
rect 4654 47772 4660 47774
rect 4724 47772 4730 47836
rect 5993 47834 6059 47837
rect 7200 47834 8000 47864
rect 5993 47832 8000 47834
rect 5993 47776 5998 47832
rect 6054 47776 8000 47832
rect 5993 47774 8000 47776
rect 5993 47771 6059 47774
rect 7200 47744 8000 47774
rect 0 47426 800 47456
rect 1577 47426 1643 47429
rect 0 47424 1643 47426
rect 0 47368 1582 47424
rect 1638 47368 1643 47424
rect 0 47366 1643 47368
rect 0 47336 800 47366
rect 1577 47363 1643 47366
rect 1909 47360 2229 47361
rect 1909 47296 1917 47360
rect 1981 47296 1997 47360
rect 2061 47296 2077 47360
rect 2141 47296 2157 47360
rect 2221 47296 2229 47360
rect 1909 47295 2229 47296
rect 3840 47360 4160 47361
rect 3840 47296 3848 47360
rect 3912 47296 3928 47360
rect 3992 47296 4008 47360
rect 4072 47296 4088 47360
rect 4152 47296 4160 47360
rect 3840 47295 4160 47296
rect 5770 47360 6090 47361
rect 5770 47296 5778 47360
rect 5842 47296 5858 47360
rect 5922 47296 5938 47360
rect 6002 47296 6018 47360
rect 6082 47296 6090 47360
rect 5770 47295 6090 47296
rect 6177 47290 6243 47293
rect 7200 47290 8000 47320
rect 6177 47288 8000 47290
rect 6177 47232 6182 47288
rect 6238 47232 8000 47288
rect 6177 47230 8000 47232
rect 6177 47227 6243 47230
rect 7200 47200 8000 47230
rect 2874 46816 3194 46817
rect 2874 46752 2882 46816
rect 2946 46752 2962 46816
rect 3026 46752 3042 46816
rect 3106 46752 3122 46816
rect 3186 46752 3194 46816
rect 2874 46751 3194 46752
rect 4805 46816 5125 46817
rect 4805 46752 4813 46816
rect 4877 46752 4893 46816
rect 4957 46752 4973 46816
rect 5037 46752 5053 46816
rect 5117 46752 5125 46816
rect 4805 46751 5125 46752
rect 5993 46746 6059 46749
rect 7200 46746 8000 46776
rect 5993 46744 8000 46746
rect 5993 46688 5998 46744
rect 6054 46688 8000 46744
rect 5993 46686 8000 46688
rect 5993 46683 6059 46686
rect 7200 46656 8000 46686
rect 0 46610 800 46640
rect 1577 46610 1643 46613
rect 0 46608 1643 46610
rect 0 46552 1582 46608
rect 1638 46552 1643 46608
rect 0 46550 1643 46552
rect 0 46520 800 46550
rect 1577 46547 1643 46550
rect 1909 46272 2229 46273
rect 1909 46208 1917 46272
rect 1981 46208 1997 46272
rect 2061 46208 2077 46272
rect 2141 46208 2157 46272
rect 2221 46208 2229 46272
rect 1909 46207 2229 46208
rect 3840 46272 4160 46273
rect 3840 46208 3848 46272
rect 3912 46208 3928 46272
rect 3992 46208 4008 46272
rect 4072 46208 4088 46272
rect 4152 46208 4160 46272
rect 3840 46207 4160 46208
rect 5770 46272 6090 46273
rect 5770 46208 5778 46272
rect 5842 46208 5858 46272
rect 5922 46208 5938 46272
rect 6002 46208 6018 46272
rect 6082 46208 6090 46272
rect 5770 46207 6090 46208
rect 6177 46066 6243 46069
rect 7200 46066 8000 46096
rect 6177 46064 8000 46066
rect 6177 46008 6182 46064
rect 6238 46008 8000 46064
rect 6177 46006 8000 46008
rect 6177 46003 6243 46006
rect 7200 45976 8000 46006
rect 0 45794 800 45824
rect 1577 45794 1643 45797
rect 0 45792 1643 45794
rect 0 45736 1582 45792
rect 1638 45736 1643 45792
rect 0 45734 1643 45736
rect 0 45704 800 45734
rect 1577 45731 1643 45734
rect 2874 45728 3194 45729
rect 2874 45664 2882 45728
rect 2946 45664 2962 45728
rect 3026 45664 3042 45728
rect 3106 45664 3122 45728
rect 3186 45664 3194 45728
rect 2874 45663 3194 45664
rect 4805 45728 5125 45729
rect 4805 45664 4813 45728
rect 4877 45664 4893 45728
rect 4957 45664 4973 45728
rect 5037 45664 5053 45728
rect 5117 45664 5125 45728
rect 4805 45663 5125 45664
rect 5993 45522 6059 45525
rect 7200 45522 8000 45552
rect 5993 45520 8000 45522
rect 5993 45464 5998 45520
rect 6054 45464 8000 45520
rect 5993 45462 8000 45464
rect 5993 45459 6059 45462
rect 7200 45432 8000 45462
rect 5206 45324 5212 45388
rect 5276 45386 5282 45388
rect 5809 45386 5875 45389
rect 5276 45384 5875 45386
rect 5276 45328 5814 45384
rect 5870 45328 5875 45384
rect 5276 45326 5875 45328
rect 5276 45324 5282 45326
rect 5809 45323 5875 45326
rect 1909 45184 2229 45185
rect 0 45114 800 45144
rect 1909 45120 1917 45184
rect 1981 45120 1997 45184
rect 2061 45120 2077 45184
rect 2141 45120 2157 45184
rect 2221 45120 2229 45184
rect 1909 45119 2229 45120
rect 3840 45184 4160 45185
rect 3840 45120 3848 45184
rect 3912 45120 3928 45184
rect 3992 45120 4008 45184
rect 4072 45120 4088 45184
rect 4152 45120 4160 45184
rect 3840 45119 4160 45120
rect 5770 45184 6090 45185
rect 5770 45120 5778 45184
rect 5842 45120 5858 45184
rect 5922 45120 5938 45184
rect 6002 45120 6018 45184
rect 6082 45120 6090 45184
rect 5770 45119 6090 45120
rect 1577 45114 1643 45117
rect 0 45112 1643 45114
rect 0 45056 1582 45112
rect 1638 45056 1643 45112
rect 0 45054 1643 45056
rect 0 45024 800 45054
rect 1577 45051 1643 45054
rect 6177 44978 6243 44981
rect 7200 44978 8000 45008
rect 6177 44976 8000 44978
rect 6177 44920 6182 44976
rect 6238 44920 8000 44976
rect 6177 44918 8000 44920
rect 6177 44915 6243 44918
rect 7200 44888 8000 44918
rect 2874 44640 3194 44641
rect 2874 44576 2882 44640
rect 2946 44576 2962 44640
rect 3026 44576 3042 44640
rect 3106 44576 3122 44640
rect 3186 44576 3194 44640
rect 2874 44575 3194 44576
rect 4805 44640 5125 44641
rect 4805 44576 4813 44640
rect 4877 44576 4893 44640
rect 4957 44576 4973 44640
rect 5037 44576 5053 44640
rect 5117 44576 5125 44640
rect 4805 44575 5125 44576
rect 5993 44434 6059 44437
rect 7200 44434 8000 44464
rect 5993 44432 8000 44434
rect 5993 44376 5998 44432
rect 6054 44376 8000 44432
rect 5993 44374 8000 44376
rect 5993 44371 6059 44374
rect 7200 44344 8000 44374
rect 0 44298 800 44328
rect 1577 44298 1643 44301
rect 0 44296 1643 44298
rect 0 44240 1582 44296
rect 1638 44240 1643 44296
rect 0 44238 1643 44240
rect 0 44208 800 44238
rect 1577 44235 1643 44238
rect 1909 44096 2229 44097
rect 1909 44032 1917 44096
rect 1981 44032 1997 44096
rect 2061 44032 2077 44096
rect 2141 44032 2157 44096
rect 2221 44032 2229 44096
rect 1909 44031 2229 44032
rect 3840 44096 4160 44097
rect 3840 44032 3848 44096
rect 3912 44032 3928 44096
rect 3992 44032 4008 44096
rect 4072 44032 4088 44096
rect 4152 44032 4160 44096
rect 3840 44031 4160 44032
rect 5770 44096 6090 44097
rect 5770 44032 5778 44096
rect 5842 44032 5858 44096
rect 5922 44032 5938 44096
rect 6002 44032 6018 44096
rect 6082 44032 6090 44096
rect 5770 44031 6090 44032
rect 5625 43890 5691 43893
rect 7200 43890 8000 43920
rect 5625 43888 8000 43890
rect 5625 43832 5630 43888
rect 5686 43832 8000 43888
rect 5625 43830 8000 43832
rect 5625 43827 5691 43830
rect 7200 43800 8000 43830
rect 3141 43754 3207 43757
rect 3366 43754 3372 43756
rect 3141 43752 3372 43754
rect 3141 43696 3146 43752
rect 3202 43696 3372 43752
rect 3141 43694 3372 43696
rect 3141 43691 3207 43694
rect 3366 43692 3372 43694
rect 3436 43692 3442 43756
rect 0 43618 800 43648
rect 1577 43618 1643 43621
rect 0 43616 1643 43618
rect 0 43560 1582 43616
rect 1638 43560 1643 43616
rect 0 43558 1643 43560
rect 0 43528 800 43558
rect 1577 43555 1643 43558
rect 2874 43552 3194 43553
rect 2874 43488 2882 43552
rect 2946 43488 2962 43552
rect 3026 43488 3042 43552
rect 3106 43488 3122 43552
rect 3186 43488 3194 43552
rect 2874 43487 3194 43488
rect 4805 43552 5125 43553
rect 4805 43488 4813 43552
rect 4877 43488 4893 43552
rect 4957 43488 4973 43552
rect 5037 43488 5053 43552
rect 5117 43488 5125 43552
rect 4805 43487 5125 43488
rect 4613 43346 4679 43349
rect 5574 43346 5580 43348
rect 4613 43344 5580 43346
rect 4613 43288 4618 43344
rect 4674 43288 5580 43344
rect 4613 43286 5580 43288
rect 4613 43283 4679 43286
rect 5574 43284 5580 43286
rect 5644 43284 5650 43348
rect 5993 43346 6059 43349
rect 7200 43346 8000 43376
rect 5993 43344 8000 43346
rect 5993 43288 5998 43344
rect 6054 43288 8000 43344
rect 5993 43286 8000 43288
rect 5993 43283 6059 43286
rect 7200 43256 8000 43286
rect 1909 43008 2229 43009
rect 1909 42944 1917 43008
rect 1981 42944 1997 43008
rect 2061 42944 2077 43008
rect 2141 42944 2157 43008
rect 2221 42944 2229 43008
rect 1909 42943 2229 42944
rect 3840 43008 4160 43009
rect 3840 42944 3848 43008
rect 3912 42944 3928 43008
rect 3992 42944 4008 43008
rect 4072 42944 4088 43008
rect 4152 42944 4160 43008
rect 3840 42943 4160 42944
rect 5770 43008 6090 43009
rect 5770 42944 5778 43008
rect 5842 42944 5858 43008
rect 5922 42944 5938 43008
rect 6002 42944 6018 43008
rect 6082 42944 6090 43008
rect 5770 42943 6090 42944
rect 0 42802 800 42832
rect 1577 42802 1643 42805
rect 0 42800 1643 42802
rect 0 42744 1582 42800
rect 1638 42744 1643 42800
rect 0 42742 1643 42744
rect 0 42712 800 42742
rect 1577 42739 1643 42742
rect 5625 42802 5691 42805
rect 7200 42802 8000 42832
rect 5625 42800 8000 42802
rect 5625 42744 5630 42800
rect 5686 42744 8000 42800
rect 5625 42742 8000 42744
rect 5625 42739 5691 42742
rect 7200 42712 8000 42742
rect 2874 42464 3194 42465
rect 2874 42400 2882 42464
rect 2946 42400 2962 42464
rect 3026 42400 3042 42464
rect 3106 42400 3122 42464
rect 3186 42400 3194 42464
rect 2874 42399 3194 42400
rect 4805 42464 5125 42465
rect 4805 42400 4813 42464
rect 4877 42400 4893 42464
rect 4957 42400 4973 42464
rect 5037 42400 5053 42464
rect 5117 42400 5125 42464
rect 4805 42399 5125 42400
rect 4654 42196 4660 42260
rect 4724 42258 4730 42260
rect 4797 42258 4863 42261
rect 4724 42256 4863 42258
rect 4724 42200 4802 42256
rect 4858 42200 4863 42256
rect 4724 42198 4863 42200
rect 4724 42196 4730 42198
rect 4797 42195 4863 42198
rect 0 42122 800 42152
rect 1577 42122 1643 42125
rect 0 42120 1643 42122
rect 0 42064 1582 42120
rect 1638 42064 1643 42120
rect 0 42062 1643 42064
rect 0 42032 800 42062
rect 1577 42059 1643 42062
rect 3550 42060 3556 42124
rect 3620 42122 3626 42124
rect 5257 42122 5323 42125
rect 3620 42120 5323 42122
rect 3620 42064 5262 42120
rect 5318 42064 5323 42120
rect 3620 42062 5323 42064
rect 3620 42060 3626 42062
rect 5257 42059 5323 42062
rect 5717 42122 5783 42125
rect 7200 42122 8000 42152
rect 5717 42120 8000 42122
rect 5717 42064 5722 42120
rect 5778 42064 8000 42120
rect 5717 42062 8000 42064
rect 5717 42059 5783 42062
rect 7200 42032 8000 42062
rect 4705 41988 4771 41989
rect 4654 41924 4660 41988
rect 4724 41986 4771 41988
rect 4724 41984 4816 41986
rect 4766 41928 4816 41984
rect 4724 41926 4816 41928
rect 4724 41924 4771 41926
rect 4705 41923 4771 41924
rect 1909 41920 2229 41921
rect 1909 41856 1917 41920
rect 1981 41856 1997 41920
rect 2061 41856 2077 41920
rect 2141 41856 2157 41920
rect 2221 41856 2229 41920
rect 1909 41855 2229 41856
rect 3840 41920 4160 41921
rect 3840 41856 3848 41920
rect 3912 41856 3928 41920
rect 3992 41856 4008 41920
rect 4072 41856 4088 41920
rect 4152 41856 4160 41920
rect 3840 41855 4160 41856
rect 5770 41920 6090 41921
rect 5770 41856 5778 41920
rect 5842 41856 5858 41920
rect 5922 41856 5938 41920
rect 6002 41856 6018 41920
rect 6082 41856 6090 41920
rect 5770 41855 6090 41856
rect 1485 41850 1551 41853
rect 4521 41852 4587 41853
rect 1485 41848 1594 41850
rect 1485 41792 1490 41848
rect 1546 41792 1594 41848
rect 1485 41787 1594 41792
rect 4470 41788 4476 41852
rect 4540 41850 4587 41852
rect 4540 41848 4632 41850
rect 4582 41792 4632 41848
rect 4540 41790 4632 41792
rect 4540 41788 4587 41790
rect 4521 41787 4587 41788
rect 1534 41445 1594 41787
rect 4337 41714 4403 41717
rect 4294 41712 4403 41714
rect 4294 41656 4342 41712
rect 4398 41656 4403 41712
rect 4294 41651 4403 41656
rect 4613 41714 4679 41717
rect 5390 41714 5396 41716
rect 4613 41712 5396 41714
rect 4613 41656 4618 41712
rect 4674 41656 5396 41712
rect 4613 41654 5396 41656
rect 4613 41651 4679 41654
rect 5390 41652 5396 41654
rect 5460 41652 5466 41716
rect 1710 41516 1716 41580
rect 1780 41578 1786 41580
rect 3509 41578 3575 41581
rect 1780 41576 3575 41578
rect 1780 41520 3514 41576
rect 3570 41520 3575 41576
rect 1780 41518 3575 41520
rect 1780 41516 1786 41518
rect 3509 41515 3575 41518
rect 1485 41440 1594 41445
rect 1485 41384 1490 41440
rect 1546 41384 1594 41440
rect 1485 41382 1594 41384
rect 1485 41379 1551 41382
rect 2874 41376 3194 41377
rect 0 41306 800 41336
rect 2874 41312 2882 41376
rect 2946 41312 2962 41376
rect 3026 41312 3042 41376
rect 3106 41312 3122 41376
rect 3186 41312 3194 41376
rect 2874 41311 3194 41312
rect 1577 41306 1643 41309
rect 0 41304 1643 41306
rect 0 41248 1582 41304
rect 1638 41248 1643 41304
rect 0 41246 1643 41248
rect 0 41216 800 41246
rect 1577 41243 1643 41246
rect 3233 41170 3299 41173
rect 3366 41170 3372 41172
rect 3233 41168 3372 41170
rect 3233 41112 3238 41168
rect 3294 41112 3372 41168
rect 3233 41110 3372 41112
rect 3233 41107 3299 41110
rect 3366 41108 3372 41110
rect 3436 41108 3442 41172
rect 4294 41034 4354 41651
rect 5257 41578 5323 41581
rect 7200 41578 8000 41608
rect 5257 41576 8000 41578
rect 5257 41520 5262 41576
rect 5318 41520 8000 41576
rect 5257 41518 8000 41520
rect 5257 41515 5323 41518
rect 7200 41488 8000 41518
rect 4805 41376 5125 41377
rect 4805 41312 4813 41376
rect 4877 41312 4893 41376
rect 4957 41312 4973 41376
rect 5037 41312 5053 41376
rect 5117 41312 5125 41376
rect 4805 41311 5125 41312
rect 4654 41244 4660 41308
rect 4724 41244 4730 41308
rect 4429 41170 4495 41173
rect 4662 41170 4722 41244
rect 4429 41168 4722 41170
rect 4429 41112 4434 41168
rect 4490 41112 4722 41168
rect 4429 41110 4722 41112
rect 4429 41107 4495 41110
rect 4470 41034 4476 41036
rect 4294 40974 4476 41034
rect 4470 40972 4476 40974
rect 4540 40972 4546 41036
rect 4981 41034 5047 41037
rect 7200 41034 8000 41064
rect 4981 41032 8000 41034
rect 4981 40976 4986 41032
rect 5042 40976 8000 41032
rect 4981 40974 8000 40976
rect 4981 40971 5047 40974
rect 7200 40944 8000 40974
rect 4245 40898 4311 40901
rect 5206 40898 5212 40900
rect 4245 40896 5212 40898
rect 4245 40840 4250 40896
rect 4306 40840 5212 40896
rect 4245 40838 5212 40840
rect 4245 40835 4311 40838
rect 5206 40836 5212 40838
rect 5276 40836 5282 40900
rect 1909 40832 2229 40833
rect 1909 40768 1917 40832
rect 1981 40768 1997 40832
rect 2061 40768 2077 40832
rect 2141 40768 2157 40832
rect 2221 40768 2229 40832
rect 1909 40767 2229 40768
rect 3840 40832 4160 40833
rect 3840 40768 3848 40832
rect 3912 40768 3928 40832
rect 3992 40768 4008 40832
rect 4072 40768 4088 40832
rect 4152 40768 4160 40832
rect 3840 40767 4160 40768
rect 5770 40832 6090 40833
rect 5770 40768 5778 40832
rect 5842 40768 5858 40832
rect 5922 40768 5938 40832
rect 6002 40768 6018 40832
rect 6082 40768 6090 40832
rect 5770 40767 6090 40768
rect 0 40490 800 40520
rect 1577 40490 1643 40493
rect 0 40488 1643 40490
rect 0 40432 1582 40488
rect 1638 40432 1643 40488
rect 0 40430 1643 40432
rect 0 40400 800 40430
rect 1577 40427 1643 40430
rect 5717 40490 5783 40493
rect 7200 40490 8000 40520
rect 5717 40488 8000 40490
rect 5717 40432 5722 40488
rect 5778 40432 8000 40488
rect 5717 40430 8000 40432
rect 5717 40427 5783 40430
rect 7200 40400 8000 40430
rect 2874 40288 3194 40289
rect 2874 40224 2882 40288
rect 2946 40224 2962 40288
rect 3026 40224 3042 40288
rect 3106 40224 3122 40288
rect 3186 40224 3194 40288
rect 2874 40223 3194 40224
rect 4805 40288 5125 40289
rect 4805 40224 4813 40288
rect 4877 40224 4893 40288
rect 4957 40224 4973 40288
rect 5037 40224 5053 40288
rect 5117 40224 5125 40288
rect 4805 40223 5125 40224
rect 5809 39946 5875 39949
rect 7200 39946 8000 39976
rect 5809 39944 8000 39946
rect 5809 39888 5814 39944
rect 5870 39888 8000 39944
rect 5809 39886 8000 39888
rect 5809 39883 5875 39886
rect 7200 39856 8000 39886
rect 0 39810 800 39840
rect 1577 39810 1643 39813
rect 0 39808 1643 39810
rect 0 39752 1582 39808
rect 1638 39752 1643 39808
rect 0 39750 1643 39752
rect 0 39720 800 39750
rect 1577 39747 1643 39750
rect 1909 39744 2229 39745
rect 1909 39680 1917 39744
rect 1981 39680 1997 39744
rect 2061 39680 2077 39744
rect 2141 39680 2157 39744
rect 2221 39680 2229 39744
rect 1909 39679 2229 39680
rect 3840 39744 4160 39745
rect 3840 39680 3848 39744
rect 3912 39680 3928 39744
rect 3992 39680 4008 39744
rect 4072 39680 4088 39744
rect 4152 39680 4160 39744
rect 3840 39679 4160 39680
rect 5770 39744 6090 39745
rect 5770 39680 5778 39744
rect 5842 39680 5858 39744
rect 5922 39680 5938 39744
rect 6002 39680 6018 39744
rect 6082 39680 6090 39744
rect 5770 39679 6090 39680
rect 6085 39402 6151 39405
rect 7200 39402 8000 39432
rect 6085 39400 8000 39402
rect 6085 39344 6090 39400
rect 6146 39344 8000 39400
rect 6085 39342 8000 39344
rect 6085 39339 6151 39342
rect 7200 39312 8000 39342
rect 2874 39200 3194 39201
rect 2874 39136 2882 39200
rect 2946 39136 2962 39200
rect 3026 39136 3042 39200
rect 3106 39136 3122 39200
rect 3186 39136 3194 39200
rect 2874 39135 3194 39136
rect 4805 39200 5125 39201
rect 4805 39136 4813 39200
rect 4877 39136 4893 39200
rect 4957 39136 4973 39200
rect 5037 39136 5053 39200
rect 5117 39136 5125 39200
rect 4805 39135 5125 39136
rect 0 38994 800 39024
rect 1577 38994 1643 38997
rect 0 38992 1643 38994
rect 0 38936 1582 38992
rect 1638 38936 1643 38992
rect 0 38934 1643 38936
rect 0 38904 800 38934
rect 1577 38931 1643 38934
rect 2630 38932 2636 38996
rect 2700 38994 2706 38996
rect 3141 38994 3207 38997
rect 2700 38992 3207 38994
rect 2700 38936 3146 38992
rect 3202 38936 3207 38992
rect 2700 38934 3207 38936
rect 2700 38932 2706 38934
rect 3141 38931 3207 38934
rect 5073 38994 5139 38997
rect 5574 38994 5580 38996
rect 5073 38992 5580 38994
rect 5073 38936 5078 38992
rect 5134 38936 5580 38992
rect 5073 38934 5580 38936
rect 5073 38931 5139 38934
rect 5574 38932 5580 38934
rect 5644 38932 5650 38996
rect 2405 38722 2471 38725
rect 2630 38722 2636 38724
rect 2405 38720 2636 38722
rect 2405 38664 2410 38720
rect 2466 38664 2636 38720
rect 2405 38662 2636 38664
rect 2405 38659 2471 38662
rect 2630 38660 2636 38662
rect 2700 38660 2706 38724
rect 6177 38722 6243 38725
rect 7200 38722 8000 38752
rect 6177 38720 8000 38722
rect 3509 38670 3575 38673
rect 3374 38668 3575 38670
rect 1909 38656 2229 38657
rect 1909 38592 1917 38656
rect 1981 38592 1997 38656
rect 2061 38592 2077 38656
rect 2141 38592 2157 38656
rect 2221 38592 2229 38656
rect 1909 38591 2229 38592
rect 3374 38612 3514 38668
rect 3570 38612 3575 38668
rect 6177 38664 6182 38720
rect 6238 38664 8000 38720
rect 6177 38662 8000 38664
rect 6177 38659 6243 38662
rect 3374 38610 3575 38612
rect 2446 38524 2452 38588
rect 2516 38586 2522 38588
rect 3374 38586 3434 38610
rect 3509 38607 3575 38610
rect 3840 38656 4160 38657
rect 3840 38592 3848 38656
rect 3912 38592 3928 38656
rect 3992 38592 4008 38656
rect 4072 38592 4088 38656
rect 4152 38592 4160 38656
rect 3840 38591 4160 38592
rect 5770 38656 6090 38657
rect 5770 38592 5778 38656
rect 5842 38592 5858 38656
rect 5922 38592 5938 38656
rect 6002 38592 6018 38656
rect 6082 38592 6090 38656
rect 7200 38632 8000 38662
rect 5770 38591 6090 38592
rect 2516 38526 3434 38586
rect 2516 38524 2522 38526
rect 2589 38450 2655 38453
rect 5625 38450 5691 38453
rect 2589 38448 5691 38450
rect 2589 38392 2594 38448
rect 2650 38392 5630 38448
rect 5686 38392 5691 38448
rect 2589 38390 5691 38392
rect 2589 38387 2655 38390
rect 5625 38387 5691 38390
rect 0 38314 800 38344
rect 1577 38314 1643 38317
rect 0 38312 1643 38314
rect 0 38256 1582 38312
rect 1638 38256 1643 38312
rect 0 38254 1643 38256
rect 0 38224 800 38254
rect 1577 38251 1643 38254
rect 3366 38252 3372 38316
rect 3436 38314 3442 38316
rect 5073 38314 5139 38317
rect 3436 38312 5139 38314
rect 3436 38256 5078 38312
rect 5134 38256 5139 38312
rect 3436 38254 5139 38256
rect 3436 38252 3442 38254
rect 5073 38251 5139 38254
rect 6085 38178 6151 38181
rect 7200 38178 8000 38208
rect 6085 38176 8000 38178
rect 6085 38120 6090 38176
rect 6146 38120 8000 38176
rect 6085 38118 8000 38120
rect 6085 38115 6151 38118
rect 2874 38112 3194 38113
rect 2874 38048 2882 38112
rect 2946 38048 2962 38112
rect 3026 38048 3042 38112
rect 3106 38048 3122 38112
rect 3186 38048 3194 38112
rect 2874 38047 3194 38048
rect 4805 38112 5125 38113
rect 4805 38048 4813 38112
rect 4877 38048 4893 38112
rect 4957 38048 4973 38112
rect 5037 38048 5053 38112
rect 5117 38048 5125 38112
rect 7200 38088 8000 38118
rect 4805 38047 5125 38048
rect 1710 37844 1716 37908
rect 1780 37906 1786 37908
rect 3509 37906 3575 37909
rect 1780 37904 3575 37906
rect 1780 37848 3514 37904
rect 3570 37848 3575 37904
rect 1780 37846 3575 37848
rect 1780 37844 1786 37846
rect 3509 37843 3575 37846
rect 4981 37770 5047 37773
rect 4981 37768 6378 37770
rect 4981 37712 4986 37768
rect 5042 37712 6378 37768
rect 4981 37710 6378 37712
rect 4981 37707 5047 37710
rect 6318 37634 6378 37710
rect 7200 37634 8000 37664
rect 6318 37574 8000 37634
rect 1909 37568 2229 37569
rect 0 37498 800 37528
rect 1909 37504 1917 37568
rect 1981 37504 1997 37568
rect 2061 37504 2077 37568
rect 2141 37504 2157 37568
rect 2221 37504 2229 37568
rect 1909 37503 2229 37504
rect 3840 37568 4160 37569
rect 3840 37504 3848 37568
rect 3912 37504 3928 37568
rect 3992 37504 4008 37568
rect 4072 37504 4088 37568
rect 4152 37504 4160 37568
rect 3840 37503 4160 37504
rect 5770 37568 6090 37569
rect 5770 37504 5778 37568
rect 5842 37504 5858 37568
rect 5922 37504 5938 37568
rect 6002 37504 6018 37568
rect 6082 37504 6090 37568
rect 7200 37544 8000 37574
rect 5770 37503 6090 37504
rect 1577 37498 1643 37501
rect 0 37496 1643 37498
rect 0 37440 1582 37496
rect 1638 37440 1643 37496
rect 0 37438 1643 37440
rect 0 37408 800 37438
rect 1577 37435 1643 37438
rect 5257 37090 5323 37093
rect 7200 37090 8000 37120
rect 5257 37088 8000 37090
rect 5257 37032 5262 37088
rect 5318 37032 8000 37088
rect 5257 37030 8000 37032
rect 5257 37027 5323 37030
rect 2874 37024 3194 37025
rect 2874 36960 2882 37024
rect 2946 36960 2962 37024
rect 3026 36960 3042 37024
rect 3106 36960 3122 37024
rect 3186 36960 3194 37024
rect 2874 36959 3194 36960
rect 4805 37024 5125 37025
rect 4805 36960 4813 37024
rect 4877 36960 4893 37024
rect 4957 36960 4973 37024
rect 5037 36960 5053 37024
rect 5117 36960 5125 37024
rect 7200 37000 8000 37030
rect 4805 36959 5125 36960
rect 2681 36956 2747 36957
rect 2630 36954 2636 36956
rect 2590 36894 2636 36954
rect 2700 36952 2747 36956
rect 2742 36896 2747 36952
rect 2630 36892 2636 36894
rect 2700 36892 2747 36896
rect 2681 36891 2747 36892
rect 0 36682 800 36712
rect 1577 36682 1643 36685
rect 0 36680 1643 36682
rect 0 36624 1582 36680
rect 1638 36624 1643 36680
rect 0 36622 1643 36624
rect 0 36592 800 36622
rect 1577 36619 1643 36622
rect 4981 36682 5047 36685
rect 4981 36680 6378 36682
rect 4981 36624 4986 36680
rect 5042 36624 6378 36680
rect 4981 36622 6378 36624
rect 4981 36619 5047 36622
rect 6318 36546 6378 36622
rect 7200 36546 8000 36576
rect 6318 36486 8000 36546
rect 1909 36480 2229 36481
rect 1909 36416 1917 36480
rect 1981 36416 1997 36480
rect 2061 36416 2077 36480
rect 2141 36416 2157 36480
rect 2221 36416 2229 36480
rect 1909 36415 2229 36416
rect 3840 36480 4160 36481
rect 3840 36416 3848 36480
rect 3912 36416 3928 36480
rect 3992 36416 4008 36480
rect 4072 36416 4088 36480
rect 4152 36416 4160 36480
rect 3840 36415 4160 36416
rect 5770 36480 6090 36481
rect 5770 36416 5778 36480
rect 5842 36416 5858 36480
rect 5922 36416 5938 36480
rect 6002 36416 6018 36480
rect 6082 36416 6090 36480
rect 7200 36456 8000 36486
rect 5770 36415 6090 36416
rect 0 36002 800 36032
rect 1301 36002 1367 36005
rect 0 36000 1367 36002
rect 0 35944 1306 36000
rect 1362 35944 1367 36000
rect 0 35942 1367 35944
rect 0 35912 800 35942
rect 1301 35939 1367 35942
rect 5257 36002 5323 36005
rect 7200 36002 8000 36032
rect 5257 36000 8000 36002
rect 5257 35944 5262 36000
rect 5318 35944 8000 36000
rect 5257 35942 8000 35944
rect 5257 35939 5323 35942
rect 2874 35936 3194 35937
rect 2874 35872 2882 35936
rect 2946 35872 2962 35936
rect 3026 35872 3042 35936
rect 3106 35872 3122 35936
rect 3186 35872 3194 35936
rect 2874 35871 3194 35872
rect 4805 35936 5125 35937
rect 4805 35872 4813 35936
rect 4877 35872 4893 35936
rect 4957 35872 4973 35936
rect 5037 35872 5053 35936
rect 5117 35872 5125 35936
rect 7200 35912 8000 35942
rect 4805 35871 5125 35872
rect 4981 35594 5047 35597
rect 4981 35592 6378 35594
rect 4981 35536 4986 35592
rect 5042 35536 6378 35592
rect 4981 35534 6378 35536
rect 4981 35531 5047 35534
rect 1909 35392 2229 35393
rect 1909 35328 1917 35392
rect 1981 35328 1997 35392
rect 2061 35328 2077 35392
rect 2141 35328 2157 35392
rect 2221 35328 2229 35392
rect 1909 35327 2229 35328
rect 3840 35392 4160 35393
rect 3840 35328 3848 35392
rect 3912 35328 3928 35392
rect 3992 35328 4008 35392
rect 4072 35328 4088 35392
rect 4152 35328 4160 35392
rect 3840 35327 4160 35328
rect 5770 35392 6090 35393
rect 5770 35328 5778 35392
rect 5842 35328 5858 35392
rect 5922 35328 5938 35392
rect 6002 35328 6018 35392
rect 6082 35328 6090 35392
rect 5770 35327 6090 35328
rect 6318 35322 6378 35534
rect 7200 35322 8000 35352
rect 6318 35262 8000 35322
rect 7200 35232 8000 35262
rect 0 35186 800 35216
rect 1393 35186 1459 35189
rect 0 35184 1459 35186
rect 0 35128 1398 35184
rect 1454 35128 1459 35184
rect 0 35126 1459 35128
rect 0 35096 800 35126
rect 1393 35123 1459 35126
rect 2874 34848 3194 34849
rect 2874 34784 2882 34848
rect 2946 34784 2962 34848
rect 3026 34784 3042 34848
rect 3106 34784 3122 34848
rect 3186 34784 3194 34848
rect 2874 34783 3194 34784
rect 4805 34848 5125 34849
rect 4805 34784 4813 34848
rect 4877 34784 4893 34848
rect 4957 34784 4973 34848
rect 5037 34784 5053 34848
rect 5117 34784 5125 34848
rect 4805 34783 5125 34784
rect 5257 34778 5323 34781
rect 7200 34778 8000 34808
rect 5257 34776 8000 34778
rect 5257 34720 5262 34776
rect 5318 34720 8000 34776
rect 5257 34718 8000 34720
rect 5257 34715 5323 34718
rect 7200 34688 8000 34718
rect 0 34506 800 34536
rect 1853 34506 1919 34509
rect 0 34504 1919 34506
rect 0 34448 1858 34504
rect 1914 34448 1919 34504
rect 0 34446 1919 34448
rect 0 34416 800 34446
rect 1853 34443 1919 34446
rect 4337 34506 4403 34509
rect 4470 34506 4476 34508
rect 4337 34504 4476 34506
rect 4337 34448 4342 34504
rect 4398 34448 4476 34504
rect 4337 34446 4476 34448
rect 4337 34443 4403 34446
rect 4470 34444 4476 34446
rect 4540 34444 4546 34508
rect 4981 34506 5047 34509
rect 4981 34504 6378 34506
rect 4981 34448 4986 34504
rect 5042 34448 6378 34504
rect 4981 34446 6378 34448
rect 4981 34443 5047 34446
rect 1669 34370 1735 34373
rect 1534 34368 1735 34370
rect 1534 34312 1674 34368
rect 1730 34312 1735 34368
rect 1534 34310 1735 34312
rect 1534 34101 1594 34310
rect 1669 34307 1735 34310
rect 1909 34304 2229 34305
rect 1909 34240 1917 34304
rect 1981 34240 1997 34304
rect 2061 34240 2077 34304
rect 2141 34240 2157 34304
rect 2221 34240 2229 34304
rect 1909 34239 2229 34240
rect 3840 34304 4160 34305
rect 3840 34240 3848 34304
rect 3912 34240 3928 34304
rect 3992 34240 4008 34304
rect 4072 34240 4088 34304
rect 4152 34240 4160 34304
rect 3840 34239 4160 34240
rect 5770 34304 6090 34305
rect 5770 34240 5778 34304
rect 5842 34240 5858 34304
rect 5922 34240 5938 34304
rect 6002 34240 6018 34304
rect 6082 34240 6090 34304
rect 5770 34239 6090 34240
rect 6318 34234 6378 34446
rect 7200 34234 8000 34264
rect 6318 34174 8000 34234
rect 7200 34144 8000 34174
rect 1534 34096 1643 34101
rect 1534 34040 1582 34096
rect 1638 34040 1643 34096
rect 1534 34038 1643 34040
rect 1577 34035 1643 34038
rect 2874 33760 3194 33761
rect 0 33690 800 33720
rect 2874 33696 2882 33760
rect 2946 33696 2962 33760
rect 3026 33696 3042 33760
rect 3106 33696 3122 33760
rect 3186 33696 3194 33760
rect 2874 33695 3194 33696
rect 4805 33760 5125 33761
rect 4805 33696 4813 33760
rect 4877 33696 4893 33760
rect 4957 33696 4973 33760
rect 5037 33696 5053 33760
rect 5117 33696 5125 33760
rect 4805 33695 5125 33696
rect 1853 33690 1919 33693
rect 0 33688 1919 33690
rect 0 33632 1858 33688
rect 1914 33632 1919 33688
rect 0 33630 1919 33632
rect 0 33600 800 33630
rect 1853 33627 1919 33630
rect 5257 33690 5323 33693
rect 7200 33690 8000 33720
rect 5257 33688 8000 33690
rect 5257 33632 5262 33688
rect 5318 33632 8000 33688
rect 5257 33630 8000 33632
rect 5257 33627 5323 33630
rect 7200 33600 8000 33630
rect 1909 33216 2229 33217
rect 1909 33152 1917 33216
rect 1981 33152 1997 33216
rect 2061 33152 2077 33216
rect 2141 33152 2157 33216
rect 2221 33152 2229 33216
rect 1909 33151 2229 33152
rect 3840 33216 4160 33217
rect 3840 33152 3848 33216
rect 3912 33152 3928 33216
rect 3992 33152 4008 33216
rect 4072 33152 4088 33216
rect 4152 33152 4160 33216
rect 3840 33151 4160 33152
rect 5770 33216 6090 33217
rect 5770 33152 5778 33216
rect 5842 33152 5858 33216
rect 5922 33152 5938 33216
rect 6002 33152 6018 33216
rect 6082 33152 6090 33216
rect 5770 33151 6090 33152
rect 7200 33146 8000 33176
rect 6318 33086 8000 33146
rect 0 33010 800 33040
rect 1393 33010 1459 33013
rect 0 33008 1459 33010
rect 0 32952 1398 33008
rect 1454 32952 1459 33008
rect 0 32950 1459 32952
rect 0 32920 800 32950
rect 1393 32947 1459 32950
rect 4981 33010 5047 33013
rect 6318 33010 6378 33086
rect 7200 33056 8000 33086
rect 4981 33008 6378 33010
rect 4981 32952 4986 33008
rect 5042 32952 6378 33008
rect 4981 32950 6378 32952
rect 4981 32947 5047 32950
rect 2037 32874 2103 32877
rect 4286 32874 4292 32876
rect 2037 32872 4292 32874
rect 2037 32816 2042 32872
rect 2098 32816 4292 32872
rect 2037 32814 4292 32816
rect 2037 32811 2103 32814
rect 4286 32812 4292 32814
rect 4356 32812 4362 32876
rect 2874 32672 3194 32673
rect 2874 32608 2882 32672
rect 2946 32608 2962 32672
rect 3026 32608 3042 32672
rect 3106 32608 3122 32672
rect 3186 32608 3194 32672
rect 2874 32607 3194 32608
rect 4805 32672 5125 32673
rect 4805 32608 4813 32672
rect 4877 32608 4893 32672
rect 4957 32608 4973 32672
rect 5037 32608 5053 32672
rect 5117 32608 5125 32672
rect 4805 32607 5125 32608
rect 5257 32602 5323 32605
rect 7200 32602 8000 32632
rect 5257 32600 8000 32602
rect 5257 32544 5262 32600
rect 5318 32544 8000 32600
rect 5257 32542 8000 32544
rect 5257 32539 5323 32542
rect 7200 32512 8000 32542
rect 4654 32268 4660 32332
rect 4724 32330 4730 32332
rect 5349 32330 5415 32333
rect 4724 32328 5415 32330
rect 4724 32272 5354 32328
rect 5410 32272 5415 32328
rect 4724 32270 5415 32272
rect 4724 32268 4730 32270
rect 5349 32267 5415 32270
rect 0 32194 800 32224
rect 1393 32194 1459 32197
rect 0 32192 1459 32194
rect 0 32136 1398 32192
rect 1454 32136 1459 32192
rect 0 32134 1459 32136
rect 0 32104 800 32134
rect 1393 32131 1459 32134
rect 1909 32128 2229 32129
rect 1909 32064 1917 32128
rect 1981 32064 1997 32128
rect 2061 32064 2077 32128
rect 2141 32064 2157 32128
rect 2221 32064 2229 32128
rect 1909 32063 2229 32064
rect 3840 32128 4160 32129
rect 3840 32064 3848 32128
rect 3912 32064 3928 32128
rect 3992 32064 4008 32128
rect 4072 32064 4088 32128
rect 4152 32064 4160 32128
rect 3840 32063 4160 32064
rect 5770 32128 6090 32129
rect 5770 32064 5778 32128
rect 5842 32064 5858 32128
rect 5922 32064 5938 32128
rect 6002 32064 6018 32128
rect 6082 32064 6090 32128
rect 5770 32063 6090 32064
rect 4981 31922 5047 31925
rect 7200 31922 8000 31952
rect 4981 31920 8000 31922
rect 4981 31864 4986 31920
rect 5042 31864 8000 31920
rect 4981 31862 8000 31864
rect 4981 31859 5047 31862
rect 7200 31832 8000 31862
rect 3550 31724 3556 31788
rect 3620 31786 3626 31788
rect 5349 31786 5415 31789
rect 3620 31784 5415 31786
rect 3620 31728 5354 31784
rect 5410 31728 5415 31784
rect 3620 31726 5415 31728
rect 3620 31724 3626 31726
rect 5349 31723 5415 31726
rect 2874 31584 3194 31585
rect 2874 31520 2882 31584
rect 2946 31520 2962 31584
rect 3026 31520 3042 31584
rect 3106 31520 3122 31584
rect 3186 31520 3194 31584
rect 2874 31519 3194 31520
rect 4805 31584 5125 31585
rect 4805 31520 4813 31584
rect 4877 31520 4893 31584
rect 4957 31520 4973 31584
rect 5037 31520 5053 31584
rect 5117 31520 5125 31584
rect 4805 31519 5125 31520
rect 0 31378 800 31408
rect 1853 31378 1919 31381
rect 0 31376 1919 31378
rect 0 31320 1858 31376
rect 1914 31320 1919 31376
rect 0 31318 1919 31320
rect 0 31288 800 31318
rect 1853 31315 1919 31318
rect 6821 31378 6887 31381
rect 7200 31378 8000 31408
rect 6821 31376 8000 31378
rect 6821 31320 6826 31376
rect 6882 31320 8000 31376
rect 6821 31318 8000 31320
rect 6821 31315 6887 31318
rect 7200 31288 8000 31318
rect 2405 31244 2471 31245
rect 2405 31240 2452 31244
rect 2516 31242 2522 31244
rect 2405 31184 2410 31240
rect 2405 31180 2452 31184
rect 2516 31182 2562 31242
rect 2516 31180 2522 31182
rect 2405 31179 2471 31180
rect 1909 31040 2229 31041
rect 1909 30976 1917 31040
rect 1981 30976 1997 31040
rect 2061 30976 2077 31040
rect 2141 30976 2157 31040
rect 2221 30976 2229 31040
rect 1909 30975 2229 30976
rect 3840 31040 4160 31041
rect 3840 30976 3848 31040
rect 3912 30976 3928 31040
rect 3992 30976 4008 31040
rect 4072 30976 4088 31040
rect 4152 30976 4160 31040
rect 3840 30975 4160 30976
rect 5770 31040 6090 31041
rect 5770 30976 5778 31040
rect 5842 30976 5858 31040
rect 5922 30976 5938 31040
rect 6002 30976 6018 31040
rect 6082 30976 6090 31040
rect 5770 30975 6090 30976
rect 6177 30834 6243 30837
rect 7200 30834 8000 30864
rect 6177 30832 8000 30834
rect 6177 30776 6182 30832
rect 6238 30776 8000 30832
rect 6177 30774 8000 30776
rect 6177 30771 6243 30774
rect 7200 30744 8000 30774
rect 0 30698 800 30728
rect 1393 30698 1459 30701
rect 0 30696 1459 30698
rect 0 30640 1398 30696
rect 1454 30640 1459 30696
rect 0 30638 1459 30640
rect 0 30608 800 30638
rect 1393 30635 1459 30638
rect 2874 30496 3194 30497
rect 2874 30432 2882 30496
rect 2946 30432 2962 30496
rect 3026 30432 3042 30496
rect 3106 30432 3122 30496
rect 3186 30432 3194 30496
rect 2874 30431 3194 30432
rect 4805 30496 5125 30497
rect 4805 30432 4813 30496
rect 4877 30432 4893 30496
rect 4957 30432 4973 30496
rect 5037 30432 5053 30496
rect 5117 30432 5125 30496
rect 4805 30431 5125 30432
rect 5441 30290 5507 30293
rect 7200 30290 8000 30320
rect 5441 30288 8000 30290
rect 5441 30232 5446 30288
rect 5502 30232 8000 30288
rect 5441 30230 8000 30232
rect 5441 30227 5507 30230
rect 7200 30200 8000 30230
rect 1909 29952 2229 29953
rect 0 29882 800 29912
rect 1909 29888 1917 29952
rect 1981 29888 1997 29952
rect 2061 29888 2077 29952
rect 2141 29888 2157 29952
rect 2221 29888 2229 29952
rect 1909 29887 2229 29888
rect 3840 29952 4160 29953
rect 3840 29888 3848 29952
rect 3912 29888 3928 29952
rect 3992 29888 4008 29952
rect 4072 29888 4088 29952
rect 4152 29888 4160 29952
rect 3840 29887 4160 29888
rect 5770 29952 6090 29953
rect 5770 29888 5778 29952
rect 5842 29888 5858 29952
rect 5922 29888 5938 29952
rect 6002 29888 6018 29952
rect 6082 29888 6090 29952
rect 5770 29887 6090 29888
rect 1393 29882 1459 29885
rect 0 29880 1459 29882
rect 0 29824 1398 29880
rect 1454 29824 1459 29880
rect 0 29822 1459 29824
rect 0 29792 800 29822
rect 1393 29819 1459 29822
rect 2865 29882 2931 29885
rect 3366 29882 3372 29884
rect 2865 29880 3372 29882
rect 2865 29824 2870 29880
rect 2926 29824 3372 29880
rect 2865 29822 3372 29824
rect 2865 29819 2931 29822
rect 3366 29820 3372 29822
rect 3436 29820 3442 29884
rect 6177 29746 6243 29749
rect 7200 29746 8000 29776
rect 6177 29744 8000 29746
rect 6177 29688 6182 29744
rect 6238 29688 8000 29744
rect 6177 29686 8000 29688
rect 6177 29683 6243 29686
rect 7200 29656 8000 29686
rect 2874 29408 3194 29409
rect 2874 29344 2882 29408
rect 2946 29344 2962 29408
rect 3026 29344 3042 29408
rect 3106 29344 3122 29408
rect 3186 29344 3194 29408
rect 2874 29343 3194 29344
rect 4805 29408 5125 29409
rect 4805 29344 4813 29408
rect 4877 29344 4893 29408
rect 4957 29344 4973 29408
rect 5037 29344 5053 29408
rect 5117 29344 5125 29408
rect 4805 29343 5125 29344
rect 0 29202 800 29232
rect 1577 29202 1643 29205
rect 0 29200 1643 29202
rect 0 29144 1582 29200
rect 1638 29144 1643 29200
rect 0 29142 1643 29144
rect 0 29112 800 29142
rect 1577 29139 1643 29142
rect 5257 29202 5323 29205
rect 7200 29202 8000 29232
rect 5257 29200 8000 29202
rect 5257 29144 5262 29200
rect 5318 29144 8000 29200
rect 5257 29142 8000 29144
rect 5257 29139 5323 29142
rect 7200 29112 8000 29142
rect 1909 28864 2229 28865
rect 1909 28800 1917 28864
rect 1981 28800 1997 28864
rect 2061 28800 2077 28864
rect 2141 28800 2157 28864
rect 2221 28800 2229 28864
rect 1909 28799 2229 28800
rect 3840 28864 4160 28865
rect 3840 28800 3848 28864
rect 3912 28800 3928 28864
rect 3992 28800 4008 28864
rect 4072 28800 4088 28864
rect 4152 28800 4160 28864
rect 3840 28799 4160 28800
rect 5770 28864 6090 28865
rect 5770 28800 5778 28864
rect 5842 28800 5858 28864
rect 5922 28800 5938 28864
rect 6002 28800 6018 28864
rect 6082 28800 6090 28864
rect 5770 28799 6090 28800
rect 4981 28658 5047 28661
rect 7200 28658 8000 28688
rect 4981 28656 8000 28658
rect 4981 28600 4986 28656
rect 5042 28600 8000 28656
rect 4981 28598 8000 28600
rect 4981 28595 5047 28598
rect 7200 28568 8000 28598
rect 0 28386 800 28416
rect 1393 28386 1459 28389
rect 0 28384 1459 28386
rect 0 28328 1398 28384
rect 1454 28328 1459 28384
rect 0 28326 1459 28328
rect 0 28296 800 28326
rect 1393 28323 1459 28326
rect 2874 28320 3194 28321
rect 2874 28256 2882 28320
rect 2946 28256 2962 28320
rect 3026 28256 3042 28320
rect 3106 28256 3122 28320
rect 3186 28256 3194 28320
rect 2874 28255 3194 28256
rect 4805 28320 5125 28321
rect 4805 28256 4813 28320
rect 4877 28256 4893 28320
rect 4957 28256 4973 28320
rect 5037 28256 5053 28320
rect 5117 28256 5125 28320
rect 4805 28255 5125 28256
rect 6085 27978 6151 27981
rect 7200 27978 8000 28008
rect 6085 27976 8000 27978
rect 6085 27920 6090 27976
rect 6146 27920 8000 27976
rect 6085 27918 8000 27920
rect 6085 27915 6151 27918
rect 7200 27888 8000 27918
rect 1909 27776 2229 27777
rect 1909 27712 1917 27776
rect 1981 27712 1997 27776
rect 2061 27712 2077 27776
rect 2141 27712 2157 27776
rect 2221 27712 2229 27776
rect 1909 27711 2229 27712
rect 3840 27776 4160 27777
rect 3840 27712 3848 27776
rect 3912 27712 3928 27776
rect 3992 27712 4008 27776
rect 4072 27712 4088 27776
rect 4152 27712 4160 27776
rect 3840 27711 4160 27712
rect 5770 27776 6090 27777
rect 5770 27712 5778 27776
rect 5842 27712 5858 27776
rect 5922 27712 5938 27776
rect 6002 27712 6018 27776
rect 6082 27712 6090 27776
rect 5770 27711 6090 27712
rect 0 27570 800 27600
rect 2773 27570 2839 27573
rect 0 27568 2839 27570
rect 0 27512 2778 27568
rect 2834 27512 2839 27568
rect 0 27510 2839 27512
rect 0 27480 800 27510
rect 2773 27507 2839 27510
rect 6177 27434 6243 27437
rect 7200 27434 8000 27464
rect 6177 27432 8000 27434
rect 6177 27376 6182 27432
rect 6238 27376 8000 27432
rect 6177 27374 8000 27376
rect 6177 27371 6243 27374
rect 7200 27344 8000 27374
rect 2874 27232 3194 27233
rect 2874 27168 2882 27232
rect 2946 27168 2962 27232
rect 3026 27168 3042 27232
rect 3106 27168 3122 27232
rect 3186 27168 3194 27232
rect 2874 27167 3194 27168
rect 4805 27232 5125 27233
rect 4805 27168 4813 27232
rect 4877 27168 4893 27232
rect 4957 27168 4973 27232
rect 5037 27168 5053 27232
rect 5117 27168 5125 27232
rect 4805 27167 5125 27168
rect 0 26890 800 26920
rect 1577 26890 1643 26893
rect 0 26888 1643 26890
rect 0 26832 1582 26888
rect 1638 26832 1643 26888
rect 0 26830 1643 26832
rect 0 26800 800 26830
rect 1577 26827 1643 26830
rect 5073 26890 5139 26893
rect 7200 26890 8000 26920
rect 5073 26888 8000 26890
rect 5073 26832 5078 26888
rect 5134 26832 8000 26888
rect 5073 26830 8000 26832
rect 5073 26827 5139 26830
rect 7200 26800 8000 26830
rect 1909 26688 2229 26689
rect 1909 26624 1917 26688
rect 1981 26624 1997 26688
rect 2061 26624 2077 26688
rect 2141 26624 2157 26688
rect 2221 26624 2229 26688
rect 1909 26623 2229 26624
rect 3840 26688 4160 26689
rect 3840 26624 3848 26688
rect 3912 26624 3928 26688
rect 3992 26624 4008 26688
rect 4072 26624 4088 26688
rect 4152 26624 4160 26688
rect 3840 26623 4160 26624
rect 5770 26688 6090 26689
rect 5770 26624 5778 26688
rect 5842 26624 5858 26688
rect 5922 26624 5938 26688
rect 6002 26624 6018 26688
rect 6082 26624 6090 26688
rect 5770 26623 6090 26624
rect 5441 26346 5507 26349
rect 7200 26346 8000 26376
rect 5441 26344 8000 26346
rect 5441 26288 5446 26344
rect 5502 26288 8000 26344
rect 5441 26286 8000 26288
rect 5441 26283 5507 26286
rect 7200 26256 8000 26286
rect 2874 26144 3194 26145
rect 0 26074 800 26104
rect 2874 26080 2882 26144
rect 2946 26080 2962 26144
rect 3026 26080 3042 26144
rect 3106 26080 3122 26144
rect 3186 26080 3194 26144
rect 2874 26079 3194 26080
rect 4805 26144 5125 26145
rect 4805 26080 4813 26144
rect 4877 26080 4893 26144
rect 4957 26080 4973 26144
rect 5037 26080 5053 26144
rect 5117 26080 5125 26144
rect 4805 26079 5125 26080
rect 1577 26074 1643 26077
rect 0 26072 1643 26074
rect 0 26016 1582 26072
rect 1638 26016 1643 26072
rect 0 26014 1643 26016
rect 0 25984 800 26014
rect 1577 26011 1643 26014
rect 6821 25802 6887 25805
rect 7200 25802 8000 25832
rect 6821 25800 8000 25802
rect 6821 25744 6826 25800
rect 6882 25744 8000 25800
rect 6821 25742 8000 25744
rect 6821 25739 6887 25742
rect 7200 25712 8000 25742
rect 1909 25600 2229 25601
rect 1909 25536 1917 25600
rect 1981 25536 1997 25600
rect 2061 25536 2077 25600
rect 2141 25536 2157 25600
rect 2221 25536 2229 25600
rect 1909 25535 2229 25536
rect 3840 25600 4160 25601
rect 3840 25536 3848 25600
rect 3912 25536 3928 25600
rect 3992 25536 4008 25600
rect 4072 25536 4088 25600
rect 4152 25536 4160 25600
rect 3840 25535 4160 25536
rect 5770 25600 6090 25601
rect 5770 25536 5778 25600
rect 5842 25536 5858 25600
rect 5922 25536 5938 25600
rect 6002 25536 6018 25600
rect 6082 25536 6090 25600
rect 5770 25535 6090 25536
rect 0 25394 800 25424
rect 1577 25394 1643 25397
rect 0 25392 1643 25394
rect 0 25336 1582 25392
rect 1638 25336 1643 25392
rect 0 25334 1643 25336
rect 0 25304 800 25334
rect 1577 25331 1643 25334
rect 6085 25258 6151 25261
rect 7200 25258 8000 25288
rect 6085 25256 8000 25258
rect 6085 25200 6090 25256
rect 6146 25200 8000 25256
rect 6085 25198 8000 25200
rect 6085 25195 6151 25198
rect 7200 25168 8000 25198
rect 2874 25056 3194 25057
rect 2874 24992 2882 25056
rect 2946 24992 2962 25056
rect 3026 24992 3042 25056
rect 3106 24992 3122 25056
rect 3186 24992 3194 25056
rect 2874 24991 3194 24992
rect 4805 25056 5125 25057
rect 4805 24992 4813 25056
rect 4877 24992 4893 25056
rect 4957 24992 4973 25056
rect 5037 24992 5053 25056
rect 5117 24992 5125 25056
rect 4805 24991 5125 24992
rect 0 24578 800 24608
rect 1577 24578 1643 24581
rect 0 24576 1643 24578
rect 0 24520 1582 24576
rect 1638 24520 1643 24576
rect 0 24518 1643 24520
rect 0 24488 800 24518
rect 1577 24515 1643 24518
rect 6177 24578 6243 24581
rect 7200 24578 8000 24608
rect 6177 24576 8000 24578
rect 6177 24520 6182 24576
rect 6238 24520 8000 24576
rect 6177 24518 8000 24520
rect 6177 24515 6243 24518
rect 1909 24512 2229 24513
rect 1909 24448 1917 24512
rect 1981 24448 1997 24512
rect 2061 24448 2077 24512
rect 2141 24448 2157 24512
rect 2221 24448 2229 24512
rect 1909 24447 2229 24448
rect 3840 24512 4160 24513
rect 3840 24448 3848 24512
rect 3912 24448 3928 24512
rect 3992 24448 4008 24512
rect 4072 24448 4088 24512
rect 4152 24448 4160 24512
rect 3840 24447 4160 24448
rect 5770 24512 6090 24513
rect 5770 24448 5778 24512
rect 5842 24448 5858 24512
rect 5922 24448 5938 24512
rect 6002 24448 6018 24512
rect 6082 24448 6090 24512
rect 7200 24488 8000 24518
rect 5770 24447 6090 24448
rect 5441 24034 5507 24037
rect 7200 24034 8000 24064
rect 5441 24032 8000 24034
rect 5441 23976 5446 24032
rect 5502 23976 8000 24032
rect 5441 23974 8000 23976
rect 5441 23971 5507 23974
rect 2874 23968 3194 23969
rect 0 23898 800 23928
rect 2874 23904 2882 23968
rect 2946 23904 2962 23968
rect 3026 23904 3042 23968
rect 3106 23904 3122 23968
rect 3186 23904 3194 23968
rect 2874 23903 3194 23904
rect 4805 23968 5125 23969
rect 4805 23904 4813 23968
rect 4877 23904 4893 23968
rect 4957 23904 4973 23968
rect 5037 23904 5053 23968
rect 5117 23904 5125 23968
rect 7200 23944 8000 23974
rect 4805 23903 5125 23904
rect 1577 23898 1643 23901
rect 0 23896 1643 23898
rect 0 23840 1582 23896
rect 1638 23840 1643 23896
rect 0 23838 1643 23840
rect 0 23808 800 23838
rect 1577 23835 1643 23838
rect 6177 23490 6243 23493
rect 7200 23490 8000 23520
rect 6177 23488 8000 23490
rect 6177 23432 6182 23488
rect 6238 23432 8000 23488
rect 6177 23430 8000 23432
rect 6177 23427 6243 23430
rect 1909 23424 2229 23425
rect 1909 23360 1917 23424
rect 1981 23360 1997 23424
rect 2061 23360 2077 23424
rect 2141 23360 2157 23424
rect 2221 23360 2229 23424
rect 1909 23359 2229 23360
rect 3840 23424 4160 23425
rect 3840 23360 3848 23424
rect 3912 23360 3928 23424
rect 3992 23360 4008 23424
rect 4072 23360 4088 23424
rect 4152 23360 4160 23424
rect 3840 23359 4160 23360
rect 5770 23424 6090 23425
rect 5770 23360 5778 23424
rect 5842 23360 5858 23424
rect 5922 23360 5938 23424
rect 6002 23360 6018 23424
rect 6082 23360 6090 23424
rect 7200 23400 8000 23430
rect 5770 23359 6090 23360
rect 0 23082 800 23112
rect 1577 23082 1643 23085
rect 0 23080 1643 23082
rect 0 23024 1582 23080
rect 1638 23024 1643 23080
rect 0 23022 1643 23024
rect 0 22992 800 23022
rect 1577 23019 1643 23022
rect 5257 22946 5323 22949
rect 7200 22946 8000 22976
rect 5257 22944 8000 22946
rect 5257 22888 5262 22944
rect 5318 22888 8000 22944
rect 5257 22886 8000 22888
rect 5257 22883 5323 22886
rect 2874 22880 3194 22881
rect 2874 22816 2882 22880
rect 2946 22816 2962 22880
rect 3026 22816 3042 22880
rect 3106 22816 3122 22880
rect 3186 22816 3194 22880
rect 2874 22815 3194 22816
rect 4805 22880 5125 22881
rect 4805 22816 4813 22880
rect 4877 22816 4893 22880
rect 4957 22816 4973 22880
rect 5037 22816 5053 22880
rect 5117 22816 5125 22880
rect 7200 22856 8000 22886
rect 4805 22815 5125 22816
rect 5165 22538 5231 22541
rect 5165 22536 6240 22538
rect 5165 22480 5170 22536
rect 5226 22480 6240 22536
rect 5165 22478 6240 22480
rect 5165 22475 5231 22478
rect 6180 22402 6240 22478
rect 7200 22402 8000 22432
rect 6180 22342 8000 22402
rect 1909 22336 2229 22337
rect 0 22266 800 22296
rect 1909 22272 1917 22336
rect 1981 22272 1997 22336
rect 2061 22272 2077 22336
rect 2141 22272 2157 22336
rect 2221 22272 2229 22336
rect 1909 22271 2229 22272
rect 3840 22336 4160 22337
rect 3840 22272 3848 22336
rect 3912 22272 3928 22336
rect 3992 22272 4008 22336
rect 4072 22272 4088 22336
rect 4152 22272 4160 22336
rect 3840 22271 4160 22272
rect 5770 22336 6090 22337
rect 5770 22272 5778 22336
rect 5842 22272 5858 22336
rect 5922 22272 5938 22336
rect 6002 22272 6018 22336
rect 6082 22272 6090 22336
rect 7200 22312 8000 22342
rect 5770 22271 6090 22272
rect 1577 22266 1643 22269
rect 0 22264 1643 22266
rect 0 22208 1582 22264
rect 1638 22208 1643 22264
rect 0 22206 1643 22208
rect 0 22176 800 22206
rect 1577 22203 1643 22206
rect 6177 21858 6243 21861
rect 7200 21858 8000 21888
rect 6177 21856 8000 21858
rect 6177 21800 6182 21856
rect 6238 21800 8000 21856
rect 6177 21798 8000 21800
rect 6177 21795 6243 21798
rect 2874 21792 3194 21793
rect 2874 21728 2882 21792
rect 2946 21728 2962 21792
rect 3026 21728 3042 21792
rect 3106 21728 3122 21792
rect 3186 21728 3194 21792
rect 2874 21727 3194 21728
rect 4805 21792 5125 21793
rect 4805 21728 4813 21792
rect 4877 21728 4893 21792
rect 4957 21728 4973 21792
rect 5037 21728 5053 21792
rect 5117 21728 5125 21792
rect 7200 21768 8000 21798
rect 4805 21727 5125 21728
rect 0 21586 800 21616
rect 1577 21586 1643 21589
rect 0 21584 1643 21586
rect 0 21528 1582 21584
rect 1638 21528 1643 21584
rect 0 21526 1643 21528
rect 0 21496 800 21526
rect 1577 21523 1643 21526
rect 1909 21248 2229 21249
rect 1909 21184 1917 21248
rect 1981 21184 1997 21248
rect 2061 21184 2077 21248
rect 2141 21184 2157 21248
rect 2221 21184 2229 21248
rect 1909 21183 2229 21184
rect 3840 21248 4160 21249
rect 3840 21184 3848 21248
rect 3912 21184 3928 21248
rect 3992 21184 4008 21248
rect 4072 21184 4088 21248
rect 4152 21184 4160 21248
rect 3840 21183 4160 21184
rect 5770 21248 6090 21249
rect 5770 21184 5778 21248
rect 5842 21184 5858 21248
rect 5922 21184 5938 21248
rect 6002 21184 6018 21248
rect 6082 21184 6090 21248
rect 5770 21183 6090 21184
rect 6177 21178 6243 21181
rect 7200 21178 8000 21208
rect 6177 21176 8000 21178
rect 6177 21120 6182 21176
rect 6238 21120 8000 21176
rect 6177 21118 8000 21120
rect 6177 21115 6243 21118
rect 7200 21088 8000 21118
rect 0 20770 800 20800
rect 1577 20770 1643 20773
rect 0 20768 1643 20770
rect 0 20712 1582 20768
rect 1638 20712 1643 20768
rect 0 20710 1643 20712
rect 0 20680 800 20710
rect 1577 20707 1643 20710
rect 2874 20704 3194 20705
rect 2874 20640 2882 20704
rect 2946 20640 2962 20704
rect 3026 20640 3042 20704
rect 3106 20640 3122 20704
rect 3186 20640 3194 20704
rect 2874 20639 3194 20640
rect 4805 20704 5125 20705
rect 4805 20640 4813 20704
rect 4877 20640 4893 20704
rect 4957 20640 4973 20704
rect 5037 20640 5053 20704
rect 5117 20640 5125 20704
rect 4805 20639 5125 20640
rect 6085 20634 6151 20637
rect 7200 20634 8000 20664
rect 6085 20632 8000 20634
rect 6085 20576 6090 20632
rect 6146 20576 8000 20632
rect 6085 20574 8000 20576
rect 6085 20571 6151 20574
rect 7200 20544 8000 20574
rect 1909 20160 2229 20161
rect 0 20090 800 20120
rect 1909 20096 1917 20160
rect 1981 20096 1997 20160
rect 2061 20096 2077 20160
rect 2141 20096 2157 20160
rect 2221 20096 2229 20160
rect 1909 20095 2229 20096
rect 3840 20160 4160 20161
rect 3840 20096 3848 20160
rect 3912 20096 3928 20160
rect 3992 20096 4008 20160
rect 4072 20096 4088 20160
rect 4152 20096 4160 20160
rect 3840 20095 4160 20096
rect 5770 20160 6090 20161
rect 5770 20096 5778 20160
rect 5842 20096 5858 20160
rect 5922 20096 5938 20160
rect 6002 20096 6018 20160
rect 6082 20096 6090 20160
rect 5770 20095 6090 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 800 20030
rect 1577 20027 1643 20030
rect 6177 20090 6243 20093
rect 7200 20090 8000 20120
rect 6177 20088 8000 20090
rect 6177 20032 6182 20088
rect 6238 20032 8000 20088
rect 6177 20030 8000 20032
rect 6177 20027 6243 20030
rect 7200 20000 8000 20030
rect 2874 19616 3194 19617
rect 2874 19552 2882 19616
rect 2946 19552 2962 19616
rect 3026 19552 3042 19616
rect 3106 19552 3122 19616
rect 3186 19552 3194 19616
rect 2874 19551 3194 19552
rect 4805 19616 5125 19617
rect 4805 19552 4813 19616
rect 4877 19552 4893 19616
rect 4957 19552 4973 19616
rect 5037 19552 5053 19616
rect 5117 19552 5125 19616
rect 4805 19551 5125 19552
rect 6085 19546 6151 19549
rect 7200 19546 8000 19576
rect 6085 19544 8000 19546
rect 6085 19488 6090 19544
rect 6146 19488 8000 19544
rect 6085 19486 8000 19488
rect 6085 19483 6151 19486
rect 7200 19456 8000 19486
rect 0 19274 800 19304
rect 1577 19274 1643 19277
rect 0 19272 1643 19274
rect 0 19216 1582 19272
rect 1638 19216 1643 19272
rect 0 19214 1643 19216
rect 0 19184 800 19214
rect 1577 19211 1643 19214
rect 1909 19072 2229 19073
rect 1909 19008 1917 19072
rect 1981 19008 1997 19072
rect 2061 19008 2077 19072
rect 2141 19008 2157 19072
rect 2221 19008 2229 19072
rect 1909 19007 2229 19008
rect 3840 19072 4160 19073
rect 3840 19008 3848 19072
rect 3912 19008 3928 19072
rect 3992 19008 4008 19072
rect 4072 19008 4088 19072
rect 4152 19008 4160 19072
rect 3840 19007 4160 19008
rect 5770 19072 6090 19073
rect 5770 19008 5778 19072
rect 5842 19008 5858 19072
rect 5922 19008 5938 19072
rect 6002 19008 6018 19072
rect 6082 19008 6090 19072
rect 5770 19007 6090 19008
rect 6453 19002 6519 19005
rect 7200 19002 8000 19032
rect 6453 19000 8000 19002
rect 6453 18944 6458 19000
rect 6514 18944 8000 19000
rect 6453 18942 8000 18944
rect 6453 18939 6519 18942
rect 7200 18912 8000 18942
rect 2874 18528 3194 18529
rect 0 18458 800 18488
rect 2874 18464 2882 18528
rect 2946 18464 2962 18528
rect 3026 18464 3042 18528
rect 3106 18464 3122 18528
rect 3186 18464 3194 18528
rect 2874 18463 3194 18464
rect 4805 18528 5125 18529
rect 4805 18464 4813 18528
rect 4877 18464 4893 18528
rect 4957 18464 4973 18528
rect 5037 18464 5053 18528
rect 5117 18464 5125 18528
rect 4805 18463 5125 18464
rect 1577 18458 1643 18461
rect 0 18456 1643 18458
rect 0 18400 1582 18456
rect 1638 18400 1643 18456
rect 0 18398 1643 18400
rect 0 18368 800 18398
rect 1577 18395 1643 18398
rect 6085 18458 6151 18461
rect 7200 18458 8000 18488
rect 6085 18456 8000 18458
rect 6085 18400 6090 18456
rect 6146 18400 8000 18456
rect 6085 18398 8000 18400
rect 6085 18395 6151 18398
rect 7200 18368 8000 18398
rect 1909 17984 2229 17985
rect 1909 17920 1917 17984
rect 1981 17920 1997 17984
rect 2061 17920 2077 17984
rect 2141 17920 2157 17984
rect 2221 17920 2229 17984
rect 1909 17919 2229 17920
rect 3840 17984 4160 17985
rect 3840 17920 3848 17984
rect 3912 17920 3928 17984
rect 3992 17920 4008 17984
rect 4072 17920 4088 17984
rect 4152 17920 4160 17984
rect 3840 17919 4160 17920
rect 5770 17984 6090 17985
rect 5770 17920 5778 17984
rect 5842 17920 5858 17984
rect 5922 17920 5938 17984
rect 6002 17920 6018 17984
rect 6082 17920 6090 17984
rect 5770 17919 6090 17920
rect 0 17778 800 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 800 17718
rect 1577 17715 1643 17718
rect 6177 17778 6243 17781
rect 7200 17778 8000 17808
rect 6177 17776 8000 17778
rect 6177 17720 6182 17776
rect 6238 17720 8000 17776
rect 6177 17718 8000 17720
rect 6177 17715 6243 17718
rect 7200 17688 8000 17718
rect 2874 17440 3194 17441
rect 2874 17376 2882 17440
rect 2946 17376 2962 17440
rect 3026 17376 3042 17440
rect 3106 17376 3122 17440
rect 3186 17376 3194 17440
rect 2874 17375 3194 17376
rect 4805 17440 5125 17441
rect 4805 17376 4813 17440
rect 4877 17376 4893 17440
rect 4957 17376 4973 17440
rect 5037 17376 5053 17440
rect 5117 17376 5125 17440
rect 4805 17375 5125 17376
rect 5441 17234 5507 17237
rect 7200 17234 8000 17264
rect 5441 17232 8000 17234
rect 5441 17176 5446 17232
rect 5502 17176 8000 17232
rect 5441 17174 8000 17176
rect 5441 17171 5507 17174
rect 7200 17144 8000 17174
rect 0 16962 800 16992
rect 1577 16962 1643 16965
rect 0 16960 1643 16962
rect 0 16904 1582 16960
rect 1638 16904 1643 16960
rect 0 16902 1643 16904
rect 0 16872 800 16902
rect 1577 16899 1643 16902
rect 1909 16896 2229 16897
rect 1909 16832 1917 16896
rect 1981 16832 1997 16896
rect 2061 16832 2077 16896
rect 2141 16832 2157 16896
rect 2221 16832 2229 16896
rect 1909 16831 2229 16832
rect 3840 16896 4160 16897
rect 3840 16832 3848 16896
rect 3912 16832 3928 16896
rect 3992 16832 4008 16896
rect 4072 16832 4088 16896
rect 4152 16832 4160 16896
rect 3840 16831 4160 16832
rect 5770 16896 6090 16897
rect 5770 16832 5778 16896
rect 5842 16832 5858 16896
rect 5922 16832 5938 16896
rect 6002 16832 6018 16896
rect 6082 16832 6090 16896
rect 5770 16831 6090 16832
rect 6177 16690 6243 16693
rect 7200 16690 8000 16720
rect 6177 16688 8000 16690
rect 6177 16632 6182 16688
rect 6238 16632 8000 16688
rect 6177 16630 8000 16632
rect 6177 16627 6243 16630
rect 7200 16600 8000 16630
rect 2874 16352 3194 16353
rect 0 16282 800 16312
rect 2874 16288 2882 16352
rect 2946 16288 2962 16352
rect 3026 16288 3042 16352
rect 3106 16288 3122 16352
rect 3186 16288 3194 16352
rect 2874 16287 3194 16288
rect 4805 16352 5125 16353
rect 4805 16288 4813 16352
rect 4877 16288 4893 16352
rect 4957 16288 4973 16352
rect 5037 16288 5053 16352
rect 5117 16288 5125 16352
rect 4805 16287 5125 16288
rect 1577 16282 1643 16285
rect 0 16280 1643 16282
rect 0 16224 1582 16280
rect 1638 16224 1643 16280
rect 0 16222 1643 16224
rect 0 16192 800 16222
rect 1577 16219 1643 16222
rect 6361 16146 6427 16149
rect 7200 16146 8000 16176
rect 6361 16144 8000 16146
rect 6361 16088 6366 16144
rect 6422 16088 8000 16144
rect 6361 16086 8000 16088
rect 6361 16083 6427 16086
rect 7200 16056 8000 16086
rect 1909 15808 2229 15809
rect 1909 15744 1917 15808
rect 1981 15744 1997 15808
rect 2061 15744 2077 15808
rect 2141 15744 2157 15808
rect 2221 15744 2229 15808
rect 1909 15743 2229 15744
rect 3840 15808 4160 15809
rect 3840 15744 3848 15808
rect 3912 15744 3928 15808
rect 3992 15744 4008 15808
rect 4072 15744 4088 15808
rect 4152 15744 4160 15808
rect 3840 15743 4160 15744
rect 5770 15808 6090 15809
rect 5770 15744 5778 15808
rect 5842 15744 5858 15808
rect 5922 15744 5938 15808
rect 6002 15744 6018 15808
rect 6082 15744 6090 15808
rect 5770 15743 6090 15744
rect 6177 15602 6243 15605
rect 7200 15602 8000 15632
rect 6177 15600 8000 15602
rect 6177 15544 6182 15600
rect 6238 15544 8000 15600
rect 6177 15542 8000 15544
rect 6177 15539 6243 15542
rect 7200 15512 8000 15542
rect 0 15466 800 15496
rect 1577 15466 1643 15469
rect 0 15464 1643 15466
rect 0 15408 1582 15464
rect 1638 15408 1643 15464
rect 0 15406 1643 15408
rect 0 15376 800 15406
rect 1577 15403 1643 15406
rect 2874 15264 3194 15265
rect 2874 15200 2882 15264
rect 2946 15200 2962 15264
rect 3026 15200 3042 15264
rect 3106 15200 3122 15264
rect 3186 15200 3194 15264
rect 2874 15199 3194 15200
rect 4805 15264 5125 15265
rect 4805 15200 4813 15264
rect 4877 15200 4893 15264
rect 4957 15200 4973 15264
rect 5037 15200 5053 15264
rect 5117 15200 5125 15264
rect 4805 15199 5125 15200
rect 5441 15058 5507 15061
rect 7200 15058 8000 15088
rect 5441 15056 8000 15058
rect 5441 15000 5446 15056
rect 5502 15000 8000 15056
rect 5441 14998 8000 15000
rect 5441 14995 5507 14998
rect 7200 14968 8000 14998
rect 0 14786 800 14816
rect 1577 14786 1643 14789
rect 0 14784 1643 14786
rect 0 14728 1582 14784
rect 1638 14728 1643 14784
rect 0 14726 1643 14728
rect 0 14696 800 14726
rect 1577 14723 1643 14726
rect 1909 14720 2229 14721
rect 1909 14656 1917 14720
rect 1981 14656 1997 14720
rect 2061 14656 2077 14720
rect 2141 14656 2157 14720
rect 2221 14656 2229 14720
rect 1909 14655 2229 14656
rect 3840 14720 4160 14721
rect 3840 14656 3848 14720
rect 3912 14656 3928 14720
rect 3992 14656 4008 14720
rect 4072 14656 4088 14720
rect 4152 14656 4160 14720
rect 3840 14655 4160 14656
rect 5770 14720 6090 14721
rect 5770 14656 5778 14720
rect 5842 14656 5858 14720
rect 5922 14656 5938 14720
rect 6002 14656 6018 14720
rect 6082 14656 6090 14720
rect 5770 14655 6090 14656
rect 6177 14514 6243 14517
rect 7200 14514 8000 14544
rect 6177 14512 8000 14514
rect 6177 14456 6182 14512
rect 6238 14456 8000 14512
rect 6177 14454 8000 14456
rect 6177 14451 6243 14454
rect 7200 14424 8000 14454
rect 2874 14176 3194 14177
rect 2874 14112 2882 14176
rect 2946 14112 2962 14176
rect 3026 14112 3042 14176
rect 3106 14112 3122 14176
rect 3186 14112 3194 14176
rect 2874 14111 3194 14112
rect 4805 14176 5125 14177
rect 4805 14112 4813 14176
rect 4877 14112 4893 14176
rect 4957 14112 4973 14176
rect 5037 14112 5053 14176
rect 5117 14112 5125 14176
rect 4805 14111 5125 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 5809 13834 5875 13837
rect 7200 13834 8000 13864
rect 5809 13832 8000 13834
rect 5809 13776 5814 13832
rect 5870 13776 8000 13832
rect 5809 13774 8000 13776
rect 5809 13771 5875 13774
rect 7200 13744 8000 13774
rect 1909 13632 2229 13633
rect 1909 13568 1917 13632
rect 1981 13568 1997 13632
rect 2061 13568 2077 13632
rect 2141 13568 2157 13632
rect 2221 13568 2229 13632
rect 1909 13567 2229 13568
rect 3840 13632 4160 13633
rect 3840 13568 3848 13632
rect 3912 13568 3928 13632
rect 3992 13568 4008 13632
rect 4072 13568 4088 13632
rect 4152 13568 4160 13632
rect 3840 13567 4160 13568
rect 5770 13632 6090 13633
rect 5770 13568 5778 13632
rect 5842 13568 5858 13632
rect 5922 13568 5938 13632
rect 6002 13568 6018 13632
rect 6082 13568 6090 13632
rect 5770 13567 6090 13568
rect 6085 13290 6151 13293
rect 7200 13290 8000 13320
rect 6085 13288 8000 13290
rect 6085 13232 6090 13288
rect 6146 13232 8000 13288
rect 6085 13230 8000 13232
rect 6085 13227 6151 13230
rect 7200 13200 8000 13230
rect 0 13154 800 13184
rect 1577 13154 1643 13157
rect 0 13152 1643 13154
rect 0 13096 1582 13152
rect 1638 13096 1643 13152
rect 0 13094 1643 13096
rect 0 13064 800 13094
rect 1577 13091 1643 13094
rect 2874 13088 3194 13089
rect 2874 13024 2882 13088
rect 2946 13024 2962 13088
rect 3026 13024 3042 13088
rect 3106 13024 3122 13088
rect 3186 13024 3194 13088
rect 2874 13023 3194 13024
rect 4805 13088 5125 13089
rect 4805 13024 4813 13088
rect 4877 13024 4893 13088
rect 4957 13024 4973 13088
rect 5037 13024 5053 13088
rect 5117 13024 5125 13088
rect 4805 13023 5125 13024
rect 5809 12746 5875 12749
rect 7200 12746 8000 12776
rect 5809 12744 8000 12746
rect 5809 12688 5814 12744
rect 5870 12688 8000 12744
rect 5809 12686 8000 12688
rect 5809 12683 5875 12686
rect 7200 12656 8000 12686
rect 1909 12544 2229 12545
rect 0 12474 800 12504
rect 1909 12480 1917 12544
rect 1981 12480 1997 12544
rect 2061 12480 2077 12544
rect 2141 12480 2157 12544
rect 2221 12480 2229 12544
rect 1909 12479 2229 12480
rect 3840 12544 4160 12545
rect 3840 12480 3848 12544
rect 3912 12480 3928 12544
rect 3992 12480 4008 12544
rect 4072 12480 4088 12544
rect 4152 12480 4160 12544
rect 3840 12479 4160 12480
rect 5770 12544 6090 12545
rect 5770 12480 5778 12544
rect 5842 12480 5858 12544
rect 5922 12480 5938 12544
rect 6002 12480 6018 12544
rect 6082 12480 6090 12544
rect 5770 12479 6090 12480
rect 1577 12474 1643 12477
rect 0 12472 1643 12474
rect 0 12416 1582 12472
rect 1638 12416 1643 12472
rect 0 12414 1643 12416
rect 0 12384 800 12414
rect 1577 12411 1643 12414
rect 6085 12202 6151 12205
rect 7200 12202 8000 12232
rect 6085 12200 8000 12202
rect 6085 12144 6090 12200
rect 6146 12144 8000 12200
rect 6085 12142 8000 12144
rect 6085 12139 6151 12142
rect 7200 12112 8000 12142
rect 2874 12000 3194 12001
rect 2874 11936 2882 12000
rect 2946 11936 2962 12000
rect 3026 11936 3042 12000
rect 3106 11936 3122 12000
rect 3186 11936 3194 12000
rect 2874 11935 3194 11936
rect 4805 12000 5125 12001
rect 4805 11936 4813 12000
rect 4877 11936 4893 12000
rect 4957 11936 4973 12000
rect 5037 11936 5053 12000
rect 5117 11936 5125 12000
rect 4805 11935 5125 11936
rect 0 11658 800 11688
rect 1577 11658 1643 11661
rect 0 11656 1643 11658
rect 0 11600 1582 11656
rect 1638 11600 1643 11656
rect 0 11598 1643 11600
rect 0 11568 800 11598
rect 1577 11595 1643 11598
rect 6177 11658 6243 11661
rect 7200 11658 8000 11688
rect 6177 11656 8000 11658
rect 6177 11600 6182 11656
rect 6238 11600 8000 11656
rect 6177 11598 8000 11600
rect 6177 11595 6243 11598
rect 7200 11568 8000 11598
rect 1909 11456 2229 11457
rect 1909 11392 1917 11456
rect 1981 11392 1997 11456
rect 2061 11392 2077 11456
rect 2141 11392 2157 11456
rect 2221 11392 2229 11456
rect 1909 11391 2229 11392
rect 3840 11456 4160 11457
rect 3840 11392 3848 11456
rect 3912 11392 3928 11456
rect 3992 11392 4008 11456
rect 4072 11392 4088 11456
rect 4152 11392 4160 11456
rect 3840 11391 4160 11392
rect 5770 11456 6090 11457
rect 5770 11392 5778 11456
rect 5842 11392 5858 11456
rect 5922 11392 5938 11456
rect 6002 11392 6018 11456
rect 6082 11392 6090 11456
rect 5770 11391 6090 11392
rect 4797 11114 4863 11117
rect 7200 11114 8000 11144
rect 4797 11112 8000 11114
rect 4797 11056 4802 11112
rect 4858 11056 8000 11112
rect 4797 11054 8000 11056
rect 4797 11051 4863 11054
rect 7200 11024 8000 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 2874 10912 3194 10913
rect 2874 10848 2882 10912
rect 2946 10848 2962 10912
rect 3026 10848 3042 10912
rect 3106 10848 3122 10912
rect 3186 10848 3194 10912
rect 2874 10847 3194 10848
rect 4805 10912 5125 10913
rect 4805 10848 4813 10912
rect 4877 10848 4893 10912
rect 4957 10848 4973 10912
rect 5037 10848 5053 10912
rect 5117 10848 5125 10912
rect 4805 10847 5125 10848
rect 5349 10570 5415 10573
rect 5349 10568 6240 10570
rect 5349 10512 5354 10568
rect 5410 10512 6240 10568
rect 5349 10510 6240 10512
rect 5349 10507 5415 10510
rect 6180 10434 6240 10510
rect 7200 10434 8000 10464
rect 6180 10374 8000 10434
rect 1909 10368 2229 10369
rect 1909 10304 1917 10368
rect 1981 10304 1997 10368
rect 2061 10304 2077 10368
rect 2141 10304 2157 10368
rect 2221 10304 2229 10368
rect 1909 10303 2229 10304
rect 3840 10368 4160 10369
rect 3840 10304 3848 10368
rect 3912 10304 3928 10368
rect 3992 10304 4008 10368
rect 4072 10304 4088 10368
rect 4152 10304 4160 10368
rect 3840 10303 4160 10304
rect 5770 10368 6090 10369
rect 5770 10304 5778 10368
rect 5842 10304 5858 10368
rect 5922 10304 5938 10368
rect 6002 10304 6018 10368
rect 6082 10304 6090 10368
rect 7200 10344 8000 10374
rect 5770 10303 6090 10304
rect 0 10162 800 10192
rect 1577 10162 1643 10165
rect 0 10160 1643 10162
rect 0 10104 1582 10160
rect 1638 10104 1643 10160
rect 0 10102 1643 10104
rect 0 10072 800 10102
rect 1577 10099 1643 10102
rect 5441 9890 5507 9893
rect 7200 9890 8000 9920
rect 5441 9888 8000 9890
rect 5441 9832 5446 9888
rect 5502 9832 8000 9888
rect 5441 9830 8000 9832
rect 5441 9827 5507 9830
rect 2874 9824 3194 9825
rect 2874 9760 2882 9824
rect 2946 9760 2962 9824
rect 3026 9760 3042 9824
rect 3106 9760 3122 9824
rect 3186 9760 3194 9824
rect 2874 9759 3194 9760
rect 4805 9824 5125 9825
rect 4805 9760 4813 9824
rect 4877 9760 4893 9824
rect 4957 9760 4973 9824
rect 5037 9760 5053 9824
rect 5117 9760 5125 9824
rect 7200 9800 8000 9830
rect 4805 9759 5125 9760
rect 5165 9482 5231 9485
rect 5165 9480 6240 9482
rect 5165 9424 5170 9480
rect 5226 9424 6240 9480
rect 5165 9422 6240 9424
rect 5165 9419 5231 9422
rect 0 9346 800 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 6180 9346 6240 9422
rect 7200 9346 8000 9376
rect 6180 9286 8000 9346
rect 0 9256 800 9286
rect 1577 9283 1643 9286
rect 1909 9280 2229 9281
rect 1909 9216 1917 9280
rect 1981 9216 1997 9280
rect 2061 9216 2077 9280
rect 2141 9216 2157 9280
rect 2221 9216 2229 9280
rect 1909 9215 2229 9216
rect 3840 9280 4160 9281
rect 3840 9216 3848 9280
rect 3912 9216 3928 9280
rect 3992 9216 4008 9280
rect 4072 9216 4088 9280
rect 4152 9216 4160 9280
rect 3840 9215 4160 9216
rect 5770 9280 6090 9281
rect 5770 9216 5778 9280
rect 5842 9216 5858 9280
rect 5922 9216 5938 9280
rect 6002 9216 6018 9280
rect 6082 9216 6090 9280
rect 7200 9256 8000 9286
rect 5770 9215 6090 9216
rect 6913 8802 6979 8805
rect 7200 8802 8000 8832
rect 6913 8800 8000 8802
rect 6913 8744 6918 8800
rect 6974 8744 8000 8800
rect 6913 8742 8000 8744
rect 6913 8739 6979 8742
rect 2874 8736 3194 8737
rect 0 8666 800 8696
rect 2874 8672 2882 8736
rect 2946 8672 2962 8736
rect 3026 8672 3042 8736
rect 3106 8672 3122 8736
rect 3186 8672 3194 8736
rect 2874 8671 3194 8672
rect 4805 8736 5125 8737
rect 4805 8672 4813 8736
rect 4877 8672 4893 8736
rect 4957 8672 4973 8736
rect 5037 8672 5053 8736
rect 5117 8672 5125 8736
rect 7200 8712 8000 8742
rect 4805 8671 5125 8672
rect 1577 8666 1643 8669
rect 0 8664 1643 8666
rect 0 8608 1582 8664
rect 1638 8608 1643 8664
rect 0 8606 1643 8608
rect 0 8576 800 8606
rect 1577 8603 1643 8606
rect 5441 8394 5507 8397
rect 5441 8392 6240 8394
rect 5441 8336 5446 8392
rect 5502 8336 6240 8392
rect 5441 8334 6240 8336
rect 5441 8331 5507 8334
rect 6180 8258 6240 8334
rect 7200 8258 8000 8288
rect 6180 8198 8000 8258
rect 1909 8192 2229 8193
rect 1909 8128 1917 8192
rect 1981 8128 1997 8192
rect 2061 8128 2077 8192
rect 2141 8128 2157 8192
rect 2221 8128 2229 8192
rect 1909 8127 2229 8128
rect 3840 8192 4160 8193
rect 3840 8128 3848 8192
rect 3912 8128 3928 8192
rect 3992 8128 4008 8192
rect 4072 8128 4088 8192
rect 4152 8128 4160 8192
rect 3840 8127 4160 8128
rect 5770 8192 6090 8193
rect 5770 8128 5778 8192
rect 5842 8128 5858 8192
rect 5922 8128 5938 8192
rect 6002 8128 6018 8192
rect 6082 8128 6090 8192
rect 7200 8168 8000 8198
rect 5770 8127 6090 8128
rect 0 7850 800 7880
rect 1577 7850 1643 7853
rect 0 7848 1643 7850
rect 0 7792 1582 7848
rect 1638 7792 1643 7848
rect 0 7790 1643 7792
rect 0 7760 800 7790
rect 1577 7787 1643 7790
rect 5349 7714 5415 7717
rect 7200 7714 8000 7744
rect 5349 7712 8000 7714
rect 5349 7656 5354 7712
rect 5410 7656 8000 7712
rect 5349 7654 8000 7656
rect 5349 7651 5415 7654
rect 2874 7648 3194 7649
rect 2874 7584 2882 7648
rect 2946 7584 2962 7648
rect 3026 7584 3042 7648
rect 3106 7584 3122 7648
rect 3186 7584 3194 7648
rect 2874 7583 3194 7584
rect 4805 7648 5125 7649
rect 4805 7584 4813 7648
rect 4877 7584 4893 7648
rect 4957 7584 4973 7648
rect 5037 7584 5053 7648
rect 5117 7584 5125 7648
rect 7200 7624 8000 7654
rect 4805 7583 5125 7584
rect 0 7170 800 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 800 7110
rect 1577 7107 1643 7110
rect 1909 7104 2229 7105
rect 1909 7040 1917 7104
rect 1981 7040 1997 7104
rect 2061 7040 2077 7104
rect 2141 7040 2157 7104
rect 2221 7040 2229 7104
rect 1909 7039 2229 7040
rect 3840 7104 4160 7105
rect 3840 7040 3848 7104
rect 3912 7040 3928 7104
rect 3992 7040 4008 7104
rect 4072 7040 4088 7104
rect 4152 7040 4160 7104
rect 3840 7039 4160 7040
rect 5770 7104 6090 7105
rect 5770 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5938 7104
rect 6002 7040 6018 7104
rect 6082 7040 6090 7104
rect 5770 7039 6090 7040
rect 7005 7034 7071 7037
rect 7200 7034 8000 7064
rect 7005 7032 8000 7034
rect 7005 6976 7010 7032
rect 7066 6976 8000 7032
rect 7005 6974 8000 6976
rect 7005 6971 7071 6974
rect 7200 6944 8000 6974
rect 2874 6560 3194 6561
rect 2874 6496 2882 6560
rect 2946 6496 2962 6560
rect 3026 6496 3042 6560
rect 3106 6496 3122 6560
rect 3186 6496 3194 6560
rect 2874 6495 3194 6496
rect 4805 6560 5125 6561
rect 4805 6496 4813 6560
rect 4877 6496 4893 6560
rect 4957 6496 4973 6560
rect 5037 6496 5053 6560
rect 5117 6496 5125 6560
rect 4805 6495 5125 6496
rect 5257 6490 5323 6493
rect 7200 6490 8000 6520
rect 5257 6488 8000 6490
rect 5257 6432 5262 6488
rect 5318 6432 8000 6488
rect 5257 6430 8000 6432
rect 5257 6427 5323 6430
rect 7200 6400 8000 6430
rect 0 6354 800 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 800 6294
rect 1577 6291 1643 6294
rect 1909 6016 2229 6017
rect 1909 5952 1917 6016
rect 1981 5952 1997 6016
rect 2061 5952 2077 6016
rect 2141 5952 2157 6016
rect 2221 5952 2229 6016
rect 1909 5951 2229 5952
rect 3840 6016 4160 6017
rect 3840 5952 3848 6016
rect 3912 5952 3928 6016
rect 3992 5952 4008 6016
rect 4072 5952 4088 6016
rect 4152 5952 4160 6016
rect 3840 5951 4160 5952
rect 5770 6016 6090 6017
rect 5770 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6018 6016
rect 6082 5952 6090 6016
rect 5770 5951 6090 5952
rect 7005 5946 7071 5949
rect 7200 5946 8000 5976
rect 7005 5944 8000 5946
rect 7005 5888 7010 5944
rect 7066 5888 8000 5944
rect 7005 5886 8000 5888
rect 7005 5883 7071 5886
rect 7200 5856 8000 5886
rect 0 5674 800 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 800 5614
rect 1577 5611 1643 5614
rect 2874 5472 3194 5473
rect 2874 5408 2882 5472
rect 2946 5408 2962 5472
rect 3026 5408 3042 5472
rect 3106 5408 3122 5472
rect 3186 5408 3194 5472
rect 2874 5407 3194 5408
rect 4805 5472 5125 5473
rect 4805 5408 4813 5472
rect 4877 5408 4893 5472
rect 4957 5408 4973 5472
rect 5037 5408 5053 5472
rect 5117 5408 5125 5472
rect 4805 5407 5125 5408
rect 7200 5402 8000 5432
rect 5214 5342 8000 5402
rect 3601 5266 3667 5269
rect 5214 5266 5274 5342
rect 7200 5312 8000 5342
rect 3601 5264 5274 5266
rect 3601 5208 3606 5264
rect 3662 5208 5274 5264
rect 3601 5206 5274 5208
rect 3601 5203 3667 5206
rect 5441 5130 5507 5133
rect 5441 5128 6378 5130
rect 5441 5072 5446 5128
rect 5502 5072 6378 5128
rect 5441 5070 6378 5072
rect 5441 5067 5507 5070
rect 1909 4928 2229 4929
rect 0 4858 800 4888
rect 1909 4864 1917 4928
rect 1981 4864 1997 4928
rect 2061 4864 2077 4928
rect 2141 4864 2157 4928
rect 2221 4864 2229 4928
rect 1909 4863 2229 4864
rect 3840 4928 4160 4929
rect 3840 4864 3848 4928
rect 3912 4864 3928 4928
rect 3992 4864 4008 4928
rect 4072 4864 4088 4928
rect 4152 4864 4160 4928
rect 3840 4863 4160 4864
rect 5770 4928 6090 4929
rect 5770 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6018 4928
rect 6082 4864 6090 4928
rect 5770 4863 6090 4864
rect 1577 4858 1643 4861
rect 0 4856 1643 4858
rect 0 4800 1582 4856
rect 1638 4800 1643 4856
rect 0 4798 1643 4800
rect 6318 4858 6378 5070
rect 7200 4858 8000 4888
rect 6318 4798 8000 4858
rect 0 4768 800 4798
rect 1577 4795 1643 4798
rect 7200 4768 8000 4798
rect 2874 4384 3194 4385
rect 2874 4320 2882 4384
rect 2946 4320 2962 4384
rect 3026 4320 3042 4384
rect 3106 4320 3122 4384
rect 3186 4320 3194 4384
rect 2874 4319 3194 4320
rect 4805 4384 5125 4385
rect 4805 4320 4813 4384
rect 4877 4320 4893 4384
rect 4957 4320 4973 4384
rect 5037 4320 5053 4384
rect 5117 4320 5125 4384
rect 4805 4319 5125 4320
rect 5257 4314 5323 4317
rect 7200 4314 8000 4344
rect 5257 4312 8000 4314
rect 5257 4256 5262 4312
rect 5318 4256 8000 4312
rect 5257 4254 8000 4256
rect 5257 4251 5323 4254
rect 7200 4224 8000 4254
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 1909 3840 2229 3841
rect 1909 3776 1917 3840
rect 1981 3776 1997 3840
rect 2061 3776 2077 3840
rect 2141 3776 2157 3840
rect 2221 3776 2229 3840
rect 1909 3775 2229 3776
rect 3840 3840 4160 3841
rect 3840 3776 3848 3840
rect 3912 3776 3928 3840
rect 3992 3776 4008 3840
rect 4072 3776 4088 3840
rect 4152 3776 4160 3840
rect 3840 3775 4160 3776
rect 5770 3840 6090 3841
rect 5770 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6018 3840
rect 6082 3776 6090 3840
rect 5770 3775 6090 3776
rect 4521 3634 4587 3637
rect 7200 3634 8000 3664
rect 4521 3632 8000 3634
rect 4521 3576 4526 3632
rect 4582 3576 8000 3632
rect 4521 3574 8000 3576
rect 4521 3571 4587 3574
rect 7200 3544 8000 3574
rect 0 3362 800 3392
rect 1577 3362 1643 3365
rect 0 3360 1643 3362
rect 0 3304 1582 3360
rect 1638 3304 1643 3360
rect 0 3302 1643 3304
rect 0 3272 800 3302
rect 1577 3299 1643 3302
rect 2874 3296 3194 3297
rect 2874 3232 2882 3296
rect 2946 3232 2962 3296
rect 3026 3232 3042 3296
rect 3106 3232 3122 3296
rect 3186 3232 3194 3296
rect 2874 3231 3194 3232
rect 4805 3296 5125 3297
rect 4805 3232 4813 3296
rect 4877 3232 4893 3296
rect 4957 3232 4973 3296
rect 5037 3232 5053 3296
rect 5117 3232 5125 3296
rect 4805 3231 5125 3232
rect 5993 3090 6059 3093
rect 7200 3090 8000 3120
rect 5993 3088 8000 3090
rect 5993 3032 5998 3088
rect 6054 3032 8000 3088
rect 5993 3030 8000 3032
rect 5993 3027 6059 3030
rect 7200 3000 8000 3030
rect 1909 2752 2229 2753
rect 1909 2688 1917 2752
rect 1981 2688 1997 2752
rect 2061 2688 2077 2752
rect 2141 2688 2157 2752
rect 2221 2688 2229 2752
rect 1909 2687 2229 2688
rect 3840 2752 4160 2753
rect 3840 2688 3848 2752
rect 3912 2688 3928 2752
rect 3992 2688 4008 2752
rect 4072 2688 4088 2752
rect 4152 2688 4160 2752
rect 3840 2687 4160 2688
rect 5770 2752 6090 2753
rect 5770 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5938 2752
rect 6002 2688 6018 2752
rect 6082 2688 6090 2752
rect 5770 2687 6090 2688
rect 0 2546 800 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 0 2456 800 2486
rect 1393 2483 1459 2486
rect 5165 2546 5231 2549
rect 7200 2546 8000 2576
rect 5165 2544 8000 2546
rect 5165 2488 5170 2544
rect 5226 2488 8000 2544
rect 5165 2486 8000 2488
rect 5165 2483 5231 2486
rect 7200 2456 8000 2486
rect 2874 2208 3194 2209
rect 2874 2144 2882 2208
rect 2946 2144 2962 2208
rect 3026 2144 3042 2208
rect 3106 2144 3122 2208
rect 3186 2144 3194 2208
rect 2874 2143 3194 2144
rect 4805 2208 5125 2209
rect 4805 2144 4813 2208
rect 4877 2144 4893 2208
rect 4957 2144 4973 2208
rect 5037 2144 5053 2208
rect 5117 2144 5125 2208
rect 4805 2143 5125 2144
rect 6177 2002 6243 2005
rect 7200 2002 8000 2032
rect 6177 2000 8000 2002
rect 6177 1944 6182 2000
rect 6238 1944 8000 2000
rect 6177 1942 8000 1944
rect 6177 1939 6243 1942
rect 7200 1912 8000 1942
rect 0 1866 800 1896
rect 1485 1866 1551 1869
rect 0 1864 1551 1866
rect 0 1808 1490 1864
rect 1546 1808 1551 1864
rect 0 1806 1551 1808
rect 0 1776 800 1806
rect 1485 1803 1551 1806
rect 5165 1458 5231 1461
rect 7200 1458 8000 1488
rect 5165 1456 8000 1458
rect 5165 1400 5170 1456
rect 5226 1400 8000 1456
rect 5165 1398 8000 1400
rect 5165 1395 5231 1398
rect 7200 1368 8000 1398
rect 0 1050 800 1080
rect 1577 1050 1643 1053
rect 0 1048 1643 1050
rect 0 992 1582 1048
rect 1638 992 1643 1048
rect 0 990 1643 992
rect 0 960 800 990
rect 1577 987 1643 990
rect 5809 914 5875 917
rect 7200 914 8000 944
rect 5809 912 8000 914
rect 5809 856 5814 912
rect 5870 856 8000 912
rect 5809 854 8000 856
rect 5809 851 5875 854
rect 7200 824 8000 854
rect 0 370 800 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 800 310
rect 2773 307 2839 310
rect 4245 370 4311 373
rect 7200 370 8000 400
rect 4245 368 8000 370
rect 4245 312 4250 368
rect 4306 312 8000 368
rect 4245 310 8000 312
rect 4245 307 4311 310
rect 7200 280 8000 310
<< via3 >>
rect 2882 57692 2946 57696
rect 2882 57636 2886 57692
rect 2886 57636 2942 57692
rect 2942 57636 2946 57692
rect 2882 57632 2946 57636
rect 2962 57692 3026 57696
rect 2962 57636 2966 57692
rect 2966 57636 3022 57692
rect 3022 57636 3026 57692
rect 2962 57632 3026 57636
rect 3042 57692 3106 57696
rect 3042 57636 3046 57692
rect 3046 57636 3102 57692
rect 3102 57636 3106 57692
rect 3042 57632 3106 57636
rect 3122 57692 3186 57696
rect 3122 57636 3126 57692
rect 3126 57636 3182 57692
rect 3182 57636 3186 57692
rect 3122 57632 3186 57636
rect 4813 57692 4877 57696
rect 4813 57636 4817 57692
rect 4817 57636 4873 57692
rect 4873 57636 4877 57692
rect 4813 57632 4877 57636
rect 4893 57692 4957 57696
rect 4893 57636 4897 57692
rect 4897 57636 4953 57692
rect 4953 57636 4957 57692
rect 4893 57632 4957 57636
rect 4973 57692 5037 57696
rect 4973 57636 4977 57692
rect 4977 57636 5033 57692
rect 5033 57636 5037 57692
rect 4973 57632 5037 57636
rect 5053 57692 5117 57696
rect 5053 57636 5057 57692
rect 5057 57636 5113 57692
rect 5113 57636 5117 57692
rect 5053 57632 5117 57636
rect 1917 57148 1981 57152
rect 1917 57092 1921 57148
rect 1921 57092 1977 57148
rect 1977 57092 1981 57148
rect 1917 57088 1981 57092
rect 1997 57148 2061 57152
rect 1997 57092 2001 57148
rect 2001 57092 2057 57148
rect 2057 57092 2061 57148
rect 1997 57088 2061 57092
rect 2077 57148 2141 57152
rect 2077 57092 2081 57148
rect 2081 57092 2137 57148
rect 2137 57092 2141 57148
rect 2077 57088 2141 57092
rect 2157 57148 2221 57152
rect 2157 57092 2161 57148
rect 2161 57092 2217 57148
rect 2217 57092 2221 57148
rect 2157 57088 2221 57092
rect 3848 57148 3912 57152
rect 3848 57092 3852 57148
rect 3852 57092 3908 57148
rect 3908 57092 3912 57148
rect 3848 57088 3912 57092
rect 3928 57148 3992 57152
rect 3928 57092 3932 57148
rect 3932 57092 3988 57148
rect 3988 57092 3992 57148
rect 3928 57088 3992 57092
rect 4008 57148 4072 57152
rect 4008 57092 4012 57148
rect 4012 57092 4068 57148
rect 4068 57092 4072 57148
rect 4008 57088 4072 57092
rect 4088 57148 4152 57152
rect 4088 57092 4092 57148
rect 4092 57092 4148 57148
rect 4148 57092 4152 57148
rect 4088 57088 4152 57092
rect 5778 57148 5842 57152
rect 5778 57092 5782 57148
rect 5782 57092 5838 57148
rect 5838 57092 5842 57148
rect 5778 57088 5842 57092
rect 5858 57148 5922 57152
rect 5858 57092 5862 57148
rect 5862 57092 5918 57148
rect 5918 57092 5922 57148
rect 5858 57088 5922 57092
rect 5938 57148 6002 57152
rect 5938 57092 5942 57148
rect 5942 57092 5998 57148
rect 5998 57092 6002 57148
rect 5938 57088 6002 57092
rect 6018 57148 6082 57152
rect 6018 57092 6022 57148
rect 6022 57092 6078 57148
rect 6078 57092 6082 57148
rect 6018 57088 6082 57092
rect 2882 56604 2946 56608
rect 2882 56548 2886 56604
rect 2886 56548 2942 56604
rect 2942 56548 2946 56604
rect 2882 56544 2946 56548
rect 2962 56604 3026 56608
rect 2962 56548 2966 56604
rect 2966 56548 3022 56604
rect 3022 56548 3026 56604
rect 2962 56544 3026 56548
rect 3042 56604 3106 56608
rect 3042 56548 3046 56604
rect 3046 56548 3102 56604
rect 3102 56548 3106 56604
rect 3042 56544 3106 56548
rect 3122 56604 3186 56608
rect 3122 56548 3126 56604
rect 3126 56548 3182 56604
rect 3182 56548 3186 56604
rect 3122 56544 3186 56548
rect 4813 56604 4877 56608
rect 4813 56548 4817 56604
rect 4817 56548 4873 56604
rect 4873 56548 4877 56604
rect 4813 56544 4877 56548
rect 4893 56604 4957 56608
rect 4893 56548 4897 56604
rect 4897 56548 4953 56604
rect 4953 56548 4957 56604
rect 4893 56544 4957 56548
rect 4973 56604 5037 56608
rect 4973 56548 4977 56604
rect 4977 56548 5033 56604
rect 5033 56548 5037 56604
rect 4973 56544 5037 56548
rect 5053 56604 5117 56608
rect 5053 56548 5057 56604
rect 5057 56548 5113 56604
rect 5113 56548 5117 56604
rect 5053 56544 5117 56548
rect 1917 56060 1981 56064
rect 1917 56004 1921 56060
rect 1921 56004 1977 56060
rect 1977 56004 1981 56060
rect 1917 56000 1981 56004
rect 1997 56060 2061 56064
rect 1997 56004 2001 56060
rect 2001 56004 2057 56060
rect 2057 56004 2061 56060
rect 1997 56000 2061 56004
rect 2077 56060 2141 56064
rect 2077 56004 2081 56060
rect 2081 56004 2137 56060
rect 2137 56004 2141 56060
rect 2077 56000 2141 56004
rect 2157 56060 2221 56064
rect 2157 56004 2161 56060
rect 2161 56004 2217 56060
rect 2217 56004 2221 56060
rect 2157 56000 2221 56004
rect 3848 56060 3912 56064
rect 3848 56004 3852 56060
rect 3852 56004 3908 56060
rect 3908 56004 3912 56060
rect 3848 56000 3912 56004
rect 3928 56060 3992 56064
rect 3928 56004 3932 56060
rect 3932 56004 3988 56060
rect 3988 56004 3992 56060
rect 3928 56000 3992 56004
rect 4008 56060 4072 56064
rect 4008 56004 4012 56060
rect 4012 56004 4068 56060
rect 4068 56004 4072 56060
rect 4008 56000 4072 56004
rect 4088 56060 4152 56064
rect 4088 56004 4092 56060
rect 4092 56004 4148 56060
rect 4148 56004 4152 56060
rect 4088 56000 4152 56004
rect 5778 56060 5842 56064
rect 5778 56004 5782 56060
rect 5782 56004 5838 56060
rect 5838 56004 5842 56060
rect 5778 56000 5842 56004
rect 5858 56060 5922 56064
rect 5858 56004 5862 56060
rect 5862 56004 5918 56060
rect 5918 56004 5922 56060
rect 5858 56000 5922 56004
rect 5938 56060 6002 56064
rect 5938 56004 5942 56060
rect 5942 56004 5998 56060
rect 5998 56004 6002 56060
rect 5938 56000 6002 56004
rect 6018 56060 6082 56064
rect 6018 56004 6022 56060
rect 6022 56004 6078 56060
rect 6078 56004 6082 56060
rect 6018 56000 6082 56004
rect 2882 55516 2946 55520
rect 2882 55460 2886 55516
rect 2886 55460 2942 55516
rect 2942 55460 2946 55516
rect 2882 55456 2946 55460
rect 2962 55516 3026 55520
rect 2962 55460 2966 55516
rect 2966 55460 3022 55516
rect 3022 55460 3026 55516
rect 2962 55456 3026 55460
rect 3042 55516 3106 55520
rect 3042 55460 3046 55516
rect 3046 55460 3102 55516
rect 3102 55460 3106 55516
rect 3042 55456 3106 55460
rect 3122 55516 3186 55520
rect 3122 55460 3126 55516
rect 3126 55460 3182 55516
rect 3182 55460 3186 55516
rect 3122 55456 3186 55460
rect 4813 55516 4877 55520
rect 4813 55460 4817 55516
rect 4817 55460 4873 55516
rect 4873 55460 4877 55516
rect 4813 55456 4877 55460
rect 4893 55516 4957 55520
rect 4893 55460 4897 55516
rect 4897 55460 4953 55516
rect 4953 55460 4957 55516
rect 4893 55456 4957 55460
rect 4973 55516 5037 55520
rect 4973 55460 4977 55516
rect 4977 55460 5033 55516
rect 5033 55460 5037 55516
rect 4973 55456 5037 55460
rect 5053 55516 5117 55520
rect 5053 55460 5057 55516
rect 5057 55460 5113 55516
rect 5113 55460 5117 55516
rect 5053 55456 5117 55460
rect 4292 55312 4356 55316
rect 4292 55256 4306 55312
rect 4306 55256 4356 55312
rect 4292 55252 4356 55256
rect 1917 54972 1981 54976
rect 1917 54916 1921 54972
rect 1921 54916 1977 54972
rect 1977 54916 1981 54972
rect 1917 54912 1981 54916
rect 1997 54972 2061 54976
rect 1997 54916 2001 54972
rect 2001 54916 2057 54972
rect 2057 54916 2061 54972
rect 1997 54912 2061 54916
rect 2077 54972 2141 54976
rect 2077 54916 2081 54972
rect 2081 54916 2137 54972
rect 2137 54916 2141 54972
rect 2077 54912 2141 54916
rect 2157 54972 2221 54976
rect 2157 54916 2161 54972
rect 2161 54916 2217 54972
rect 2217 54916 2221 54972
rect 2157 54912 2221 54916
rect 3848 54972 3912 54976
rect 3848 54916 3852 54972
rect 3852 54916 3908 54972
rect 3908 54916 3912 54972
rect 3848 54912 3912 54916
rect 3928 54972 3992 54976
rect 3928 54916 3932 54972
rect 3932 54916 3988 54972
rect 3988 54916 3992 54972
rect 3928 54912 3992 54916
rect 4008 54972 4072 54976
rect 4008 54916 4012 54972
rect 4012 54916 4068 54972
rect 4068 54916 4072 54972
rect 4008 54912 4072 54916
rect 4088 54972 4152 54976
rect 4088 54916 4092 54972
rect 4092 54916 4148 54972
rect 4148 54916 4152 54972
rect 4088 54912 4152 54916
rect 5778 54972 5842 54976
rect 5778 54916 5782 54972
rect 5782 54916 5838 54972
rect 5838 54916 5842 54972
rect 5778 54912 5842 54916
rect 5858 54972 5922 54976
rect 5858 54916 5862 54972
rect 5862 54916 5918 54972
rect 5918 54916 5922 54972
rect 5858 54912 5922 54916
rect 5938 54972 6002 54976
rect 5938 54916 5942 54972
rect 5942 54916 5998 54972
rect 5998 54916 6002 54972
rect 5938 54912 6002 54916
rect 6018 54972 6082 54976
rect 6018 54916 6022 54972
rect 6022 54916 6078 54972
rect 6078 54916 6082 54972
rect 6018 54912 6082 54916
rect 2882 54428 2946 54432
rect 2882 54372 2886 54428
rect 2886 54372 2942 54428
rect 2942 54372 2946 54428
rect 2882 54368 2946 54372
rect 2962 54428 3026 54432
rect 2962 54372 2966 54428
rect 2966 54372 3022 54428
rect 3022 54372 3026 54428
rect 2962 54368 3026 54372
rect 3042 54428 3106 54432
rect 3042 54372 3046 54428
rect 3046 54372 3102 54428
rect 3102 54372 3106 54428
rect 3042 54368 3106 54372
rect 3122 54428 3186 54432
rect 3122 54372 3126 54428
rect 3126 54372 3182 54428
rect 3182 54372 3186 54428
rect 3122 54368 3186 54372
rect 4813 54428 4877 54432
rect 4813 54372 4817 54428
rect 4817 54372 4873 54428
rect 4873 54372 4877 54428
rect 4813 54368 4877 54372
rect 4893 54428 4957 54432
rect 4893 54372 4897 54428
rect 4897 54372 4953 54428
rect 4953 54372 4957 54428
rect 4893 54368 4957 54372
rect 4973 54428 5037 54432
rect 4973 54372 4977 54428
rect 4977 54372 5033 54428
rect 5033 54372 5037 54428
rect 4973 54368 5037 54372
rect 5053 54428 5117 54432
rect 5053 54372 5057 54428
rect 5057 54372 5113 54428
rect 5113 54372 5117 54428
rect 5053 54368 5117 54372
rect 1917 53884 1981 53888
rect 1917 53828 1921 53884
rect 1921 53828 1977 53884
rect 1977 53828 1981 53884
rect 1917 53824 1981 53828
rect 1997 53884 2061 53888
rect 1997 53828 2001 53884
rect 2001 53828 2057 53884
rect 2057 53828 2061 53884
rect 1997 53824 2061 53828
rect 2077 53884 2141 53888
rect 2077 53828 2081 53884
rect 2081 53828 2137 53884
rect 2137 53828 2141 53884
rect 2077 53824 2141 53828
rect 2157 53884 2221 53888
rect 2157 53828 2161 53884
rect 2161 53828 2217 53884
rect 2217 53828 2221 53884
rect 2157 53824 2221 53828
rect 3848 53884 3912 53888
rect 3848 53828 3852 53884
rect 3852 53828 3908 53884
rect 3908 53828 3912 53884
rect 3848 53824 3912 53828
rect 3928 53884 3992 53888
rect 3928 53828 3932 53884
rect 3932 53828 3988 53884
rect 3988 53828 3992 53884
rect 3928 53824 3992 53828
rect 4008 53884 4072 53888
rect 4008 53828 4012 53884
rect 4012 53828 4068 53884
rect 4068 53828 4072 53884
rect 4008 53824 4072 53828
rect 4088 53884 4152 53888
rect 4088 53828 4092 53884
rect 4092 53828 4148 53884
rect 4148 53828 4152 53884
rect 4088 53824 4152 53828
rect 5778 53884 5842 53888
rect 5778 53828 5782 53884
rect 5782 53828 5838 53884
rect 5838 53828 5842 53884
rect 5778 53824 5842 53828
rect 5858 53884 5922 53888
rect 5858 53828 5862 53884
rect 5862 53828 5918 53884
rect 5918 53828 5922 53884
rect 5858 53824 5922 53828
rect 5938 53884 6002 53888
rect 5938 53828 5942 53884
rect 5942 53828 5998 53884
rect 5998 53828 6002 53884
rect 5938 53824 6002 53828
rect 6018 53884 6082 53888
rect 6018 53828 6022 53884
rect 6022 53828 6078 53884
rect 6078 53828 6082 53884
rect 6018 53824 6082 53828
rect 2882 53340 2946 53344
rect 2882 53284 2886 53340
rect 2886 53284 2942 53340
rect 2942 53284 2946 53340
rect 2882 53280 2946 53284
rect 2962 53340 3026 53344
rect 2962 53284 2966 53340
rect 2966 53284 3022 53340
rect 3022 53284 3026 53340
rect 2962 53280 3026 53284
rect 3042 53340 3106 53344
rect 3042 53284 3046 53340
rect 3046 53284 3102 53340
rect 3102 53284 3106 53340
rect 3042 53280 3106 53284
rect 3122 53340 3186 53344
rect 3122 53284 3126 53340
rect 3126 53284 3182 53340
rect 3182 53284 3186 53340
rect 3122 53280 3186 53284
rect 4813 53340 4877 53344
rect 4813 53284 4817 53340
rect 4817 53284 4873 53340
rect 4873 53284 4877 53340
rect 4813 53280 4877 53284
rect 4893 53340 4957 53344
rect 4893 53284 4897 53340
rect 4897 53284 4953 53340
rect 4953 53284 4957 53340
rect 4893 53280 4957 53284
rect 4973 53340 5037 53344
rect 4973 53284 4977 53340
rect 4977 53284 5033 53340
rect 5033 53284 5037 53340
rect 4973 53280 5037 53284
rect 5053 53340 5117 53344
rect 5053 53284 5057 53340
rect 5057 53284 5113 53340
rect 5113 53284 5117 53340
rect 5053 53280 5117 53284
rect 1917 52796 1981 52800
rect 1917 52740 1921 52796
rect 1921 52740 1977 52796
rect 1977 52740 1981 52796
rect 1917 52736 1981 52740
rect 1997 52796 2061 52800
rect 1997 52740 2001 52796
rect 2001 52740 2057 52796
rect 2057 52740 2061 52796
rect 1997 52736 2061 52740
rect 2077 52796 2141 52800
rect 2077 52740 2081 52796
rect 2081 52740 2137 52796
rect 2137 52740 2141 52796
rect 2077 52736 2141 52740
rect 2157 52796 2221 52800
rect 2157 52740 2161 52796
rect 2161 52740 2217 52796
rect 2217 52740 2221 52796
rect 2157 52736 2221 52740
rect 3848 52796 3912 52800
rect 3848 52740 3852 52796
rect 3852 52740 3908 52796
rect 3908 52740 3912 52796
rect 3848 52736 3912 52740
rect 3928 52796 3992 52800
rect 3928 52740 3932 52796
rect 3932 52740 3988 52796
rect 3988 52740 3992 52796
rect 3928 52736 3992 52740
rect 4008 52796 4072 52800
rect 4008 52740 4012 52796
rect 4012 52740 4068 52796
rect 4068 52740 4072 52796
rect 4008 52736 4072 52740
rect 4088 52796 4152 52800
rect 4088 52740 4092 52796
rect 4092 52740 4148 52796
rect 4148 52740 4152 52796
rect 4088 52736 4152 52740
rect 5778 52796 5842 52800
rect 5778 52740 5782 52796
rect 5782 52740 5838 52796
rect 5838 52740 5842 52796
rect 5778 52736 5842 52740
rect 5858 52796 5922 52800
rect 5858 52740 5862 52796
rect 5862 52740 5918 52796
rect 5918 52740 5922 52796
rect 5858 52736 5922 52740
rect 5938 52796 6002 52800
rect 5938 52740 5942 52796
rect 5942 52740 5998 52796
rect 5998 52740 6002 52796
rect 5938 52736 6002 52740
rect 6018 52796 6082 52800
rect 6018 52740 6022 52796
rect 6022 52740 6078 52796
rect 6078 52740 6082 52796
rect 6018 52736 6082 52740
rect 2882 52252 2946 52256
rect 2882 52196 2886 52252
rect 2886 52196 2942 52252
rect 2942 52196 2946 52252
rect 2882 52192 2946 52196
rect 2962 52252 3026 52256
rect 2962 52196 2966 52252
rect 2966 52196 3022 52252
rect 3022 52196 3026 52252
rect 2962 52192 3026 52196
rect 3042 52252 3106 52256
rect 3042 52196 3046 52252
rect 3046 52196 3102 52252
rect 3102 52196 3106 52252
rect 3042 52192 3106 52196
rect 3122 52252 3186 52256
rect 3122 52196 3126 52252
rect 3126 52196 3182 52252
rect 3182 52196 3186 52252
rect 3122 52192 3186 52196
rect 4813 52252 4877 52256
rect 4813 52196 4817 52252
rect 4817 52196 4873 52252
rect 4873 52196 4877 52252
rect 4813 52192 4877 52196
rect 4893 52252 4957 52256
rect 4893 52196 4897 52252
rect 4897 52196 4953 52252
rect 4953 52196 4957 52252
rect 4893 52192 4957 52196
rect 4973 52252 5037 52256
rect 4973 52196 4977 52252
rect 4977 52196 5033 52252
rect 5033 52196 5037 52252
rect 4973 52192 5037 52196
rect 5053 52252 5117 52256
rect 5053 52196 5057 52252
rect 5057 52196 5113 52252
rect 5113 52196 5117 52252
rect 5053 52192 5117 52196
rect 1917 51708 1981 51712
rect 1917 51652 1921 51708
rect 1921 51652 1977 51708
rect 1977 51652 1981 51708
rect 1917 51648 1981 51652
rect 1997 51708 2061 51712
rect 1997 51652 2001 51708
rect 2001 51652 2057 51708
rect 2057 51652 2061 51708
rect 1997 51648 2061 51652
rect 2077 51708 2141 51712
rect 2077 51652 2081 51708
rect 2081 51652 2137 51708
rect 2137 51652 2141 51708
rect 2077 51648 2141 51652
rect 2157 51708 2221 51712
rect 2157 51652 2161 51708
rect 2161 51652 2217 51708
rect 2217 51652 2221 51708
rect 2157 51648 2221 51652
rect 3848 51708 3912 51712
rect 3848 51652 3852 51708
rect 3852 51652 3908 51708
rect 3908 51652 3912 51708
rect 3848 51648 3912 51652
rect 3928 51708 3992 51712
rect 3928 51652 3932 51708
rect 3932 51652 3988 51708
rect 3988 51652 3992 51708
rect 3928 51648 3992 51652
rect 4008 51708 4072 51712
rect 4008 51652 4012 51708
rect 4012 51652 4068 51708
rect 4068 51652 4072 51708
rect 4008 51648 4072 51652
rect 4088 51708 4152 51712
rect 4088 51652 4092 51708
rect 4092 51652 4148 51708
rect 4148 51652 4152 51708
rect 4088 51648 4152 51652
rect 5778 51708 5842 51712
rect 5778 51652 5782 51708
rect 5782 51652 5838 51708
rect 5838 51652 5842 51708
rect 5778 51648 5842 51652
rect 5858 51708 5922 51712
rect 5858 51652 5862 51708
rect 5862 51652 5918 51708
rect 5918 51652 5922 51708
rect 5858 51648 5922 51652
rect 5938 51708 6002 51712
rect 5938 51652 5942 51708
rect 5942 51652 5998 51708
rect 5998 51652 6002 51708
rect 5938 51648 6002 51652
rect 6018 51708 6082 51712
rect 6018 51652 6022 51708
rect 6022 51652 6078 51708
rect 6078 51652 6082 51708
rect 6018 51648 6082 51652
rect 2882 51164 2946 51168
rect 2882 51108 2886 51164
rect 2886 51108 2942 51164
rect 2942 51108 2946 51164
rect 2882 51104 2946 51108
rect 2962 51164 3026 51168
rect 2962 51108 2966 51164
rect 2966 51108 3022 51164
rect 3022 51108 3026 51164
rect 2962 51104 3026 51108
rect 3042 51164 3106 51168
rect 3042 51108 3046 51164
rect 3046 51108 3102 51164
rect 3102 51108 3106 51164
rect 3042 51104 3106 51108
rect 3122 51164 3186 51168
rect 3122 51108 3126 51164
rect 3126 51108 3182 51164
rect 3182 51108 3186 51164
rect 3122 51104 3186 51108
rect 4813 51164 4877 51168
rect 4813 51108 4817 51164
rect 4817 51108 4873 51164
rect 4873 51108 4877 51164
rect 4813 51104 4877 51108
rect 4893 51164 4957 51168
rect 4893 51108 4897 51164
rect 4897 51108 4953 51164
rect 4953 51108 4957 51164
rect 4893 51104 4957 51108
rect 4973 51164 5037 51168
rect 4973 51108 4977 51164
rect 4977 51108 5033 51164
rect 5033 51108 5037 51164
rect 4973 51104 5037 51108
rect 5053 51164 5117 51168
rect 5053 51108 5057 51164
rect 5057 51108 5113 51164
rect 5113 51108 5117 51164
rect 5053 51104 5117 51108
rect 1917 50620 1981 50624
rect 1917 50564 1921 50620
rect 1921 50564 1977 50620
rect 1977 50564 1981 50620
rect 1917 50560 1981 50564
rect 1997 50620 2061 50624
rect 1997 50564 2001 50620
rect 2001 50564 2057 50620
rect 2057 50564 2061 50620
rect 1997 50560 2061 50564
rect 2077 50620 2141 50624
rect 2077 50564 2081 50620
rect 2081 50564 2137 50620
rect 2137 50564 2141 50620
rect 2077 50560 2141 50564
rect 2157 50620 2221 50624
rect 2157 50564 2161 50620
rect 2161 50564 2217 50620
rect 2217 50564 2221 50620
rect 2157 50560 2221 50564
rect 3848 50620 3912 50624
rect 3848 50564 3852 50620
rect 3852 50564 3908 50620
rect 3908 50564 3912 50620
rect 3848 50560 3912 50564
rect 3928 50620 3992 50624
rect 3928 50564 3932 50620
rect 3932 50564 3988 50620
rect 3988 50564 3992 50620
rect 3928 50560 3992 50564
rect 4008 50620 4072 50624
rect 4008 50564 4012 50620
rect 4012 50564 4068 50620
rect 4068 50564 4072 50620
rect 4008 50560 4072 50564
rect 4088 50620 4152 50624
rect 4088 50564 4092 50620
rect 4092 50564 4148 50620
rect 4148 50564 4152 50620
rect 4088 50560 4152 50564
rect 5778 50620 5842 50624
rect 5778 50564 5782 50620
rect 5782 50564 5838 50620
rect 5838 50564 5842 50620
rect 5778 50560 5842 50564
rect 5858 50620 5922 50624
rect 5858 50564 5862 50620
rect 5862 50564 5918 50620
rect 5918 50564 5922 50620
rect 5858 50560 5922 50564
rect 5938 50620 6002 50624
rect 5938 50564 5942 50620
rect 5942 50564 5998 50620
rect 5998 50564 6002 50620
rect 5938 50560 6002 50564
rect 6018 50620 6082 50624
rect 6018 50564 6022 50620
rect 6022 50564 6078 50620
rect 6078 50564 6082 50620
rect 6018 50560 6082 50564
rect 2882 50076 2946 50080
rect 2882 50020 2886 50076
rect 2886 50020 2942 50076
rect 2942 50020 2946 50076
rect 2882 50016 2946 50020
rect 2962 50076 3026 50080
rect 2962 50020 2966 50076
rect 2966 50020 3022 50076
rect 3022 50020 3026 50076
rect 2962 50016 3026 50020
rect 3042 50076 3106 50080
rect 3042 50020 3046 50076
rect 3046 50020 3102 50076
rect 3102 50020 3106 50076
rect 3042 50016 3106 50020
rect 3122 50076 3186 50080
rect 3122 50020 3126 50076
rect 3126 50020 3182 50076
rect 3182 50020 3186 50076
rect 3122 50016 3186 50020
rect 4813 50076 4877 50080
rect 4813 50020 4817 50076
rect 4817 50020 4873 50076
rect 4873 50020 4877 50076
rect 4813 50016 4877 50020
rect 4893 50076 4957 50080
rect 4893 50020 4897 50076
rect 4897 50020 4953 50076
rect 4953 50020 4957 50076
rect 4893 50016 4957 50020
rect 4973 50076 5037 50080
rect 4973 50020 4977 50076
rect 4977 50020 5033 50076
rect 5033 50020 5037 50076
rect 4973 50016 5037 50020
rect 5053 50076 5117 50080
rect 5053 50020 5057 50076
rect 5057 50020 5113 50076
rect 5113 50020 5117 50076
rect 5053 50016 5117 50020
rect 1917 49532 1981 49536
rect 1917 49476 1921 49532
rect 1921 49476 1977 49532
rect 1977 49476 1981 49532
rect 1917 49472 1981 49476
rect 1997 49532 2061 49536
rect 1997 49476 2001 49532
rect 2001 49476 2057 49532
rect 2057 49476 2061 49532
rect 1997 49472 2061 49476
rect 2077 49532 2141 49536
rect 2077 49476 2081 49532
rect 2081 49476 2137 49532
rect 2137 49476 2141 49532
rect 2077 49472 2141 49476
rect 2157 49532 2221 49536
rect 2157 49476 2161 49532
rect 2161 49476 2217 49532
rect 2217 49476 2221 49532
rect 2157 49472 2221 49476
rect 3848 49532 3912 49536
rect 3848 49476 3852 49532
rect 3852 49476 3908 49532
rect 3908 49476 3912 49532
rect 3848 49472 3912 49476
rect 3928 49532 3992 49536
rect 3928 49476 3932 49532
rect 3932 49476 3988 49532
rect 3988 49476 3992 49532
rect 3928 49472 3992 49476
rect 4008 49532 4072 49536
rect 4008 49476 4012 49532
rect 4012 49476 4068 49532
rect 4068 49476 4072 49532
rect 4008 49472 4072 49476
rect 4088 49532 4152 49536
rect 4088 49476 4092 49532
rect 4092 49476 4148 49532
rect 4148 49476 4152 49532
rect 4088 49472 4152 49476
rect 5778 49532 5842 49536
rect 5778 49476 5782 49532
rect 5782 49476 5838 49532
rect 5838 49476 5842 49532
rect 5778 49472 5842 49476
rect 5858 49532 5922 49536
rect 5858 49476 5862 49532
rect 5862 49476 5918 49532
rect 5918 49476 5922 49532
rect 5858 49472 5922 49476
rect 5938 49532 6002 49536
rect 5938 49476 5942 49532
rect 5942 49476 5998 49532
rect 5998 49476 6002 49532
rect 5938 49472 6002 49476
rect 6018 49532 6082 49536
rect 6018 49476 6022 49532
rect 6022 49476 6078 49532
rect 6078 49476 6082 49532
rect 6018 49472 6082 49476
rect 2882 48988 2946 48992
rect 2882 48932 2886 48988
rect 2886 48932 2942 48988
rect 2942 48932 2946 48988
rect 2882 48928 2946 48932
rect 2962 48988 3026 48992
rect 2962 48932 2966 48988
rect 2966 48932 3022 48988
rect 3022 48932 3026 48988
rect 2962 48928 3026 48932
rect 3042 48988 3106 48992
rect 3042 48932 3046 48988
rect 3046 48932 3102 48988
rect 3102 48932 3106 48988
rect 3042 48928 3106 48932
rect 3122 48988 3186 48992
rect 3122 48932 3126 48988
rect 3126 48932 3182 48988
rect 3182 48932 3186 48988
rect 3122 48928 3186 48932
rect 4813 48988 4877 48992
rect 4813 48932 4817 48988
rect 4817 48932 4873 48988
rect 4873 48932 4877 48988
rect 4813 48928 4877 48932
rect 4893 48988 4957 48992
rect 4893 48932 4897 48988
rect 4897 48932 4953 48988
rect 4953 48932 4957 48988
rect 4893 48928 4957 48932
rect 4973 48988 5037 48992
rect 4973 48932 4977 48988
rect 4977 48932 5033 48988
rect 5033 48932 5037 48988
rect 4973 48928 5037 48932
rect 5053 48988 5117 48992
rect 5053 48932 5057 48988
rect 5057 48932 5113 48988
rect 5113 48932 5117 48988
rect 5053 48928 5117 48932
rect 1917 48444 1981 48448
rect 1917 48388 1921 48444
rect 1921 48388 1977 48444
rect 1977 48388 1981 48444
rect 1917 48384 1981 48388
rect 1997 48444 2061 48448
rect 1997 48388 2001 48444
rect 2001 48388 2057 48444
rect 2057 48388 2061 48444
rect 1997 48384 2061 48388
rect 2077 48444 2141 48448
rect 2077 48388 2081 48444
rect 2081 48388 2137 48444
rect 2137 48388 2141 48444
rect 2077 48384 2141 48388
rect 2157 48444 2221 48448
rect 2157 48388 2161 48444
rect 2161 48388 2217 48444
rect 2217 48388 2221 48444
rect 2157 48384 2221 48388
rect 3848 48444 3912 48448
rect 3848 48388 3852 48444
rect 3852 48388 3908 48444
rect 3908 48388 3912 48444
rect 3848 48384 3912 48388
rect 3928 48444 3992 48448
rect 3928 48388 3932 48444
rect 3932 48388 3988 48444
rect 3988 48388 3992 48444
rect 3928 48384 3992 48388
rect 4008 48444 4072 48448
rect 4008 48388 4012 48444
rect 4012 48388 4068 48444
rect 4068 48388 4072 48444
rect 4008 48384 4072 48388
rect 4088 48444 4152 48448
rect 4088 48388 4092 48444
rect 4092 48388 4148 48444
rect 4148 48388 4152 48444
rect 4088 48384 4152 48388
rect 5778 48444 5842 48448
rect 5778 48388 5782 48444
rect 5782 48388 5838 48444
rect 5838 48388 5842 48444
rect 5778 48384 5842 48388
rect 5858 48444 5922 48448
rect 5858 48388 5862 48444
rect 5862 48388 5918 48444
rect 5918 48388 5922 48444
rect 5858 48384 5922 48388
rect 5938 48444 6002 48448
rect 5938 48388 5942 48444
rect 5942 48388 5998 48444
rect 5998 48388 6002 48444
rect 5938 48384 6002 48388
rect 6018 48444 6082 48448
rect 6018 48388 6022 48444
rect 6022 48388 6078 48444
rect 6078 48388 6082 48444
rect 6018 48384 6082 48388
rect 2636 48044 2700 48108
rect 5396 48044 5460 48108
rect 2882 47900 2946 47904
rect 2882 47844 2886 47900
rect 2886 47844 2942 47900
rect 2942 47844 2946 47900
rect 2882 47840 2946 47844
rect 2962 47900 3026 47904
rect 2962 47844 2966 47900
rect 2966 47844 3022 47900
rect 3022 47844 3026 47900
rect 2962 47840 3026 47844
rect 3042 47900 3106 47904
rect 3042 47844 3046 47900
rect 3046 47844 3102 47900
rect 3102 47844 3106 47900
rect 3042 47840 3106 47844
rect 3122 47900 3186 47904
rect 3122 47844 3126 47900
rect 3126 47844 3182 47900
rect 3182 47844 3186 47900
rect 3122 47840 3186 47844
rect 4813 47900 4877 47904
rect 4813 47844 4817 47900
rect 4817 47844 4873 47900
rect 4873 47844 4877 47900
rect 4813 47840 4877 47844
rect 4893 47900 4957 47904
rect 4893 47844 4897 47900
rect 4897 47844 4953 47900
rect 4953 47844 4957 47900
rect 4893 47840 4957 47844
rect 4973 47900 5037 47904
rect 4973 47844 4977 47900
rect 4977 47844 5033 47900
rect 5033 47844 5037 47900
rect 4973 47840 5037 47844
rect 5053 47900 5117 47904
rect 5053 47844 5057 47900
rect 5057 47844 5113 47900
rect 5113 47844 5117 47900
rect 5053 47840 5117 47844
rect 4660 47772 4724 47836
rect 1917 47356 1981 47360
rect 1917 47300 1921 47356
rect 1921 47300 1977 47356
rect 1977 47300 1981 47356
rect 1917 47296 1981 47300
rect 1997 47356 2061 47360
rect 1997 47300 2001 47356
rect 2001 47300 2057 47356
rect 2057 47300 2061 47356
rect 1997 47296 2061 47300
rect 2077 47356 2141 47360
rect 2077 47300 2081 47356
rect 2081 47300 2137 47356
rect 2137 47300 2141 47356
rect 2077 47296 2141 47300
rect 2157 47356 2221 47360
rect 2157 47300 2161 47356
rect 2161 47300 2217 47356
rect 2217 47300 2221 47356
rect 2157 47296 2221 47300
rect 3848 47356 3912 47360
rect 3848 47300 3852 47356
rect 3852 47300 3908 47356
rect 3908 47300 3912 47356
rect 3848 47296 3912 47300
rect 3928 47356 3992 47360
rect 3928 47300 3932 47356
rect 3932 47300 3988 47356
rect 3988 47300 3992 47356
rect 3928 47296 3992 47300
rect 4008 47356 4072 47360
rect 4008 47300 4012 47356
rect 4012 47300 4068 47356
rect 4068 47300 4072 47356
rect 4008 47296 4072 47300
rect 4088 47356 4152 47360
rect 4088 47300 4092 47356
rect 4092 47300 4148 47356
rect 4148 47300 4152 47356
rect 4088 47296 4152 47300
rect 5778 47356 5842 47360
rect 5778 47300 5782 47356
rect 5782 47300 5838 47356
rect 5838 47300 5842 47356
rect 5778 47296 5842 47300
rect 5858 47356 5922 47360
rect 5858 47300 5862 47356
rect 5862 47300 5918 47356
rect 5918 47300 5922 47356
rect 5858 47296 5922 47300
rect 5938 47356 6002 47360
rect 5938 47300 5942 47356
rect 5942 47300 5998 47356
rect 5998 47300 6002 47356
rect 5938 47296 6002 47300
rect 6018 47356 6082 47360
rect 6018 47300 6022 47356
rect 6022 47300 6078 47356
rect 6078 47300 6082 47356
rect 6018 47296 6082 47300
rect 2882 46812 2946 46816
rect 2882 46756 2886 46812
rect 2886 46756 2942 46812
rect 2942 46756 2946 46812
rect 2882 46752 2946 46756
rect 2962 46812 3026 46816
rect 2962 46756 2966 46812
rect 2966 46756 3022 46812
rect 3022 46756 3026 46812
rect 2962 46752 3026 46756
rect 3042 46812 3106 46816
rect 3042 46756 3046 46812
rect 3046 46756 3102 46812
rect 3102 46756 3106 46812
rect 3042 46752 3106 46756
rect 3122 46812 3186 46816
rect 3122 46756 3126 46812
rect 3126 46756 3182 46812
rect 3182 46756 3186 46812
rect 3122 46752 3186 46756
rect 4813 46812 4877 46816
rect 4813 46756 4817 46812
rect 4817 46756 4873 46812
rect 4873 46756 4877 46812
rect 4813 46752 4877 46756
rect 4893 46812 4957 46816
rect 4893 46756 4897 46812
rect 4897 46756 4953 46812
rect 4953 46756 4957 46812
rect 4893 46752 4957 46756
rect 4973 46812 5037 46816
rect 4973 46756 4977 46812
rect 4977 46756 5033 46812
rect 5033 46756 5037 46812
rect 4973 46752 5037 46756
rect 5053 46812 5117 46816
rect 5053 46756 5057 46812
rect 5057 46756 5113 46812
rect 5113 46756 5117 46812
rect 5053 46752 5117 46756
rect 1917 46268 1981 46272
rect 1917 46212 1921 46268
rect 1921 46212 1977 46268
rect 1977 46212 1981 46268
rect 1917 46208 1981 46212
rect 1997 46268 2061 46272
rect 1997 46212 2001 46268
rect 2001 46212 2057 46268
rect 2057 46212 2061 46268
rect 1997 46208 2061 46212
rect 2077 46268 2141 46272
rect 2077 46212 2081 46268
rect 2081 46212 2137 46268
rect 2137 46212 2141 46268
rect 2077 46208 2141 46212
rect 2157 46268 2221 46272
rect 2157 46212 2161 46268
rect 2161 46212 2217 46268
rect 2217 46212 2221 46268
rect 2157 46208 2221 46212
rect 3848 46268 3912 46272
rect 3848 46212 3852 46268
rect 3852 46212 3908 46268
rect 3908 46212 3912 46268
rect 3848 46208 3912 46212
rect 3928 46268 3992 46272
rect 3928 46212 3932 46268
rect 3932 46212 3988 46268
rect 3988 46212 3992 46268
rect 3928 46208 3992 46212
rect 4008 46268 4072 46272
rect 4008 46212 4012 46268
rect 4012 46212 4068 46268
rect 4068 46212 4072 46268
rect 4008 46208 4072 46212
rect 4088 46268 4152 46272
rect 4088 46212 4092 46268
rect 4092 46212 4148 46268
rect 4148 46212 4152 46268
rect 4088 46208 4152 46212
rect 5778 46268 5842 46272
rect 5778 46212 5782 46268
rect 5782 46212 5838 46268
rect 5838 46212 5842 46268
rect 5778 46208 5842 46212
rect 5858 46268 5922 46272
rect 5858 46212 5862 46268
rect 5862 46212 5918 46268
rect 5918 46212 5922 46268
rect 5858 46208 5922 46212
rect 5938 46268 6002 46272
rect 5938 46212 5942 46268
rect 5942 46212 5998 46268
rect 5998 46212 6002 46268
rect 5938 46208 6002 46212
rect 6018 46268 6082 46272
rect 6018 46212 6022 46268
rect 6022 46212 6078 46268
rect 6078 46212 6082 46268
rect 6018 46208 6082 46212
rect 2882 45724 2946 45728
rect 2882 45668 2886 45724
rect 2886 45668 2942 45724
rect 2942 45668 2946 45724
rect 2882 45664 2946 45668
rect 2962 45724 3026 45728
rect 2962 45668 2966 45724
rect 2966 45668 3022 45724
rect 3022 45668 3026 45724
rect 2962 45664 3026 45668
rect 3042 45724 3106 45728
rect 3042 45668 3046 45724
rect 3046 45668 3102 45724
rect 3102 45668 3106 45724
rect 3042 45664 3106 45668
rect 3122 45724 3186 45728
rect 3122 45668 3126 45724
rect 3126 45668 3182 45724
rect 3182 45668 3186 45724
rect 3122 45664 3186 45668
rect 4813 45724 4877 45728
rect 4813 45668 4817 45724
rect 4817 45668 4873 45724
rect 4873 45668 4877 45724
rect 4813 45664 4877 45668
rect 4893 45724 4957 45728
rect 4893 45668 4897 45724
rect 4897 45668 4953 45724
rect 4953 45668 4957 45724
rect 4893 45664 4957 45668
rect 4973 45724 5037 45728
rect 4973 45668 4977 45724
rect 4977 45668 5033 45724
rect 5033 45668 5037 45724
rect 4973 45664 5037 45668
rect 5053 45724 5117 45728
rect 5053 45668 5057 45724
rect 5057 45668 5113 45724
rect 5113 45668 5117 45724
rect 5053 45664 5117 45668
rect 5212 45324 5276 45388
rect 1917 45180 1981 45184
rect 1917 45124 1921 45180
rect 1921 45124 1977 45180
rect 1977 45124 1981 45180
rect 1917 45120 1981 45124
rect 1997 45180 2061 45184
rect 1997 45124 2001 45180
rect 2001 45124 2057 45180
rect 2057 45124 2061 45180
rect 1997 45120 2061 45124
rect 2077 45180 2141 45184
rect 2077 45124 2081 45180
rect 2081 45124 2137 45180
rect 2137 45124 2141 45180
rect 2077 45120 2141 45124
rect 2157 45180 2221 45184
rect 2157 45124 2161 45180
rect 2161 45124 2217 45180
rect 2217 45124 2221 45180
rect 2157 45120 2221 45124
rect 3848 45180 3912 45184
rect 3848 45124 3852 45180
rect 3852 45124 3908 45180
rect 3908 45124 3912 45180
rect 3848 45120 3912 45124
rect 3928 45180 3992 45184
rect 3928 45124 3932 45180
rect 3932 45124 3988 45180
rect 3988 45124 3992 45180
rect 3928 45120 3992 45124
rect 4008 45180 4072 45184
rect 4008 45124 4012 45180
rect 4012 45124 4068 45180
rect 4068 45124 4072 45180
rect 4008 45120 4072 45124
rect 4088 45180 4152 45184
rect 4088 45124 4092 45180
rect 4092 45124 4148 45180
rect 4148 45124 4152 45180
rect 4088 45120 4152 45124
rect 5778 45180 5842 45184
rect 5778 45124 5782 45180
rect 5782 45124 5838 45180
rect 5838 45124 5842 45180
rect 5778 45120 5842 45124
rect 5858 45180 5922 45184
rect 5858 45124 5862 45180
rect 5862 45124 5918 45180
rect 5918 45124 5922 45180
rect 5858 45120 5922 45124
rect 5938 45180 6002 45184
rect 5938 45124 5942 45180
rect 5942 45124 5998 45180
rect 5998 45124 6002 45180
rect 5938 45120 6002 45124
rect 6018 45180 6082 45184
rect 6018 45124 6022 45180
rect 6022 45124 6078 45180
rect 6078 45124 6082 45180
rect 6018 45120 6082 45124
rect 2882 44636 2946 44640
rect 2882 44580 2886 44636
rect 2886 44580 2942 44636
rect 2942 44580 2946 44636
rect 2882 44576 2946 44580
rect 2962 44636 3026 44640
rect 2962 44580 2966 44636
rect 2966 44580 3022 44636
rect 3022 44580 3026 44636
rect 2962 44576 3026 44580
rect 3042 44636 3106 44640
rect 3042 44580 3046 44636
rect 3046 44580 3102 44636
rect 3102 44580 3106 44636
rect 3042 44576 3106 44580
rect 3122 44636 3186 44640
rect 3122 44580 3126 44636
rect 3126 44580 3182 44636
rect 3182 44580 3186 44636
rect 3122 44576 3186 44580
rect 4813 44636 4877 44640
rect 4813 44580 4817 44636
rect 4817 44580 4873 44636
rect 4873 44580 4877 44636
rect 4813 44576 4877 44580
rect 4893 44636 4957 44640
rect 4893 44580 4897 44636
rect 4897 44580 4953 44636
rect 4953 44580 4957 44636
rect 4893 44576 4957 44580
rect 4973 44636 5037 44640
rect 4973 44580 4977 44636
rect 4977 44580 5033 44636
rect 5033 44580 5037 44636
rect 4973 44576 5037 44580
rect 5053 44636 5117 44640
rect 5053 44580 5057 44636
rect 5057 44580 5113 44636
rect 5113 44580 5117 44636
rect 5053 44576 5117 44580
rect 1917 44092 1981 44096
rect 1917 44036 1921 44092
rect 1921 44036 1977 44092
rect 1977 44036 1981 44092
rect 1917 44032 1981 44036
rect 1997 44092 2061 44096
rect 1997 44036 2001 44092
rect 2001 44036 2057 44092
rect 2057 44036 2061 44092
rect 1997 44032 2061 44036
rect 2077 44092 2141 44096
rect 2077 44036 2081 44092
rect 2081 44036 2137 44092
rect 2137 44036 2141 44092
rect 2077 44032 2141 44036
rect 2157 44092 2221 44096
rect 2157 44036 2161 44092
rect 2161 44036 2217 44092
rect 2217 44036 2221 44092
rect 2157 44032 2221 44036
rect 3848 44092 3912 44096
rect 3848 44036 3852 44092
rect 3852 44036 3908 44092
rect 3908 44036 3912 44092
rect 3848 44032 3912 44036
rect 3928 44092 3992 44096
rect 3928 44036 3932 44092
rect 3932 44036 3988 44092
rect 3988 44036 3992 44092
rect 3928 44032 3992 44036
rect 4008 44092 4072 44096
rect 4008 44036 4012 44092
rect 4012 44036 4068 44092
rect 4068 44036 4072 44092
rect 4008 44032 4072 44036
rect 4088 44092 4152 44096
rect 4088 44036 4092 44092
rect 4092 44036 4148 44092
rect 4148 44036 4152 44092
rect 4088 44032 4152 44036
rect 5778 44092 5842 44096
rect 5778 44036 5782 44092
rect 5782 44036 5838 44092
rect 5838 44036 5842 44092
rect 5778 44032 5842 44036
rect 5858 44092 5922 44096
rect 5858 44036 5862 44092
rect 5862 44036 5918 44092
rect 5918 44036 5922 44092
rect 5858 44032 5922 44036
rect 5938 44092 6002 44096
rect 5938 44036 5942 44092
rect 5942 44036 5998 44092
rect 5998 44036 6002 44092
rect 5938 44032 6002 44036
rect 6018 44092 6082 44096
rect 6018 44036 6022 44092
rect 6022 44036 6078 44092
rect 6078 44036 6082 44092
rect 6018 44032 6082 44036
rect 3372 43692 3436 43756
rect 2882 43548 2946 43552
rect 2882 43492 2886 43548
rect 2886 43492 2942 43548
rect 2942 43492 2946 43548
rect 2882 43488 2946 43492
rect 2962 43548 3026 43552
rect 2962 43492 2966 43548
rect 2966 43492 3022 43548
rect 3022 43492 3026 43548
rect 2962 43488 3026 43492
rect 3042 43548 3106 43552
rect 3042 43492 3046 43548
rect 3046 43492 3102 43548
rect 3102 43492 3106 43548
rect 3042 43488 3106 43492
rect 3122 43548 3186 43552
rect 3122 43492 3126 43548
rect 3126 43492 3182 43548
rect 3182 43492 3186 43548
rect 3122 43488 3186 43492
rect 4813 43548 4877 43552
rect 4813 43492 4817 43548
rect 4817 43492 4873 43548
rect 4873 43492 4877 43548
rect 4813 43488 4877 43492
rect 4893 43548 4957 43552
rect 4893 43492 4897 43548
rect 4897 43492 4953 43548
rect 4953 43492 4957 43548
rect 4893 43488 4957 43492
rect 4973 43548 5037 43552
rect 4973 43492 4977 43548
rect 4977 43492 5033 43548
rect 5033 43492 5037 43548
rect 4973 43488 5037 43492
rect 5053 43548 5117 43552
rect 5053 43492 5057 43548
rect 5057 43492 5113 43548
rect 5113 43492 5117 43548
rect 5053 43488 5117 43492
rect 5580 43284 5644 43348
rect 1917 43004 1981 43008
rect 1917 42948 1921 43004
rect 1921 42948 1977 43004
rect 1977 42948 1981 43004
rect 1917 42944 1981 42948
rect 1997 43004 2061 43008
rect 1997 42948 2001 43004
rect 2001 42948 2057 43004
rect 2057 42948 2061 43004
rect 1997 42944 2061 42948
rect 2077 43004 2141 43008
rect 2077 42948 2081 43004
rect 2081 42948 2137 43004
rect 2137 42948 2141 43004
rect 2077 42944 2141 42948
rect 2157 43004 2221 43008
rect 2157 42948 2161 43004
rect 2161 42948 2217 43004
rect 2217 42948 2221 43004
rect 2157 42944 2221 42948
rect 3848 43004 3912 43008
rect 3848 42948 3852 43004
rect 3852 42948 3908 43004
rect 3908 42948 3912 43004
rect 3848 42944 3912 42948
rect 3928 43004 3992 43008
rect 3928 42948 3932 43004
rect 3932 42948 3988 43004
rect 3988 42948 3992 43004
rect 3928 42944 3992 42948
rect 4008 43004 4072 43008
rect 4008 42948 4012 43004
rect 4012 42948 4068 43004
rect 4068 42948 4072 43004
rect 4008 42944 4072 42948
rect 4088 43004 4152 43008
rect 4088 42948 4092 43004
rect 4092 42948 4148 43004
rect 4148 42948 4152 43004
rect 4088 42944 4152 42948
rect 5778 43004 5842 43008
rect 5778 42948 5782 43004
rect 5782 42948 5838 43004
rect 5838 42948 5842 43004
rect 5778 42944 5842 42948
rect 5858 43004 5922 43008
rect 5858 42948 5862 43004
rect 5862 42948 5918 43004
rect 5918 42948 5922 43004
rect 5858 42944 5922 42948
rect 5938 43004 6002 43008
rect 5938 42948 5942 43004
rect 5942 42948 5998 43004
rect 5998 42948 6002 43004
rect 5938 42944 6002 42948
rect 6018 43004 6082 43008
rect 6018 42948 6022 43004
rect 6022 42948 6078 43004
rect 6078 42948 6082 43004
rect 6018 42944 6082 42948
rect 2882 42460 2946 42464
rect 2882 42404 2886 42460
rect 2886 42404 2942 42460
rect 2942 42404 2946 42460
rect 2882 42400 2946 42404
rect 2962 42460 3026 42464
rect 2962 42404 2966 42460
rect 2966 42404 3022 42460
rect 3022 42404 3026 42460
rect 2962 42400 3026 42404
rect 3042 42460 3106 42464
rect 3042 42404 3046 42460
rect 3046 42404 3102 42460
rect 3102 42404 3106 42460
rect 3042 42400 3106 42404
rect 3122 42460 3186 42464
rect 3122 42404 3126 42460
rect 3126 42404 3182 42460
rect 3182 42404 3186 42460
rect 3122 42400 3186 42404
rect 4813 42460 4877 42464
rect 4813 42404 4817 42460
rect 4817 42404 4873 42460
rect 4873 42404 4877 42460
rect 4813 42400 4877 42404
rect 4893 42460 4957 42464
rect 4893 42404 4897 42460
rect 4897 42404 4953 42460
rect 4953 42404 4957 42460
rect 4893 42400 4957 42404
rect 4973 42460 5037 42464
rect 4973 42404 4977 42460
rect 4977 42404 5033 42460
rect 5033 42404 5037 42460
rect 4973 42400 5037 42404
rect 5053 42460 5117 42464
rect 5053 42404 5057 42460
rect 5057 42404 5113 42460
rect 5113 42404 5117 42460
rect 5053 42400 5117 42404
rect 4660 42196 4724 42260
rect 3556 42060 3620 42124
rect 4660 41984 4724 41988
rect 4660 41928 4710 41984
rect 4710 41928 4724 41984
rect 4660 41924 4724 41928
rect 1917 41916 1981 41920
rect 1917 41860 1921 41916
rect 1921 41860 1977 41916
rect 1977 41860 1981 41916
rect 1917 41856 1981 41860
rect 1997 41916 2061 41920
rect 1997 41860 2001 41916
rect 2001 41860 2057 41916
rect 2057 41860 2061 41916
rect 1997 41856 2061 41860
rect 2077 41916 2141 41920
rect 2077 41860 2081 41916
rect 2081 41860 2137 41916
rect 2137 41860 2141 41916
rect 2077 41856 2141 41860
rect 2157 41916 2221 41920
rect 2157 41860 2161 41916
rect 2161 41860 2217 41916
rect 2217 41860 2221 41916
rect 2157 41856 2221 41860
rect 3848 41916 3912 41920
rect 3848 41860 3852 41916
rect 3852 41860 3908 41916
rect 3908 41860 3912 41916
rect 3848 41856 3912 41860
rect 3928 41916 3992 41920
rect 3928 41860 3932 41916
rect 3932 41860 3988 41916
rect 3988 41860 3992 41916
rect 3928 41856 3992 41860
rect 4008 41916 4072 41920
rect 4008 41860 4012 41916
rect 4012 41860 4068 41916
rect 4068 41860 4072 41916
rect 4008 41856 4072 41860
rect 4088 41916 4152 41920
rect 4088 41860 4092 41916
rect 4092 41860 4148 41916
rect 4148 41860 4152 41916
rect 4088 41856 4152 41860
rect 5778 41916 5842 41920
rect 5778 41860 5782 41916
rect 5782 41860 5838 41916
rect 5838 41860 5842 41916
rect 5778 41856 5842 41860
rect 5858 41916 5922 41920
rect 5858 41860 5862 41916
rect 5862 41860 5918 41916
rect 5918 41860 5922 41916
rect 5858 41856 5922 41860
rect 5938 41916 6002 41920
rect 5938 41860 5942 41916
rect 5942 41860 5998 41916
rect 5998 41860 6002 41916
rect 5938 41856 6002 41860
rect 6018 41916 6082 41920
rect 6018 41860 6022 41916
rect 6022 41860 6078 41916
rect 6078 41860 6082 41916
rect 6018 41856 6082 41860
rect 4476 41848 4540 41852
rect 4476 41792 4526 41848
rect 4526 41792 4540 41848
rect 4476 41788 4540 41792
rect 5396 41652 5460 41716
rect 1716 41516 1780 41580
rect 2882 41372 2946 41376
rect 2882 41316 2886 41372
rect 2886 41316 2942 41372
rect 2942 41316 2946 41372
rect 2882 41312 2946 41316
rect 2962 41372 3026 41376
rect 2962 41316 2966 41372
rect 2966 41316 3022 41372
rect 3022 41316 3026 41372
rect 2962 41312 3026 41316
rect 3042 41372 3106 41376
rect 3042 41316 3046 41372
rect 3046 41316 3102 41372
rect 3102 41316 3106 41372
rect 3042 41312 3106 41316
rect 3122 41372 3186 41376
rect 3122 41316 3126 41372
rect 3126 41316 3182 41372
rect 3182 41316 3186 41372
rect 3122 41312 3186 41316
rect 3372 41108 3436 41172
rect 4813 41372 4877 41376
rect 4813 41316 4817 41372
rect 4817 41316 4873 41372
rect 4873 41316 4877 41372
rect 4813 41312 4877 41316
rect 4893 41372 4957 41376
rect 4893 41316 4897 41372
rect 4897 41316 4953 41372
rect 4953 41316 4957 41372
rect 4893 41312 4957 41316
rect 4973 41372 5037 41376
rect 4973 41316 4977 41372
rect 4977 41316 5033 41372
rect 5033 41316 5037 41372
rect 4973 41312 5037 41316
rect 5053 41372 5117 41376
rect 5053 41316 5057 41372
rect 5057 41316 5113 41372
rect 5113 41316 5117 41372
rect 5053 41312 5117 41316
rect 4660 41244 4724 41308
rect 4476 40972 4540 41036
rect 5212 40836 5276 40900
rect 1917 40828 1981 40832
rect 1917 40772 1921 40828
rect 1921 40772 1977 40828
rect 1977 40772 1981 40828
rect 1917 40768 1981 40772
rect 1997 40828 2061 40832
rect 1997 40772 2001 40828
rect 2001 40772 2057 40828
rect 2057 40772 2061 40828
rect 1997 40768 2061 40772
rect 2077 40828 2141 40832
rect 2077 40772 2081 40828
rect 2081 40772 2137 40828
rect 2137 40772 2141 40828
rect 2077 40768 2141 40772
rect 2157 40828 2221 40832
rect 2157 40772 2161 40828
rect 2161 40772 2217 40828
rect 2217 40772 2221 40828
rect 2157 40768 2221 40772
rect 3848 40828 3912 40832
rect 3848 40772 3852 40828
rect 3852 40772 3908 40828
rect 3908 40772 3912 40828
rect 3848 40768 3912 40772
rect 3928 40828 3992 40832
rect 3928 40772 3932 40828
rect 3932 40772 3988 40828
rect 3988 40772 3992 40828
rect 3928 40768 3992 40772
rect 4008 40828 4072 40832
rect 4008 40772 4012 40828
rect 4012 40772 4068 40828
rect 4068 40772 4072 40828
rect 4008 40768 4072 40772
rect 4088 40828 4152 40832
rect 4088 40772 4092 40828
rect 4092 40772 4148 40828
rect 4148 40772 4152 40828
rect 4088 40768 4152 40772
rect 5778 40828 5842 40832
rect 5778 40772 5782 40828
rect 5782 40772 5838 40828
rect 5838 40772 5842 40828
rect 5778 40768 5842 40772
rect 5858 40828 5922 40832
rect 5858 40772 5862 40828
rect 5862 40772 5918 40828
rect 5918 40772 5922 40828
rect 5858 40768 5922 40772
rect 5938 40828 6002 40832
rect 5938 40772 5942 40828
rect 5942 40772 5998 40828
rect 5998 40772 6002 40828
rect 5938 40768 6002 40772
rect 6018 40828 6082 40832
rect 6018 40772 6022 40828
rect 6022 40772 6078 40828
rect 6078 40772 6082 40828
rect 6018 40768 6082 40772
rect 2882 40284 2946 40288
rect 2882 40228 2886 40284
rect 2886 40228 2942 40284
rect 2942 40228 2946 40284
rect 2882 40224 2946 40228
rect 2962 40284 3026 40288
rect 2962 40228 2966 40284
rect 2966 40228 3022 40284
rect 3022 40228 3026 40284
rect 2962 40224 3026 40228
rect 3042 40284 3106 40288
rect 3042 40228 3046 40284
rect 3046 40228 3102 40284
rect 3102 40228 3106 40284
rect 3042 40224 3106 40228
rect 3122 40284 3186 40288
rect 3122 40228 3126 40284
rect 3126 40228 3182 40284
rect 3182 40228 3186 40284
rect 3122 40224 3186 40228
rect 4813 40284 4877 40288
rect 4813 40228 4817 40284
rect 4817 40228 4873 40284
rect 4873 40228 4877 40284
rect 4813 40224 4877 40228
rect 4893 40284 4957 40288
rect 4893 40228 4897 40284
rect 4897 40228 4953 40284
rect 4953 40228 4957 40284
rect 4893 40224 4957 40228
rect 4973 40284 5037 40288
rect 4973 40228 4977 40284
rect 4977 40228 5033 40284
rect 5033 40228 5037 40284
rect 4973 40224 5037 40228
rect 5053 40284 5117 40288
rect 5053 40228 5057 40284
rect 5057 40228 5113 40284
rect 5113 40228 5117 40284
rect 5053 40224 5117 40228
rect 1917 39740 1981 39744
rect 1917 39684 1921 39740
rect 1921 39684 1977 39740
rect 1977 39684 1981 39740
rect 1917 39680 1981 39684
rect 1997 39740 2061 39744
rect 1997 39684 2001 39740
rect 2001 39684 2057 39740
rect 2057 39684 2061 39740
rect 1997 39680 2061 39684
rect 2077 39740 2141 39744
rect 2077 39684 2081 39740
rect 2081 39684 2137 39740
rect 2137 39684 2141 39740
rect 2077 39680 2141 39684
rect 2157 39740 2221 39744
rect 2157 39684 2161 39740
rect 2161 39684 2217 39740
rect 2217 39684 2221 39740
rect 2157 39680 2221 39684
rect 3848 39740 3912 39744
rect 3848 39684 3852 39740
rect 3852 39684 3908 39740
rect 3908 39684 3912 39740
rect 3848 39680 3912 39684
rect 3928 39740 3992 39744
rect 3928 39684 3932 39740
rect 3932 39684 3988 39740
rect 3988 39684 3992 39740
rect 3928 39680 3992 39684
rect 4008 39740 4072 39744
rect 4008 39684 4012 39740
rect 4012 39684 4068 39740
rect 4068 39684 4072 39740
rect 4008 39680 4072 39684
rect 4088 39740 4152 39744
rect 4088 39684 4092 39740
rect 4092 39684 4148 39740
rect 4148 39684 4152 39740
rect 4088 39680 4152 39684
rect 5778 39740 5842 39744
rect 5778 39684 5782 39740
rect 5782 39684 5838 39740
rect 5838 39684 5842 39740
rect 5778 39680 5842 39684
rect 5858 39740 5922 39744
rect 5858 39684 5862 39740
rect 5862 39684 5918 39740
rect 5918 39684 5922 39740
rect 5858 39680 5922 39684
rect 5938 39740 6002 39744
rect 5938 39684 5942 39740
rect 5942 39684 5998 39740
rect 5998 39684 6002 39740
rect 5938 39680 6002 39684
rect 6018 39740 6082 39744
rect 6018 39684 6022 39740
rect 6022 39684 6078 39740
rect 6078 39684 6082 39740
rect 6018 39680 6082 39684
rect 2882 39196 2946 39200
rect 2882 39140 2886 39196
rect 2886 39140 2942 39196
rect 2942 39140 2946 39196
rect 2882 39136 2946 39140
rect 2962 39196 3026 39200
rect 2962 39140 2966 39196
rect 2966 39140 3022 39196
rect 3022 39140 3026 39196
rect 2962 39136 3026 39140
rect 3042 39196 3106 39200
rect 3042 39140 3046 39196
rect 3046 39140 3102 39196
rect 3102 39140 3106 39196
rect 3042 39136 3106 39140
rect 3122 39196 3186 39200
rect 3122 39140 3126 39196
rect 3126 39140 3182 39196
rect 3182 39140 3186 39196
rect 3122 39136 3186 39140
rect 4813 39196 4877 39200
rect 4813 39140 4817 39196
rect 4817 39140 4873 39196
rect 4873 39140 4877 39196
rect 4813 39136 4877 39140
rect 4893 39196 4957 39200
rect 4893 39140 4897 39196
rect 4897 39140 4953 39196
rect 4953 39140 4957 39196
rect 4893 39136 4957 39140
rect 4973 39196 5037 39200
rect 4973 39140 4977 39196
rect 4977 39140 5033 39196
rect 5033 39140 5037 39196
rect 4973 39136 5037 39140
rect 5053 39196 5117 39200
rect 5053 39140 5057 39196
rect 5057 39140 5113 39196
rect 5113 39140 5117 39196
rect 5053 39136 5117 39140
rect 2636 38932 2700 38996
rect 5580 38932 5644 38996
rect 2636 38660 2700 38724
rect 1917 38652 1981 38656
rect 1917 38596 1921 38652
rect 1921 38596 1977 38652
rect 1977 38596 1981 38652
rect 1917 38592 1981 38596
rect 1997 38652 2061 38656
rect 1997 38596 2001 38652
rect 2001 38596 2057 38652
rect 2057 38596 2061 38652
rect 1997 38592 2061 38596
rect 2077 38652 2141 38656
rect 2077 38596 2081 38652
rect 2081 38596 2137 38652
rect 2137 38596 2141 38652
rect 2077 38592 2141 38596
rect 2157 38652 2221 38656
rect 2157 38596 2161 38652
rect 2161 38596 2217 38652
rect 2217 38596 2221 38652
rect 2157 38592 2221 38596
rect 2452 38524 2516 38588
rect 3848 38652 3912 38656
rect 3848 38596 3852 38652
rect 3852 38596 3908 38652
rect 3908 38596 3912 38652
rect 3848 38592 3912 38596
rect 3928 38652 3992 38656
rect 3928 38596 3932 38652
rect 3932 38596 3988 38652
rect 3988 38596 3992 38652
rect 3928 38592 3992 38596
rect 4008 38652 4072 38656
rect 4008 38596 4012 38652
rect 4012 38596 4068 38652
rect 4068 38596 4072 38652
rect 4008 38592 4072 38596
rect 4088 38652 4152 38656
rect 4088 38596 4092 38652
rect 4092 38596 4148 38652
rect 4148 38596 4152 38652
rect 4088 38592 4152 38596
rect 5778 38652 5842 38656
rect 5778 38596 5782 38652
rect 5782 38596 5838 38652
rect 5838 38596 5842 38652
rect 5778 38592 5842 38596
rect 5858 38652 5922 38656
rect 5858 38596 5862 38652
rect 5862 38596 5918 38652
rect 5918 38596 5922 38652
rect 5858 38592 5922 38596
rect 5938 38652 6002 38656
rect 5938 38596 5942 38652
rect 5942 38596 5998 38652
rect 5998 38596 6002 38652
rect 5938 38592 6002 38596
rect 6018 38652 6082 38656
rect 6018 38596 6022 38652
rect 6022 38596 6078 38652
rect 6078 38596 6082 38652
rect 6018 38592 6082 38596
rect 3372 38252 3436 38316
rect 2882 38108 2946 38112
rect 2882 38052 2886 38108
rect 2886 38052 2942 38108
rect 2942 38052 2946 38108
rect 2882 38048 2946 38052
rect 2962 38108 3026 38112
rect 2962 38052 2966 38108
rect 2966 38052 3022 38108
rect 3022 38052 3026 38108
rect 2962 38048 3026 38052
rect 3042 38108 3106 38112
rect 3042 38052 3046 38108
rect 3046 38052 3102 38108
rect 3102 38052 3106 38108
rect 3042 38048 3106 38052
rect 3122 38108 3186 38112
rect 3122 38052 3126 38108
rect 3126 38052 3182 38108
rect 3182 38052 3186 38108
rect 3122 38048 3186 38052
rect 4813 38108 4877 38112
rect 4813 38052 4817 38108
rect 4817 38052 4873 38108
rect 4873 38052 4877 38108
rect 4813 38048 4877 38052
rect 4893 38108 4957 38112
rect 4893 38052 4897 38108
rect 4897 38052 4953 38108
rect 4953 38052 4957 38108
rect 4893 38048 4957 38052
rect 4973 38108 5037 38112
rect 4973 38052 4977 38108
rect 4977 38052 5033 38108
rect 5033 38052 5037 38108
rect 4973 38048 5037 38052
rect 5053 38108 5117 38112
rect 5053 38052 5057 38108
rect 5057 38052 5113 38108
rect 5113 38052 5117 38108
rect 5053 38048 5117 38052
rect 1716 37844 1780 37908
rect 1917 37564 1981 37568
rect 1917 37508 1921 37564
rect 1921 37508 1977 37564
rect 1977 37508 1981 37564
rect 1917 37504 1981 37508
rect 1997 37564 2061 37568
rect 1997 37508 2001 37564
rect 2001 37508 2057 37564
rect 2057 37508 2061 37564
rect 1997 37504 2061 37508
rect 2077 37564 2141 37568
rect 2077 37508 2081 37564
rect 2081 37508 2137 37564
rect 2137 37508 2141 37564
rect 2077 37504 2141 37508
rect 2157 37564 2221 37568
rect 2157 37508 2161 37564
rect 2161 37508 2217 37564
rect 2217 37508 2221 37564
rect 2157 37504 2221 37508
rect 3848 37564 3912 37568
rect 3848 37508 3852 37564
rect 3852 37508 3908 37564
rect 3908 37508 3912 37564
rect 3848 37504 3912 37508
rect 3928 37564 3992 37568
rect 3928 37508 3932 37564
rect 3932 37508 3988 37564
rect 3988 37508 3992 37564
rect 3928 37504 3992 37508
rect 4008 37564 4072 37568
rect 4008 37508 4012 37564
rect 4012 37508 4068 37564
rect 4068 37508 4072 37564
rect 4008 37504 4072 37508
rect 4088 37564 4152 37568
rect 4088 37508 4092 37564
rect 4092 37508 4148 37564
rect 4148 37508 4152 37564
rect 4088 37504 4152 37508
rect 5778 37564 5842 37568
rect 5778 37508 5782 37564
rect 5782 37508 5838 37564
rect 5838 37508 5842 37564
rect 5778 37504 5842 37508
rect 5858 37564 5922 37568
rect 5858 37508 5862 37564
rect 5862 37508 5918 37564
rect 5918 37508 5922 37564
rect 5858 37504 5922 37508
rect 5938 37564 6002 37568
rect 5938 37508 5942 37564
rect 5942 37508 5998 37564
rect 5998 37508 6002 37564
rect 5938 37504 6002 37508
rect 6018 37564 6082 37568
rect 6018 37508 6022 37564
rect 6022 37508 6078 37564
rect 6078 37508 6082 37564
rect 6018 37504 6082 37508
rect 2882 37020 2946 37024
rect 2882 36964 2886 37020
rect 2886 36964 2942 37020
rect 2942 36964 2946 37020
rect 2882 36960 2946 36964
rect 2962 37020 3026 37024
rect 2962 36964 2966 37020
rect 2966 36964 3022 37020
rect 3022 36964 3026 37020
rect 2962 36960 3026 36964
rect 3042 37020 3106 37024
rect 3042 36964 3046 37020
rect 3046 36964 3102 37020
rect 3102 36964 3106 37020
rect 3042 36960 3106 36964
rect 3122 37020 3186 37024
rect 3122 36964 3126 37020
rect 3126 36964 3182 37020
rect 3182 36964 3186 37020
rect 3122 36960 3186 36964
rect 4813 37020 4877 37024
rect 4813 36964 4817 37020
rect 4817 36964 4873 37020
rect 4873 36964 4877 37020
rect 4813 36960 4877 36964
rect 4893 37020 4957 37024
rect 4893 36964 4897 37020
rect 4897 36964 4953 37020
rect 4953 36964 4957 37020
rect 4893 36960 4957 36964
rect 4973 37020 5037 37024
rect 4973 36964 4977 37020
rect 4977 36964 5033 37020
rect 5033 36964 5037 37020
rect 4973 36960 5037 36964
rect 5053 37020 5117 37024
rect 5053 36964 5057 37020
rect 5057 36964 5113 37020
rect 5113 36964 5117 37020
rect 5053 36960 5117 36964
rect 2636 36952 2700 36956
rect 2636 36896 2686 36952
rect 2686 36896 2700 36952
rect 2636 36892 2700 36896
rect 1917 36476 1981 36480
rect 1917 36420 1921 36476
rect 1921 36420 1977 36476
rect 1977 36420 1981 36476
rect 1917 36416 1981 36420
rect 1997 36476 2061 36480
rect 1997 36420 2001 36476
rect 2001 36420 2057 36476
rect 2057 36420 2061 36476
rect 1997 36416 2061 36420
rect 2077 36476 2141 36480
rect 2077 36420 2081 36476
rect 2081 36420 2137 36476
rect 2137 36420 2141 36476
rect 2077 36416 2141 36420
rect 2157 36476 2221 36480
rect 2157 36420 2161 36476
rect 2161 36420 2217 36476
rect 2217 36420 2221 36476
rect 2157 36416 2221 36420
rect 3848 36476 3912 36480
rect 3848 36420 3852 36476
rect 3852 36420 3908 36476
rect 3908 36420 3912 36476
rect 3848 36416 3912 36420
rect 3928 36476 3992 36480
rect 3928 36420 3932 36476
rect 3932 36420 3988 36476
rect 3988 36420 3992 36476
rect 3928 36416 3992 36420
rect 4008 36476 4072 36480
rect 4008 36420 4012 36476
rect 4012 36420 4068 36476
rect 4068 36420 4072 36476
rect 4008 36416 4072 36420
rect 4088 36476 4152 36480
rect 4088 36420 4092 36476
rect 4092 36420 4148 36476
rect 4148 36420 4152 36476
rect 4088 36416 4152 36420
rect 5778 36476 5842 36480
rect 5778 36420 5782 36476
rect 5782 36420 5838 36476
rect 5838 36420 5842 36476
rect 5778 36416 5842 36420
rect 5858 36476 5922 36480
rect 5858 36420 5862 36476
rect 5862 36420 5918 36476
rect 5918 36420 5922 36476
rect 5858 36416 5922 36420
rect 5938 36476 6002 36480
rect 5938 36420 5942 36476
rect 5942 36420 5998 36476
rect 5998 36420 6002 36476
rect 5938 36416 6002 36420
rect 6018 36476 6082 36480
rect 6018 36420 6022 36476
rect 6022 36420 6078 36476
rect 6078 36420 6082 36476
rect 6018 36416 6082 36420
rect 2882 35932 2946 35936
rect 2882 35876 2886 35932
rect 2886 35876 2942 35932
rect 2942 35876 2946 35932
rect 2882 35872 2946 35876
rect 2962 35932 3026 35936
rect 2962 35876 2966 35932
rect 2966 35876 3022 35932
rect 3022 35876 3026 35932
rect 2962 35872 3026 35876
rect 3042 35932 3106 35936
rect 3042 35876 3046 35932
rect 3046 35876 3102 35932
rect 3102 35876 3106 35932
rect 3042 35872 3106 35876
rect 3122 35932 3186 35936
rect 3122 35876 3126 35932
rect 3126 35876 3182 35932
rect 3182 35876 3186 35932
rect 3122 35872 3186 35876
rect 4813 35932 4877 35936
rect 4813 35876 4817 35932
rect 4817 35876 4873 35932
rect 4873 35876 4877 35932
rect 4813 35872 4877 35876
rect 4893 35932 4957 35936
rect 4893 35876 4897 35932
rect 4897 35876 4953 35932
rect 4953 35876 4957 35932
rect 4893 35872 4957 35876
rect 4973 35932 5037 35936
rect 4973 35876 4977 35932
rect 4977 35876 5033 35932
rect 5033 35876 5037 35932
rect 4973 35872 5037 35876
rect 5053 35932 5117 35936
rect 5053 35876 5057 35932
rect 5057 35876 5113 35932
rect 5113 35876 5117 35932
rect 5053 35872 5117 35876
rect 1917 35388 1981 35392
rect 1917 35332 1921 35388
rect 1921 35332 1977 35388
rect 1977 35332 1981 35388
rect 1917 35328 1981 35332
rect 1997 35388 2061 35392
rect 1997 35332 2001 35388
rect 2001 35332 2057 35388
rect 2057 35332 2061 35388
rect 1997 35328 2061 35332
rect 2077 35388 2141 35392
rect 2077 35332 2081 35388
rect 2081 35332 2137 35388
rect 2137 35332 2141 35388
rect 2077 35328 2141 35332
rect 2157 35388 2221 35392
rect 2157 35332 2161 35388
rect 2161 35332 2217 35388
rect 2217 35332 2221 35388
rect 2157 35328 2221 35332
rect 3848 35388 3912 35392
rect 3848 35332 3852 35388
rect 3852 35332 3908 35388
rect 3908 35332 3912 35388
rect 3848 35328 3912 35332
rect 3928 35388 3992 35392
rect 3928 35332 3932 35388
rect 3932 35332 3988 35388
rect 3988 35332 3992 35388
rect 3928 35328 3992 35332
rect 4008 35388 4072 35392
rect 4008 35332 4012 35388
rect 4012 35332 4068 35388
rect 4068 35332 4072 35388
rect 4008 35328 4072 35332
rect 4088 35388 4152 35392
rect 4088 35332 4092 35388
rect 4092 35332 4148 35388
rect 4148 35332 4152 35388
rect 4088 35328 4152 35332
rect 5778 35388 5842 35392
rect 5778 35332 5782 35388
rect 5782 35332 5838 35388
rect 5838 35332 5842 35388
rect 5778 35328 5842 35332
rect 5858 35388 5922 35392
rect 5858 35332 5862 35388
rect 5862 35332 5918 35388
rect 5918 35332 5922 35388
rect 5858 35328 5922 35332
rect 5938 35388 6002 35392
rect 5938 35332 5942 35388
rect 5942 35332 5998 35388
rect 5998 35332 6002 35388
rect 5938 35328 6002 35332
rect 6018 35388 6082 35392
rect 6018 35332 6022 35388
rect 6022 35332 6078 35388
rect 6078 35332 6082 35388
rect 6018 35328 6082 35332
rect 2882 34844 2946 34848
rect 2882 34788 2886 34844
rect 2886 34788 2942 34844
rect 2942 34788 2946 34844
rect 2882 34784 2946 34788
rect 2962 34844 3026 34848
rect 2962 34788 2966 34844
rect 2966 34788 3022 34844
rect 3022 34788 3026 34844
rect 2962 34784 3026 34788
rect 3042 34844 3106 34848
rect 3042 34788 3046 34844
rect 3046 34788 3102 34844
rect 3102 34788 3106 34844
rect 3042 34784 3106 34788
rect 3122 34844 3186 34848
rect 3122 34788 3126 34844
rect 3126 34788 3182 34844
rect 3182 34788 3186 34844
rect 3122 34784 3186 34788
rect 4813 34844 4877 34848
rect 4813 34788 4817 34844
rect 4817 34788 4873 34844
rect 4873 34788 4877 34844
rect 4813 34784 4877 34788
rect 4893 34844 4957 34848
rect 4893 34788 4897 34844
rect 4897 34788 4953 34844
rect 4953 34788 4957 34844
rect 4893 34784 4957 34788
rect 4973 34844 5037 34848
rect 4973 34788 4977 34844
rect 4977 34788 5033 34844
rect 5033 34788 5037 34844
rect 4973 34784 5037 34788
rect 5053 34844 5117 34848
rect 5053 34788 5057 34844
rect 5057 34788 5113 34844
rect 5113 34788 5117 34844
rect 5053 34784 5117 34788
rect 4476 34444 4540 34508
rect 1917 34300 1981 34304
rect 1917 34244 1921 34300
rect 1921 34244 1977 34300
rect 1977 34244 1981 34300
rect 1917 34240 1981 34244
rect 1997 34300 2061 34304
rect 1997 34244 2001 34300
rect 2001 34244 2057 34300
rect 2057 34244 2061 34300
rect 1997 34240 2061 34244
rect 2077 34300 2141 34304
rect 2077 34244 2081 34300
rect 2081 34244 2137 34300
rect 2137 34244 2141 34300
rect 2077 34240 2141 34244
rect 2157 34300 2221 34304
rect 2157 34244 2161 34300
rect 2161 34244 2217 34300
rect 2217 34244 2221 34300
rect 2157 34240 2221 34244
rect 3848 34300 3912 34304
rect 3848 34244 3852 34300
rect 3852 34244 3908 34300
rect 3908 34244 3912 34300
rect 3848 34240 3912 34244
rect 3928 34300 3992 34304
rect 3928 34244 3932 34300
rect 3932 34244 3988 34300
rect 3988 34244 3992 34300
rect 3928 34240 3992 34244
rect 4008 34300 4072 34304
rect 4008 34244 4012 34300
rect 4012 34244 4068 34300
rect 4068 34244 4072 34300
rect 4008 34240 4072 34244
rect 4088 34300 4152 34304
rect 4088 34244 4092 34300
rect 4092 34244 4148 34300
rect 4148 34244 4152 34300
rect 4088 34240 4152 34244
rect 5778 34300 5842 34304
rect 5778 34244 5782 34300
rect 5782 34244 5838 34300
rect 5838 34244 5842 34300
rect 5778 34240 5842 34244
rect 5858 34300 5922 34304
rect 5858 34244 5862 34300
rect 5862 34244 5918 34300
rect 5918 34244 5922 34300
rect 5858 34240 5922 34244
rect 5938 34300 6002 34304
rect 5938 34244 5942 34300
rect 5942 34244 5998 34300
rect 5998 34244 6002 34300
rect 5938 34240 6002 34244
rect 6018 34300 6082 34304
rect 6018 34244 6022 34300
rect 6022 34244 6078 34300
rect 6078 34244 6082 34300
rect 6018 34240 6082 34244
rect 2882 33756 2946 33760
rect 2882 33700 2886 33756
rect 2886 33700 2942 33756
rect 2942 33700 2946 33756
rect 2882 33696 2946 33700
rect 2962 33756 3026 33760
rect 2962 33700 2966 33756
rect 2966 33700 3022 33756
rect 3022 33700 3026 33756
rect 2962 33696 3026 33700
rect 3042 33756 3106 33760
rect 3042 33700 3046 33756
rect 3046 33700 3102 33756
rect 3102 33700 3106 33756
rect 3042 33696 3106 33700
rect 3122 33756 3186 33760
rect 3122 33700 3126 33756
rect 3126 33700 3182 33756
rect 3182 33700 3186 33756
rect 3122 33696 3186 33700
rect 4813 33756 4877 33760
rect 4813 33700 4817 33756
rect 4817 33700 4873 33756
rect 4873 33700 4877 33756
rect 4813 33696 4877 33700
rect 4893 33756 4957 33760
rect 4893 33700 4897 33756
rect 4897 33700 4953 33756
rect 4953 33700 4957 33756
rect 4893 33696 4957 33700
rect 4973 33756 5037 33760
rect 4973 33700 4977 33756
rect 4977 33700 5033 33756
rect 5033 33700 5037 33756
rect 4973 33696 5037 33700
rect 5053 33756 5117 33760
rect 5053 33700 5057 33756
rect 5057 33700 5113 33756
rect 5113 33700 5117 33756
rect 5053 33696 5117 33700
rect 1917 33212 1981 33216
rect 1917 33156 1921 33212
rect 1921 33156 1977 33212
rect 1977 33156 1981 33212
rect 1917 33152 1981 33156
rect 1997 33212 2061 33216
rect 1997 33156 2001 33212
rect 2001 33156 2057 33212
rect 2057 33156 2061 33212
rect 1997 33152 2061 33156
rect 2077 33212 2141 33216
rect 2077 33156 2081 33212
rect 2081 33156 2137 33212
rect 2137 33156 2141 33212
rect 2077 33152 2141 33156
rect 2157 33212 2221 33216
rect 2157 33156 2161 33212
rect 2161 33156 2217 33212
rect 2217 33156 2221 33212
rect 2157 33152 2221 33156
rect 3848 33212 3912 33216
rect 3848 33156 3852 33212
rect 3852 33156 3908 33212
rect 3908 33156 3912 33212
rect 3848 33152 3912 33156
rect 3928 33212 3992 33216
rect 3928 33156 3932 33212
rect 3932 33156 3988 33212
rect 3988 33156 3992 33212
rect 3928 33152 3992 33156
rect 4008 33212 4072 33216
rect 4008 33156 4012 33212
rect 4012 33156 4068 33212
rect 4068 33156 4072 33212
rect 4008 33152 4072 33156
rect 4088 33212 4152 33216
rect 4088 33156 4092 33212
rect 4092 33156 4148 33212
rect 4148 33156 4152 33212
rect 4088 33152 4152 33156
rect 5778 33212 5842 33216
rect 5778 33156 5782 33212
rect 5782 33156 5838 33212
rect 5838 33156 5842 33212
rect 5778 33152 5842 33156
rect 5858 33212 5922 33216
rect 5858 33156 5862 33212
rect 5862 33156 5918 33212
rect 5918 33156 5922 33212
rect 5858 33152 5922 33156
rect 5938 33212 6002 33216
rect 5938 33156 5942 33212
rect 5942 33156 5998 33212
rect 5998 33156 6002 33212
rect 5938 33152 6002 33156
rect 6018 33212 6082 33216
rect 6018 33156 6022 33212
rect 6022 33156 6078 33212
rect 6078 33156 6082 33212
rect 6018 33152 6082 33156
rect 4292 32812 4356 32876
rect 2882 32668 2946 32672
rect 2882 32612 2886 32668
rect 2886 32612 2942 32668
rect 2942 32612 2946 32668
rect 2882 32608 2946 32612
rect 2962 32668 3026 32672
rect 2962 32612 2966 32668
rect 2966 32612 3022 32668
rect 3022 32612 3026 32668
rect 2962 32608 3026 32612
rect 3042 32668 3106 32672
rect 3042 32612 3046 32668
rect 3046 32612 3102 32668
rect 3102 32612 3106 32668
rect 3042 32608 3106 32612
rect 3122 32668 3186 32672
rect 3122 32612 3126 32668
rect 3126 32612 3182 32668
rect 3182 32612 3186 32668
rect 3122 32608 3186 32612
rect 4813 32668 4877 32672
rect 4813 32612 4817 32668
rect 4817 32612 4873 32668
rect 4873 32612 4877 32668
rect 4813 32608 4877 32612
rect 4893 32668 4957 32672
rect 4893 32612 4897 32668
rect 4897 32612 4953 32668
rect 4953 32612 4957 32668
rect 4893 32608 4957 32612
rect 4973 32668 5037 32672
rect 4973 32612 4977 32668
rect 4977 32612 5033 32668
rect 5033 32612 5037 32668
rect 4973 32608 5037 32612
rect 5053 32668 5117 32672
rect 5053 32612 5057 32668
rect 5057 32612 5113 32668
rect 5113 32612 5117 32668
rect 5053 32608 5117 32612
rect 4660 32268 4724 32332
rect 1917 32124 1981 32128
rect 1917 32068 1921 32124
rect 1921 32068 1977 32124
rect 1977 32068 1981 32124
rect 1917 32064 1981 32068
rect 1997 32124 2061 32128
rect 1997 32068 2001 32124
rect 2001 32068 2057 32124
rect 2057 32068 2061 32124
rect 1997 32064 2061 32068
rect 2077 32124 2141 32128
rect 2077 32068 2081 32124
rect 2081 32068 2137 32124
rect 2137 32068 2141 32124
rect 2077 32064 2141 32068
rect 2157 32124 2221 32128
rect 2157 32068 2161 32124
rect 2161 32068 2217 32124
rect 2217 32068 2221 32124
rect 2157 32064 2221 32068
rect 3848 32124 3912 32128
rect 3848 32068 3852 32124
rect 3852 32068 3908 32124
rect 3908 32068 3912 32124
rect 3848 32064 3912 32068
rect 3928 32124 3992 32128
rect 3928 32068 3932 32124
rect 3932 32068 3988 32124
rect 3988 32068 3992 32124
rect 3928 32064 3992 32068
rect 4008 32124 4072 32128
rect 4008 32068 4012 32124
rect 4012 32068 4068 32124
rect 4068 32068 4072 32124
rect 4008 32064 4072 32068
rect 4088 32124 4152 32128
rect 4088 32068 4092 32124
rect 4092 32068 4148 32124
rect 4148 32068 4152 32124
rect 4088 32064 4152 32068
rect 5778 32124 5842 32128
rect 5778 32068 5782 32124
rect 5782 32068 5838 32124
rect 5838 32068 5842 32124
rect 5778 32064 5842 32068
rect 5858 32124 5922 32128
rect 5858 32068 5862 32124
rect 5862 32068 5918 32124
rect 5918 32068 5922 32124
rect 5858 32064 5922 32068
rect 5938 32124 6002 32128
rect 5938 32068 5942 32124
rect 5942 32068 5998 32124
rect 5998 32068 6002 32124
rect 5938 32064 6002 32068
rect 6018 32124 6082 32128
rect 6018 32068 6022 32124
rect 6022 32068 6078 32124
rect 6078 32068 6082 32124
rect 6018 32064 6082 32068
rect 3556 31724 3620 31788
rect 2882 31580 2946 31584
rect 2882 31524 2886 31580
rect 2886 31524 2942 31580
rect 2942 31524 2946 31580
rect 2882 31520 2946 31524
rect 2962 31580 3026 31584
rect 2962 31524 2966 31580
rect 2966 31524 3022 31580
rect 3022 31524 3026 31580
rect 2962 31520 3026 31524
rect 3042 31580 3106 31584
rect 3042 31524 3046 31580
rect 3046 31524 3102 31580
rect 3102 31524 3106 31580
rect 3042 31520 3106 31524
rect 3122 31580 3186 31584
rect 3122 31524 3126 31580
rect 3126 31524 3182 31580
rect 3182 31524 3186 31580
rect 3122 31520 3186 31524
rect 4813 31580 4877 31584
rect 4813 31524 4817 31580
rect 4817 31524 4873 31580
rect 4873 31524 4877 31580
rect 4813 31520 4877 31524
rect 4893 31580 4957 31584
rect 4893 31524 4897 31580
rect 4897 31524 4953 31580
rect 4953 31524 4957 31580
rect 4893 31520 4957 31524
rect 4973 31580 5037 31584
rect 4973 31524 4977 31580
rect 4977 31524 5033 31580
rect 5033 31524 5037 31580
rect 4973 31520 5037 31524
rect 5053 31580 5117 31584
rect 5053 31524 5057 31580
rect 5057 31524 5113 31580
rect 5113 31524 5117 31580
rect 5053 31520 5117 31524
rect 2452 31240 2516 31244
rect 2452 31184 2466 31240
rect 2466 31184 2516 31240
rect 2452 31180 2516 31184
rect 1917 31036 1981 31040
rect 1917 30980 1921 31036
rect 1921 30980 1977 31036
rect 1977 30980 1981 31036
rect 1917 30976 1981 30980
rect 1997 31036 2061 31040
rect 1997 30980 2001 31036
rect 2001 30980 2057 31036
rect 2057 30980 2061 31036
rect 1997 30976 2061 30980
rect 2077 31036 2141 31040
rect 2077 30980 2081 31036
rect 2081 30980 2137 31036
rect 2137 30980 2141 31036
rect 2077 30976 2141 30980
rect 2157 31036 2221 31040
rect 2157 30980 2161 31036
rect 2161 30980 2217 31036
rect 2217 30980 2221 31036
rect 2157 30976 2221 30980
rect 3848 31036 3912 31040
rect 3848 30980 3852 31036
rect 3852 30980 3908 31036
rect 3908 30980 3912 31036
rect 3848 30976 3912 30980
rect 3928 31036 3992 31040
rect 3928 30980 3932 31036
rect 3932 30980 3988 31036
rect 3988 30980 3992 31036
rect 3928 30976 3992 30980
rect 4008 31036 4072 31040
rect 4008 30980 4012 31036
rect 4012 30980 4068 31036
rect 4068 30980 4072 31036
rect 4008 30976 4072 30980
rect 4088 31036 4152 31040
rect 4088 30980 4092 31036
rect 4092 30980 4148 31036
rect 4148 30980 4152 31036
rect 4088 30976 4152 30980
rect 5778 31036 5842 31040
rect 5778 30980 5782 31036
rect 5782 30980 5838 31036
rect 5838 30980 5842 31036
rect 5778 30976 5842 30980
rect 5858 31036 5922 31040
rect 5858 30980 5862 31036
rect 5862 30980 5918 31036
rect 5918 30980 5922 31036
rect 5858 30976 5922 30980
rect 5938 31036 6002 31040
rect 5938 30980 5942 31036
rect 5942 30980 5998 31036
rect 5998 30980 6002 31036
rect 5938 30976 6002 30980
rect 6018 31036 6082 31040
rect 6018 30980 6022 31036
rect 6022 30980 6078 31036
rect 6078 30980 6082 31036
rect 6018 30976 6082 30980
rect 2882 30492 2946 30496
rect 2882 30436 2886 30492
rect 2886 30436 2942 30492
rect 2942 30436 2946 30492
rect 2882 30432 2946 30436
rect 2962 30492 3026 30496
rect 2962 30436 2966 30492
rect 2966 30436 3022 30492
rect 3022 30436 3026 30492
rect 2962 30432 3026 30436
rect 3042 30492 3106 30496
rect 3042 30436 3046 30492
rect 3046 30436 3102 30492
rect 3102 30436 3106 30492
rect 3042 30432 3106 30436
rect 3122 30492 3186 30496
rect 3122 30436 3126 30492
rect 3126 30436 3182 30492
rect 3182 30436 3186 30492
rect 3122 30432 3186 30436
rect 4813 30492 4877 30496
rect 4813 30436 4817 30492
rect 4817 30436 4873 30492
rect 4873 30436 4877 30492
rect 4813 30432 4877 30436
rect 4893 30492 4957 30496
rect 4893 30436 4897 30492
rect 4897 30436 4953 30492
rect 4953 30436 4957 30492
rect 4893 30432 4957 30436
rect 4973 30492 5037 30496
rect 4973 30436 4977 30492
rect 4977 30436 5033 30492
rect 5033 30436 5037 30492
rect 4973 30432 5037 30436
rect 5053 30492 5117 30496
rect 5053 30436 5057 30492
rect 5057 30436 5113 30492
rect 5113 30436 5117 30492
rect 5053 30432 5117 30436
rect 1917 29948 1981 29952
rect 1917 29892 1921 29948
rect 1921 29892 1977 29948
rect 1977 29892 1981 29948
rect 1917 29888 1981 29892
rect 1997 29948 2061 29952
rect 1997 29892 2001 29948
rect 2001 29892 2057 29948
rect 2057 29892 2061 29948
rect 1997 29888 2061 29892
rect 2077 29948 2141 29952
rect 2077 29892 2081 29948
rect 2081 29892 2137 29948
rect 2137 29892 2141 29948
rect 2077 29888 2141 29892
rect 2157 29948 2221 29952
rect 2157 29892 2161 29948
rect 2161 29892 2217 29948
rect 2217 29892 2221 29948
rect 2157 29888 2221 29892
rect 3848 29948 3912 29952
rect 3848 29892 3852 29948
rect 3852 29892 3908 29948
rect 3908 29892 3912 29948
rect 3848 29888 3912 29892
rect 3928 29948 3992 29952
rect 3928 29892 3932 29948
rect 3932 29892 3988 29948
rect 3988 29892 3992 29948
rect 3928 29888 3992 29892
rect 4008 29948 4072 29952
rect 4008 29892 4012 29948
rect 4012 29892 4068 29948
rect 4068 29892 4072 29948
rect 4008 29888 4072 29892
rect 4088 29948 4152 29952
rect 4088 29892 4092 29948
rect 4092 29892 4148 29948
rect 4148 29892 4152 29948
rect 4088 29888 4152 29892
rect 5778 29948 5842 29952
rect 5778 29892 5782 29948
rect 5782 29892 5838 29948
rect 5838 29892 5842 29948
rect 5778 29888 5842 29892
rect 5858 29948 5922 29952
rect 5858 29892 5862 29948
rect 5862 29892 5918 29948
rect 5918 29892 5922 29948
rect 5858 29888 5922 29892
rect 5938 29948 6002 29952
rect 5938 29892 5942 29948
rect 5942 29892 5998 29948
rect 5998 29892 6002 29948
rect 5938 29888 6002 29892
rect 6018 29948 6082 29952
rect 6018 29892 6022 29948
rect 6022 29892 6078 29948
rect 6078 29892 6082 29948
rect 6018 29888 6082 29892
rect 3372 29820 3436 29884
rect 2882 29404 2946 29408
rect 2882 29348 2886 29404
rect 2886 29348 2942 29404
rect 2942 29348 2946 29404
rect 2882 29344 2946 29348
rect 2962 29404 3026 29408
rect 2962 29348 2966 29404
rect 2966 29348 3022 29404
rect 3022 29348 3026 29404
rect 2962 29344 3026 29348
rect 3042 29404 3106 29408
rect 3042 29348 3046 29404
rect 3046 29348 3102 29404
rect 3102 29348 3106 29404
rect 3042 29344 3106 29348
rect 3122 29404 3186 29408
rect 3122 29348 3126 29404
rect 3126 29348 3182 29404
rect 3182 29348 3186 29404
rect 3122 29344 3186 29348
rect 4813 29404 4877 29408
rect 4813 29348 4817 29404
rect 4817 29348 4873 29404
rect 4873 29348 4877 29404
rect 4813 29344 4877 29348
rect 4893 29404 4957 29408
rect 4893 29348 4897 29404
rect 4897 29348 4953 29404
rect 4953 29348 4957 29404
rect 4893 29344 4957 29348
rect 4973 29404 5037 29408
rect 4973 29348 4977 29404
rect 4977 29348 5033 29404
rect 5033 29348 5037 29404
rect 4973 29344 5037 29348
rect 5053 29404 5117 29408
rect 5053 29348 5057 29404
rect 5057 29348 5113 29404
rect 5113 29348 5117 29404
rect 5053 29344 5117 29348
rect 1917 28860 1981 28864
rect 1917 28804 1921 28860
rect 1921 28804 1977 28860
rect 1977 28804 1981 28860
rect 1917 28800 1981 28804
rect 1997 28860 2061 28864
rect 1997 28804 2001 28860
rect 2001 28804 2057 28860
rect 2057 28804 2061 28860
rect 1997 28800 2061 28804
rect 2077 28860 2141 28864
rect 2077 28804 2081 28860
rect 2081 28804 2137 28860
rect 2137 28804 2141 28860
rect 2077 28800 2141 28804
rect 2157 28860 2221 28864
rect 2157 28804 2161 28860
rect 2161 28804 2217 28860
rect 2217 28804 2221 28860
rect 2157 28800 2221 28804
rect 3848 28860 3912 28864
rect 3848 28804 3852 28860
rect 3852 28804 3908 28860
rect 3908 28804 3912 28860
rect 3848 28800 3912 28804
rect 3928 28860 3992 28864
rect 3928 28804 3932 28860
rect 3932 28804 3988 28860
rect 3988 28804 3992 28860
rect 3928 28800 3992 28804
rect 4008 28860 4072 28864
rect 4008 28804 4012 28860
rect 4012 28804 4068 28860
rect 4068 28804 4072 28860
rect 4008 28800 4072 28804
rect 4088 28860 4152 28864
rect 4088 28804 4092 28860
rect 4092 28804 4148 28860
rect 4148 28804 4152 28860
rect 4088 28800 4152 28804
rect 5778 28860 5842 28864
rect 5778 28804 5782 28860
rect 5782 28804 5838 28860
rect 5838 28804 5842 28860
rect 5778 28800 5842 28804
rect 5858 28860 5922 28864
rect 5858 28804 5862 28860
rect 5862 28804 5918 28860
rect 5918 28804 5922 28860
rect 5858 28800 5922 28804
rect 5938 28860 6002 28864
rect 5938 28804 5942 28860
rect 5942 28804 5998 28860
rect 5998 28804 6002 28860
rect 5938 28800 6002 28804
rect 6018 28860 6082 28864
rect 6018 28804 6022 28860
rect 6022 28804 6078 28860
rect 6078 28804 6082 28860
rect 6018 28800 6082 28804
rect 2882 28316 2946 28320
rect 2882 28260 2886 28316
rect 2886 28260 2942 28316
rect 2942 28260 2946 28316
rect 2882 28256 2946 28260
rect 2962 28316 3026 28320
rect 2962 28260 2966 28316
rect 2966 28260 3022 28316
rect 3022 28260 3026 28316
rect 2962 28256 3026 28260
rect 3042 28316 3106 28320
rect 3042 28260 3046 28316
rect 3046 28260 3102 28316
rect 3102 28260 3106 28316
rect 3042 28256 3106 28260
rect 3122 28316 3186 28320
rect 3122 28260 3126 28316
rect 3126 28260 3182 28316
rect 3182 28260 3186 28316
rect 3122 28256 3186 28260
rect 4813 28316 4877 28320
rect 4813 28260 4817 28316
rect 4817 28260 4873 28316
rect 4873 28260 4877 28316
rect 4813 28256 4877 28260
rect 4893 28316 4957 28320
rect 4893 28260 4897 28316
rect 4897 28260 4953 28316
rect 4953 28260 4957 28316
rect 4893 28256 4957 28260
rect 4973 28316 5037 28320
rect 4973 28260 4977 28316
rect 4977 28260 5033 28316
rect 5033 28260 5037 28316
rect 4973 28256 5037 28260
rect 5053 28316 5117 28320
rect 5053 28260 5057 28316
rect 5057 28260 5113 28316
rect 5113 28260 5117 28316
rect 5053 28256 5117 28260
rect 1917 27772 1981 27776
rect 1917 27716 1921 27772
rect 1921 27716 1977 27772
rect 1977 27716 1981 27772
rect 1917 27712 1981 27716
rect 1997 27772 2061 27776
rect 1997 27716 2001 27772
rect 2001 27716 2057 27772
rect 2057 27716 2061 27772
rect 1997 27712 2061 27716
rect 2077 27772 2141 27776
rect 2077 27716 2081 27772
rect 2081 27716 2137 27772
rect 2137 27716 2141 27772
rect 2077 27712 2141 27716
rect 2157 27772 2221 27776
rect 2157 27716 2161 27772
rect 2161 27716 2217 27772
rect 2217 27716 2221 27772
rect 2157 27712 2221 27716
rect 3848 27772 3912 27776
rect 3848 27716 3852 27772
rect 3852 27716 3908 27772
rect 3908 27716 3912 27772
rect 3848 27712 3912 27716
rect 3928 27772 3992 27776
rect 3928 27716 3932 27772
rect 3932 27716 3988 27772
rect 3988 27716 3992 27772
rect 3928 27712 3992 27716
rect 4008 27772 4072 27776
rect 4008 27716 4012 27772
rect 4012 27716 4068 27772
rect 4068 27716 4072 27772
rect 4008 27712 4072 27716
rect 4088 27772 4152 27776
rect 4088 27716 4092 27772
rect 4092 27716 4148 27772
rect 4148 27716 4152 27772
rect 4088 27712 4152 27716
rect 5778 27772 5842 27776
rect 5778 27716 5782 27772
rect 5782 27716 5838 27772
rect 5838 27716 5842 27772
rect 5778 27712 5842 27716
rect 5858 27772 5922 27776
rect 5858 27716 5862 27772
rect 5862 27716 5918 27772
rect 5918 27716 5922 27772
rect 5858 27712 5922 27716
rect 5938 27772 6002 27776
rect 5938 27716 5942 27772
rect 5942 27716 5998 27772
rect 5998 27716 6002 27772
rect 5938 27712 6002 27716
rect 6018 27772 6082 27776
rect 6018 27716 6022 27772
rect 6022 27716 6078 27772
rect 6078 27716 6082 27772
rect 6018 27712 6082 27716
rect 2882 27228 2946 27232
rect 2882 27172 2886 27228
rect 2886 27172 2942 27228
rect 2942 27172 2946 27228
rect 2882 27168 2946 27172
rect 2962 27228 3026 27232
rect 2962 27172 2966 27228
rect 2966 27172 3022 27228
rect 3022 27172 3026 27228
rect 2962 27168 3026 27172
rect 3042 27228 3106 27232
rect 3042 27172 3046 27228
rect 3046 27172 3102 27228
rect 3102 27172 3106 27228
rect 3042 27168 3106 27172
rect 3122 27228 3186 27232
rect 3122 27172 3126 27228
rect 3126 27172 3182 27228
rect 3182 27172 3186 27228
rect 3122 27168 3186 27172
rect 4813 27228 4877 27232
rect 4813 27172 4817 27228
rect 4817 27172 4873 27228
rect 4873 27172 4877 27228
rect 4813 27168 4877 27172
rect 4893 27228 4957 27232
rect 4893 27172 4897 27228
rect 4897 27172 4953 27228
rect 4953 27172 4957 27228
rect 4893 27168 4957 27172
rect 4973 27228 5037 27232
rect 4973 27172 4977 27228
rect 4977 27172 5033 27228
rect 5033 27172 5037 27228
rect 4973 27168 5037 27172
rect 5053 27228 5117 27232
rect 5053 27172 5057 27228
rect 5057 27172 5113 27228
rect 5113 27172 5117 27228
rect 5053 27168 5117 27172
rect 1917 26684 1981 26688
rect 1917 26628 1921 26684
rect 1921 26628 1977 26684
rect 1977 26628 1981 26684
rect 1917 26624 1981 26628
rect 1997 26684 2061 26688
rect 1997 26628 2001 26684
rect 2001 26628 2057 26684
rect 2057 26628 2061 26684
rect 1997 26624 2061 26628
rect 2077 26684 2141 26688
rect 2077 26628 2081 26684
rect 2081 26628 2137 26684
rect 2137 26628 2141 26684
rect 2077 26624 2141 26628
rect 2157 26684 2221 26688
rect 2157 26628 2161 26684
rect 2161 26628 2217 26684
rect 2217 26628 2221 26684
rect 2157 26624 2221 26628
rect 3848 26684 3912 26688
rect 3848 26628 3852 26684
rect 3852 26628 3908 26684
rect 3908 26628 3912 26684
rect 3848 26624 3912 26628
rect 3928 26684 3992 26688
rect 3928 26628 3932 26684
rect 3932 26628 3988 26684
rect 3988 26628 3992 26684
rect 3928 26624 3992 26628
rect 4008 26684 4072 26688
rect 4008 26628 4012 26684
rect 4012 26628 4068 26684
rect 4068 26628 4072 26684
rect 4008 26624 4072 26628
rect 4088 26684 4152 26688
rect 4088 26628 4092 26684
rect 4092 26628 4148 26684
rect 4148 26628 4152 26684
rect 4088 26624 4152 26628
rect 5778 26684 5842 26688
rect 5778 26628 5782 26684
rect 5782 26628 5838 26684
rect 5838 26628 5842 26684
rect 5778 26624 5842 26628
rect 5858 26684 5922 26688
rect 5858 26628 5862 26684
rect 5862 26628 5918 26684
rect 5918 26628 5922 26684
rect 5858 26624 5922 26628
rect 5938 26684 6002 26688
rect 5938 26628 5942 26684
rect 5942 26628 5998 26684
rect 5998 26628 6002 26684
rect 5938 26624 6002 26628
rect 6018 26684 6082 26688
rect 6018 26628 6022 26684
rect 6022 26628 6078 26684
rect 6078 26628 6082 26684
rect 6018 26624 6082 26628
rect 2882 26140 2946 26144
rect 2882 26084 2886 26140
rect 2886 26084 2942 26140
rect 2942 26084 2946 26140
rect 2882 26080 2946 26084
rect 2962 26140 3026 26144
rect 2962 26084 2966 26140
rect 2966 26084 3022 26140
rect 3022 26084 3026 26140
rect 2962 26080 3026 26084
rect 3042 26140 3106 26144
rect 3042 26084 3046 26140
rect 3046 26084 3102 26140
rect 3102 26084 3106 26140
rect 3042 26080 3106 26084
rect 3122 26140 3186 26144
rect 3122 26084 3126 26140
rect 3126 26084 3182 26140
rect 3182 26084 3186 26140
rect 3122 26080 3186 26084
rect 4813 26140 4877 26144
rect 4813 26084 4817 26140
rect 4817 26084 4873 26140
rect 4873 26084 4877 26140
rect 4813 26080 4877 26084
rect 4893 26140 4957 26144
rect 4893 26084 4897 26140
rect 4897 26084 4953 26140
rect 4953 26084 4957 26140
rect 4893 26080 4957 26084
rect 4973 26140 5037 26144
rect 4973 26084 4977 26140
rect 4977 26084 5033 26140
rect 5033 26084 5037 26140
rect 4973 26080 5037 26084
rect 5053 26140 5117 26144
rect 5053 26084 5057 26140
rect 5057 26084 5113 26140
rect 5113 26084 5117 26140
rect 5053 26080 5117 26084
rect 1917 25596 1981 25600
rect 1917 25540 1921 25596
rect 1921 25540 1977 25596
rect 1977 25540 1981 25596
rect 1917 25536 1981 25540
rect 1997 25596 2061 25600
rect 1997 25540 2001 25596
rect 2001 25540 2057 25596
rect 2057 25540 2061 25596
rect 1997 25536 2061 25540
rect 2077 25596 2141 25600
rect 2077 25540 2081 25596
rect 2081 25540 2137 25596
rect 2137 25540 2141 25596
rect 2077 25536 2141 25540
rect 2157 25596 2221 25600
rect 2157 25540 2161 25596
rect 2161 25540 2217 25596
rect 2217 25540 2221 25596
rect 2157 25536 2221 25540
rect 3848 25596 3912 25600
rect 3848 25540 3852 25596
rect 3852 25540 3908 25596
rect 3908 25540 3912 25596
rect 3848 25536 3912 25540
rect 3928 25596 3992 25600
rect 3928 25540 3932 25596
rect 3932 25540 3988 25596
rect 3988 25540 3992 25596
rect 3928 25536 3992 25540
rect 4008 25596 4072 25600
rect 4008 25540 4012 25596
rect 4012 25540 4068 25596
rect 4068 25540 4072 25596
rect 4008 25536 4072 25540
rect 4088 25596 4152 25600
rect 4088 25540 4092 25596
rect 4092 25540 4148 25596
rect 4148 25540 4152 25596
rect 4088 25536 4152 25540
rect 5778 25596 5842 25600
rect 5778 25540 5782 25596
rect 5782 25540 5838 25596
rect 5838 25540 5842 25596
rect 5778 25536 5842 25540
rect 5858 25596 5922 25600
rect 5858 25540 5862 25596
rect 5862 25540 5918 25596
rect 5918 25540 5922 25596
rect 5858 25536 5922 25540
rect 5938 25596 6002 25600
rect 5938 25540 5942 25596
rect 5942 25540 5998 25596
rect 5998 25540 6002 25596
rect 5938 25536 6002 25540
rect 6018 25596 6082 25600
rect 6018 25540 6022 25596
rect 6022 25540 6078 25596
rect 6078 25540 6082 25596
rect 6018 25536 6082 25540
rect 2882 25052 2946 25056
rect 2882 24996 2886 25052
rect 2886 24996 2942 25052
rect 2942 24996 2946 25052
rect 2882 24992 2946 24996
rect 2962 25052 3026 25056
rect 2962 24996 2966 25052
rect 2966 24996 3022 25052
rect 3022 24996 3026 25052
rect 2962 24992 3026 24996
rect 3042 25052 3106 25056
rect 3042 24996 3046 25052
rect 3046 24996 3102 25052
rect 3102 24996 3106 25052
rect 3042 24992 3106 24996
rect 3122 25052 3186 25056
rect 3122 24996 3126 25052
rect 3126 24996 3182 25052
rect 3182 24996 3186 25052
rect 3122 24992 3186 24996
rect 4813 25052 4877 25056
rect 4813 24996 4817 25052
rect 4817 24996 4873 25052
rect 4873 24996 4877 25052
rect 4813 24992 4877 24996
rect 4893 25052 4957 25056
rect 4893 24996 4897 25052
rect 4897 24996 4953 25052
rect 4953 24996 4957 25052
rect 4893 24992 4957 24996
rect 4973 25052 5037 25056
rect 4973 24996 4977 25052
rect 4977 24996 5033 25052
rect 5033 24996 5037 25052
rect 4973 24992 5037 24996
rect 5053 25052 5117 25056
rect 5053 24996 5057 25052
rect 5057 24996 5113 25052
rect 5113 24996 5117 25052
rect 5053 24992 5117 24996
rect 1917 24508 1981 24512
rect 1917 24452 1921 24508
rect 1921 24452 1977 24508
rect 1977 24452 1981 24508
rect 1917 24448 1981 24452
rect 1997 24508 2061 24512
rect 1997 24452 2001 24508
rect 2001 24452 2057 24508
rect 2057 24452 2061 24508
rect 1997 24448 2061 24452
rect 2077 24508 2141 24512
rect 2077 24452 2081 24508
rect 2081 24452 2137 24508
rect 2137 24452 2141 24508
rect 2077 24448 2141 24452
rect 2157 24508 2221 24512
rect 2157 24452 2161 24508
rect 2161 24452 2217 24508
rect 2217 24452 2221 24508
rect 2157 24448 2221 24452
rect 3848 24508 3912 24512
rect 3848 24452 3852 24508
rect 3852 24452 3908 24508
rect 3908 24452 3912 24508
rect 3848 24448 3912 24452
rect 3928 24508 3992 24512
rect 3928 24452 3932 24508
rect 3932 24452 3988 24508
rect 3988 24452 3992 24508
rect 3928 24448 3992 24452
rect 4008 24508 4072 24512
rect 4008 24452 4012 24508
rect 4012 24452 4068 24508
rect 4068 24452 4072 24508
rect 4008 24448 4072 24452
rect 4088 24508 4152 24512
rect 4088 24452 4092 24508
rect 4092 24452 4148 24508
rect 4148 24452 4152 24508
rect 4088 24448 4152 24452
rect 5778 24508 5842 24512
rect 5778 24452 5782 24508
rect 5782 24452 5838 24508
rect 5838 24452 5842 24508
rect 5778 24448 5842 24452
rect 5858 24508 5922 24512
rect 5858 24452 5862 24508
rect 5862 24452 5918 24508
rect 5918 24452 5922 24508
rect 5858 24448 5922 24452
rect 5938 24508 6002 24512
rect 5938 24452 5942 24508
rect 5942 24452 5998 24508
rect 5998 24452 6002 24508
rect 5938 24448 6002 24452
rect 6018 24508 6082 24512
rect 6018 24452 6022 24508
rect 6022 24452 6078 24508
rect 6078 24452 6082 24508
rect 6018 24448 6082 24452
rect 2882 23964 2946 23968
rect 2882 23908 2886 23964
rect 2886 23908 2942 23964
rect 2942 23908 2946 23964
rect 2882 23904 2946 23908
rect 2962 23964 3026 23968
rect 2962 23908 2966 23964
rect 2966 23908 3022 23964
rect 3022 23908 3026 23964
rect 2962 23904 3026 23908
rect 3042 23964 3106 23968
rect 3042 23908 3046 23964
rect 3046 23908 3102 23964
rect 3102 23908 3106 23964
rect 3042 23904 3106 23908
rect 3122 23964 3186 23968
rect 3122 23908 3126 23964
rect 3126 23908 3182 23964
rect 3182 23908 3186 23964
rect 3122 23904 3186 23908
rect 4813 23964 4877 23968
rect 4813 23908 4817 23964
rect 4817 23908 4873 23964
rect 4873 23908 4877 23964
rect 4813 23904 4877 23908
rect 4893 23964 4957 23968
rect 4893 23908 4897 23964
rect 4897 23908 4953 23964
rect 4953 23908 4957 23964
rect 4893 23904 4957 23908
rect 4973 23964 5037 23968
rect 4973 23908 4977 23964
rect 4977 23908 5033 23964
rect 5033 23908 5037 23964
rect 4973 23904 5037 23908
rect 5053 23964 5117 23968
rect 5053 23908 5057 23964
rect 5057 23908 5113 23964
rect 5113 23908 5117 23964
rect 5053 23904 5117 23908
rect 1917 23420 1981 23424
rect 1917 23364 1921 23420
rect 1921 23364 1977 23420
rect 1977 23364 1981 23420
rect 1917 23360 1981 23364
rect 1997 23420 2061 23424
rect 1997 23364 2001 23420
rect 2001 23364 2057 23420
rect 2057 23364 2061 23420
rect 1997 23360 2061 23364
rect 2077 23420 2141 23424
rect 2077 23364 2081 23420
rect 2081 23364 2137 23420
rect 2137 23364 2141 23420
rect 2077 23360 2141 23364
rect 2157 23420 2221 23424
rect 2157 23364 2161 23420
rect 2161 23364 2217 23420
rect 2217 23364 2221 23420
rect 2157 23360 2221 23364
rect 3848 23420 3912 23424
rect 3848 23364 3852 23420
rect 3852 23364 3908 23420
rect 3908 23364 3912 23420
rect 3848 23360 3912 23364
rect 3928 23420 3992 23424
rect 3928 23364 3932 23420
rect 3932 23364 3988 23420
rect 3988 23364 3992 23420
rect 3928 23360 3992 23364
rect 4008 23420 4072 23424
rect 4008 23364 4012 23420
rect 4012 23364 4068 23420
rect 4068 23364 4072 23420
rect 4008 23360 4072 23364
rect 4088 23420 4152 23424
rect 4088 23364 4092 23420
rect 4092 23364 4148 23420
rect 4148 23364 4152 23420
rect 4088 23360 4152 23364
rect 5778 23420 5842 23424
rect 5778 23364 5782 23420
rect 5782 23364 5838 23420
rect 5838 23364 5842 23420
rect 5778 23360 5842 23364
rect 5858 23420 5922 23424
rect 5858 23364 5862 23420
rect 5862 23364 5918 23420
rect 5918 23364 5922 23420
rect 5858 23360 5922 23364
rect 5938 23420 6002 23424
rect 5938 23364 5942 23420
rect 5942 23364 5998 23420
rect 5998 23364 6002 23420
rect 5938 23360 6002 23364
rect 6018 23420 6082 23424
rect 6018 23364 6022 23420
rect 6022 23364 6078 23420
rect 6078 23364 6082 23420
rect 6018 23360 6082 23364
rect 2882 22876 2946 22880
rect 2882 22820 2886 22876
rect 2886 22820 2942 22876
rect 2942 22820 2946 22876
rect 2882 22816 2946 22820
rect 2962 22876 3026 22880
rect 2962 22820 2966 22876
rect 2966 22820 3022 22876
rect 3022 22820 3026 22876
rect 2962 22816 3026 22820
rect 3042 22876 3106 22880
rect 3042 22820 3046 22876
rect 3046 22820 3102 22876
rect 3102 22820 3106 22876
rect 3042 22816 3106 22820
rect 3122 22876 3186 22880
rect 3122 22820 3126 22876
rect 3126 22820 3182 22876
rect 3182 22820 3186 22876
rect 3122 22816 3186 22820
rect 4813 22876 4877 22880
rect 4813 22820 4817 22876
rect 4817 22820 4873 22876
rect 4873 22820 4877 22876
rect 4813 22816 4877 22820
rect 4893 22876 4957 22880
rect 4893 22820 4897 22876
rect 4897 22820 4953 22876
rect 4953 22820 4957 22876
rect 4893 22816 4957 22820
rect 4973 22876 5037 22880
rect 4973 22820 4977 22876
rect 4977 22820 5033 22876
rect 5033 22820 5037 22876
rect 4973 22816 5037 22820
rect 5053 22876 5117 22880
rect 5053 22820 5057 22876
rect 5057 22820 5113 22876
rect 5113 22820 5117 22876
rect 5053 22816 5117 22820
rect 1917 22332 1981 22336
rect 1917 22276 1921 22332
rect 1921 22276 1977 22332
rect 1977 22276 1981 22332
rect 1917 22272 1981 22276
rect 1997 22332 2061 22336
rect 1997 22276 2001 22332
rect 2001 22276 2057 22332
rect 2057 22276 2061 22332
rect 1997 22272 2061 22276
rect 2077 22332 2141 22336
rect 2077 22276 2081 22332
rect 2081 22276 2137 22332
rect 2137 22276 2141 22332
rect 2077 22272 2141 22276
rect 2157 22332 2221 22336
rect 2157 22276 2161 22332
rect 2161 22276 2217 22332
rect 2217 22276 2221 22332
rect 2157 22272 2221 22276
rect 3848 22332 3912 22336
rect 3848 22276 3852 22332
rect 3852 22276 3908 22332
rect 3908 22276 3912 22332
rect 3848 22272 3912 22276
rect 3928 22332 3992 22336
rect 3928 22276 3932 22332
rect 3932 22276 3988 22332
rect 3988 22276 3992 22332
rect 3928 22272 3992 22276
rect 4008 22332 4072 22336
rect 4008 22276 4012 22332
rect 4012 22276 4068 22332
rect 4068 22276 4072 22332
rect 4008 22272 4072 22276
rect 4088 22332 4152 22336
rect 4088 22276 4092 22332
rect 4092 22276 4148 22332
rect 4148 22276 4152 22332
rect 4088 22272 4152 22276
rect 5778 22332 5842 22336
rect 5778 22276 5782 22332
rect 5782 22276 5838 22332
rect 5838 22276 5842 22332
rect 5778 22272 5842 22276
rect 5858 22332 5922 22336
rect 5858 22276 5862 22332
rect 5862 22276 5918 22332
rect 5918 22276 5922 22332
rect 5858 22272 5922 22276
rect 5938 22332 6002 22336
rect 5938 22276 5942 22332
rect 5942 22276 5998 22332
rect 5998 22276 6002 22332
rect 5938 22272 6002 22276
rect 6018 22332 6082 22336
rect 6018 22276 6022 22332
rect 6022 22276 6078 22332
rect 6078 22276 6082 22332
rect 6018 22272 6082 22276
rect 2882 21788 2946 21792
rect 2882 21732 2886 21788
rect 2886 21732 2942 21788
rect 2942 21732 2946 21788
rect 2882 21728 2946 21732
rect 2962 21788 3026 21792
rect 2962 21732 2966 21788
rect 2966 21732 3022 21788
rect 3022 21732 3026 21788
rect 2962 21728 3026 21732
rect 3042 21788 3106 21792
rect 3042 21732 3046 21788
rect 3046 21732 3102 21788
rect 3102 21732 3106 21788
rect 3042 21728 3106 21732
rect 3122 21788 3186 21792
rect 3122 21732 3126 21788
rect 3126 21732 3182 21788
rect 3182 21732 3186 21788
rect 3122 21728 3186 21732
rect 4813 21788 4877 21792
rect 4813 21732 4817 21788
rect 4817 21732 4873 21788
rect 4873 21732 4877 21788
rect 4813 21728 4877 21732
rect 4893 21788 4957 21792
rect 4893 21732 4897 21788
rect 4897 21732 4953 21788
rect 4953 21732 4957 21788
rect 4893 21728 4957 21732
rect 4973 21788 5037 21792
rect 4973 21732 4977 21788
rect 4977 21732 5033 21788
rect 5033 21732 5037 21788
rect 4973 21728 5037 21732
rect 5053 21788 5117 21792
rect 5053 21732 5057 21788
rect 5057 21732 5113 21788
rect 5113 21732 5117 21788
rect 5053 21728 5117 21732
rect 1917 21244 1981 21248
rect 1917 21188 1921 21244
rect 1921 21188 1977 21244
rect 1977 21188 1981 21244
rect 1917 21184 1981 21188
rect 1997 21244 2061 21248
rect 1997 21188 2001 21244
rect 2001 21188 2057 21244
rect 2057 21188 2061 21244
rect 1997 21184 2061 21188
rect 2077 21244 2141 21248
rect 2077 21188 2081 21244
rect 2081 21188 2137 21244
rect 2137 21188 2141 21244
rect 2077 21184 2141 21188
rect 2157 21244 2221 21248
rect 2157 21188 2161 21244
rect 2161 21188 2217 21244
rect 2217 21188 2221 21244
rect 2157 21184 2221 21188
rect 3848 21244 3912 21248
rect 3848 21188 3852 21244
rect 3852 21188 3908 21244
rect 3908 21188 3912 21244
rect 3848 21184 3912 21188
rect 3928 21244 3992 21248
rect 3928 21188 3932 21244
rect 3932 21188 3988 21244
rect 3988 21188 3992 21244
rect 3928 21184 3992 21188
rect 4008 21244 4072 21248
rect 4008 21188 4012 21244
rect 4012 21188 4068 21244
rect 4068 21188 4072 21244
rect 4008 21184 4072 21188
rect 4088 21244 4152 21248
rect 4088 21188 4092 21244
rect 4092 21188 4148 21244
rect 4148 21188 4152 21244
rect 4088 21184 4152 21188
rect 5778 21244 5842 21248
rect 5778 21188 5782 21244
rect 5782 21188 5838 21244
rect 5838 21188 5842 21244
rect 5778 21184 5842 21188
rect 5858 21244 5922 21248
rect 5858 21188 5862 21244
rect 5862 21188 5918 21244
rect 5918 21188 5922 21244
rect 5858 21184 5922 21188
rect 5938 21244 6002 21248
rect 5938 21188 5942 21244
rect 5942 21188 5998 21244
rect 5998 21188 6002 21244
rect 5938 21184 6002 21188
rect 6018 21244 6082 21248
rect 6018 21188 6022 21244
rect 6022 21188 6078 21244
rect 6078 21188 6082 21244
rect 6018 21184 6082 21188
rect 2882 20700 2946 20704
rect 2882 20644 2886 20700
rect 2886 20644 2942 20700
rect 2942 20644 2946 20700
rect 2882 20640 2946 20644
rect 2962 20700 3026 20704
rect 2962 20644 2966 20700
rect 2966 20644 3022 20700
rect 3022 20644 3026 20700
rect 2962 20640 3026 20644
rect 3042 20700 3106 20704
rect 3042 20644 3046 20700
rect 3046 20644 3102 20700
rect 3102 20644 3106 20700
rect 3042 20640 3106 20644
rect 3122 20700 3186 20704
rect 3122 20644 3126 20700
rect 3126 20644 3182 20700
rect 3182 20644 3186 20700
rect 3122 20640 3186 20644
rect 4813 20700 4877 20704
rect 4813 20644 4817 20700
rect 4817 20644 4873 20700
rect 4873 20644 4877 20700
rect 4813 20640 4877 20644
rect 4893 20700 4957 20704
rect 4893 20644 4897 20700
rect 4897 20644 4953 20700
rect 4953 20644 4957 20700
rect 4893 20640 4957 20644
rect 4973 20700 5037 20704
rect 4973 20644 4977 20700
rect 4977 20644 5033 20700
rect 5033 20644 5037 20700
rect 4973 20640 5037 20644
rect 5053 20700 5117 20704
rect 5053 20644 5057 20700
rect 5057 20644 5113 20700
rect 5113 20644 5117 20700
rect 5053 20640 5117 20644
rect 1917 20156 1981 20160
rect 1917 20100 1921 20156
rect 1921 20100 1977 20156
rect 1977 20100 1981 20156
rect 1917 20096 1981 20100
rect 1997 20156 2061 20160
rect 1997 20100 2001 20156
rect 2001 20100 2057 20156
rect 2057 20100 2061 20156
rect 1997 20096 2061 20100
rect 2077 20156 2141 20160
rect 2077 20100 2081 20156
rect 2081 20100 2137 20156
rect 2137 20100 2141 20156
rect 2077 20096 2141 20100
rect 2157 20156 2221 20160
rect 2157 20100 2161 20156
rect 2161 20100 2217 20156
rect 2217 20100 2221 20156
rect 2157 20096 2221 20100
rect 3848 20156 3912 20160
rect 3848 20100 3852 20156
rect 3852 20100 3908 20156
rect 3908 20100 3912 20156
rect 3848 20096 3912 20100
rect 3928 20156 3992 20160
rect 3928 20100 3932 20156
rect 3932 20100 3988 20156
rect 3988 20100 3992 20156
rect 3928 20096 3992 20100
rect 4008 20156 4072 20160
rect 4008 20100 4012 20156
rect 4012 20100 4068 20156
rect 4068 20100 4072 20156
rect 4008 20096 4072 20100
rect 4088 20156 4152 20160
rect 4088 20100 4092 20156
rect 4092 20100 4148 20156
rect 4148 20100 4152 20156
rect 4088 20096 4152 20100
rect 5778 20156 5842 20160
rect 5778 20100 5782 20156
rect 5782 20100 5838 20156
rect 5838 20100 5842 20156
rect 5778 20096 5842 20100
rect 5858 20156 5922 20160
rect 5858 20100 5862 20156
rect 5862 20100 5918 20156
rect 5918 20100 5922 20156
rect 5858 20096 5922 20100
rect 5938 20156 6002 20160
rect 5938 20100 5942 20156
rect 5942 20100 5998 20156
rect 5998 20100 6002 20156
rect 5938 20096 6002 20100
rect 6018 20156 6082 20160
rect 6018 20100 6022 20156
rect 6022 20100 6078 20156
rect 6078 20100 6082 20156
rect 6018 20096 6082 20100
rect 2882 19612 2946 19616
rect 2882 19556 2886 19612
rect 2886 19556 2942 19612
rect 2942 19556 2946 19612
rect 2882 19552 2946 19556
rect 2962 19612 3026 19616
rect 2962 19556 2966 19612
rect 2966 19556 3022 19612
rect 3022 19556 3026 19612
rect 2962 19552 3026 19556
rect 3042 19612 3106 19616
rect 3042 19556 3046 19612
rect 3046 19556 3102 19612
rect 3102 19556 3106 19612
rect 3042 19552 3106 19556
rect 3122 19612 3186 19616
rect 3122 19556 3126 19612
rect 3126 19556 3182 19612
rect 3182 19556 3186 19612
rect 3122 19552 3186 19556
rect 4813 19612 4877 19616
rect 4813 19556 4817 19612
rect 4817 19556 4873 19612
rect 4873 19556 4877 19612
rect 4813 19552 4877 19556
rect 4893 19612 4957 19616
rect 4893 19556 4897 19612
rect 4897 19556 4953 19612
rect 4953 19556 4957 19612
rect 4893 19552 4957 19556
rect 4973 19612 5037 19616
rect 4973 19556 4977 19612
rect 4977 19556 5033 19612
rect 5033 19556 5037 19612
rect 4973 19552 5037 19556
rect 5053 19612 5117 19616
rect 5053 19556 5057 19612
rect 5057 19556 5113 19612
rect 5113 19556 5117 19612
rect 5053 19552 5117 19556
rect 1917 19068 1981 19072
rect 1917 19012 1921 19068
rect 1921 19012 1977 19068
rect 1977 19012 1981 19068
rect 1917 19008 1981 19012
rect 1997 19068 2061 19072
rect 1997 19012 2001 19068
rect 2001 19012 2057 19068
rect 2057 19012 2061 19068
rect 1997 19008 2061 19012
rect 2077 19068 2141 19072
rect 2077 19012 2081 19068
rect 2081 19012 2137 19068
rect 2137 19012 2141 19068
rect 2077 19008 2141 19012
rect 2157 19068 2221 19072
rect 2157 19012 2161 19068
rect 2161 19012 2217 19068
rect 2217 19012 2221 19068
rect 2157 19008 2221 19012
rect 3848 19068 3912 19072
rect 3848 19012 3852 19068
rect 3852 19012 3908 19068
rect 3908 19012 3912 19068
rect 3848 19008 3912 19012
rect 3928 19068 3992 19072
rect 3928 19012 3932 19068
rect 3932 19012 3988 19068
rect 3988 19012 3992 19068
rect 3928 19008 3992 19012
rect 4008 19068 4072 19072
rect 4008 19012 4012 19068
rect 4012 19012 4068 19068
rect 4068 19012 4072 19068
rect 4008 19008 4072 19012
rect 4088 19068 4152 19072
rect 4088 19012 4092 19068
rect 4092 19012 4148 19068
rect 4148 19012 4152 19068
rect 4088 19008 4152 19012
rect 5778 19068 5842 19072
rect 5778 19012 5782 19068
rect 5782 19012 5838 19068
rect 5838 19012 5842 19068
rect 5778 19008 5842 19012
rect 5858 19068 5922 19072
rect 5858 19012 5862 19068
rect 5862 19012 5918 19068
rect 5918 19012 5922 19068
rect 5858 19008 5922 19012
rect 5938 19068 6002 19072
rect 5938 19012 5942 19068
rect 5942 19012 5998 19068
rect 5998 19012 6002 19068
rect 5938 19008 6002 19012
rect 6018 19068 6082 19072
rect 6018 19012 6022 19068
rect 6022 19012 6078 19068
rect 6078 19012 6082 19068
rect 6018 19008 6082 19012
rect 2882 18524 2946 18528
rect 2882 18468 2886 18524
rect 2886 18468 2942 18524
rect 2942 18468 2946 18524
rect 2882 18464 2946 18468
rect 2962 18524 3026 18528
rect 2962 18468 2966 18524
rect 2966 18468 3022 18524
rect 3022 18468 3026 18524
rect 2962 18464 3026 18468
rect 3042 18524 3106 18528
rect 3042 18468 3046 18524
rect 3046 18468 3102 18524
rect 3102 18468 3106 18524
rect 3042 18464 3106 18468
rect 3122 18524 3186 18528
rect 3122 18468 3126 18524
rect 3126 18468 3182 18524
rect 3182 18468 3186 18524
rect 3122 18464 3186 18468
rect 4813 18524 4877 18528
rect 4813 18468 4817 18524
rect 4817 18468 4873 18524
rect 4873 18468 4877 18524
rect 4813 18464 4877 18468
rect 4893 18524 4957 18528
rect 4893 18468 4897 18524
rect 4897 18468 4953 18524
rect 4953 18468 4957 18524
rect 4893 18464 4957 18468
rect 4973 18524 5037 18528
rect 4973 18468 4977 18524
rect 4977 18468 5033 18524
rect 5033 18468 5037 18524
rect 4973 18464 5037 18468
rect 5053 18524 5117 18528
rect 5053 18468 5057 18524
rect 5057 18468 5113 18524
rect 5113 18468 5117 18524
rect 5053 18464 5117 18468
rect 1917 17980 1981 17984
rect 1917 17924 1921 17980
rect 1921 17924 1977 17980
rect 1977 17924 1981 17980
rect 1917 17920 1981 17924
rect 1997 17980 2061 17984
rect 1997 17924 2001 17980
rect 2001 17924 2057 17980
rect 2057 17924 2061 17980
rect 1997 17920 2061 17924
rect 2077 17980 2141 17984
rect 2077 17924 2081 17980
rect 2081 17924 2137 17980
rect 2137 17924 2141 17980
rect 2077 17920 2141 17924
rect 2157 17980 2221 17984
rect 2157 17924 2161 17980
rect 2161 17924 2217 17980
rect 2217 17924 2221 17980
rect 2157 17920 2221 17924
rect 3848 17980 3912 17984
rect 3848 17924 3852 17980
rect 3852 17924 3908 17980
rect 3908 17924 3912 17980
rect 3848 17920 3912 17924
rect 3928 17980 3992 17984
rect 3928 17924 3932 17980
rect 3932 17924 3988 17980
rect 3988 17924 3992 17980
rect 3928 17920 3992 17924
rect 4008 17980 4072 17984
rect 4008 17924 4012 17980
rect 4012 17924 4068 17980
rect 4068 17924 4072 17980
rect 4008 17920 4072 17924
rect 4088 17980 4152 17984
rect 4088 17924 4092 17980
rect 4092 17924 4148 17980
rect 4148 17924 4152 17980
rect 4088 17920 4152 17924
rect 5778 17980 5842 17984
rect 5778 17924 5782 17980
rect 5782 17924 5838 17980
rect 5838 17924 5842 17980
rect 5778 17920 5842 17924
rect 5858 17980 5922 17984
rect 5858 17924 5862 17980
rect 5862 17924 5918 17980
rect 5918 17924 5922 17980
rect 5858 17920 5922 17924
rect 5938 17980 6002 17984
rect 5938 17924 5942 17980
rect 5942 17924 5998 17980
rect 5998 17924 6002 17980
rect 5938 17920 6002 17924
rect 6018 17980 6082 17984
rect 6018 17924 6022 17980
rect 6022 17924 6078 17980
rect 6078 17924 6082 17980
rect 6018 17920 6082 17924
rect 2882 17436 2946 17440
rect 2882 17380 2886 17436
rect 2886 17380 2942 17436
rect 2942 17380 2946 17436
rect 2882 17376 2946 17380
rect 2962 17436 3026 17440
rect 2962 17380 2966 17436
rect 2966 17380 3022 17436
rect 3022 17380 3026 17436
rect 2962 17376 3026 17380
rect 3042 17436 3106 17440
rect 3042 17380 3046 17436
rect 3046 17380 3102 17436
rect 3102 17380 3106 17436
rect 3042 17376 3106 17380
rect 3122 17436 3186 17440
rect 3122 17380 3126 17436
rect 3126 17380 3182 17436
rect 3182 17380 3186 17436
rect 3122 17376 3186 17380
rect 4813 17436 4877 17440
rect 4813 17380 4817 17436
rect 4817 17380 4873 17436
rect 4873 17380 4877 17436
rect 4813 17376 4877 17380
rect 4893 17436 4957 17440
rect 4893 17380 4897 17436
rect 4897 17380 4953 17436
rect 4953 17380 4957 17436
rect 4893 17376 4957 17380
rect 4973 17436 5037 17440
rect 4973 17380 4977 17436
rect 4977 17380 5033 17436
rect 5033 17380 5037 17436
rect 4973 17376 5037 17380
rect 5053 17436 5117 17440
rect 5053 17380 5057 17436
rect 5057 17380 5113 17436
rect 5113 17380 5117 17436
rect 5053 17376 5117 17380
rect 1917 16892 1981 16896
rect 1917 16836 1921 16892
rect 1921 16836 1977 16892
rect 1977 16836 1981 16892
rect 1917 16832 1981 16836
rect 1997 16892 2061 16896
rect 1997 16836 2001 16892
rect 2001 16836 2057 16892
rect 2057 16836 2061 16892
rect 1997 16832 2061 16836
rect 2077 16892 2141 16896
rect 2077 16836 2081 16892
rect 2081 16836 2137 16892
rect 2137 16836 2141 16892
rect 2077 16832 2141 16836
rect 2157 16892 2221 16896
rect 2157 16836 2161 16892
rect 2161 16836 2217 16892
rect 2217 16836 2221 16892
rect 2157 16832 2221 16836
rect 3848 16892 3912 16896
rect 3848 16836 3852 16892
rect 3852 16836 3908 16892
rect 3908 16836 3912 16892
rect 3848 16832 3912 16836
rect 3928 16892 3992 16896
rect 3928 16836 3932 16892
rect 3932 16836 3988 16892
rect 3988 16836 3992 16892
rect 3928 16832 3992 16836
rect 4008 16892 4072 16896
rect 4008 16836 4012 16892
rect 4012 16836 4068 16892
rect 4068 16836 4072 16892
rect 4008 16832 4072 16836
rect 4088 16892 4152 16896
rect 4088 16836 4092 16892
rect 4092 16836 4148 16892
rect 4148 16836 4152 16892
rect 4088 16832 4152 16836
rect 5778 16892 5842 16896
rect 5778 16836 5782 16892
rect 5782 16836 5838 16892
rect 5838 16836 5842 16892
rect 5778 16832 5842 16836
rect 5858 16892 5922 16896
rect 5858 16836 5862 16892
rect 5862 16836 5918 16892
rect 5918 16836 5922 16892
rect 5858 16832 5922 16836
rect 5938 16892 6002 16896
rect 5938 16836 5942 16892
rect 5942 16836 5998 16892
rect 5998 16836 6002 16892
rect 5938 16832 6002 16836
rect 6018 16892 6082 16896
rect 6018 16836 6022 16892
rect 6022 16836 6078 16892
rect 6078 16836 6082 16892
rect 6018 16832 6082 16836
rect 2882 16348 2946 16352
rect 2882 16292 2886 16348
rect 2886 16292 2942 16348
rect 2942 16292 2946 16348
rect 2882 16288 2946 16292
rect 2962 16348 3026 16352
rect 2962 16292 2966 16348
rect 2966 16292 3022 16348
rect 3022 16292 3026 16348
rect 2962 16288 3026 16292
rect 3042 16348 3106 16352
rect 3042 16292 3046 16348
rect 3046 16292 3102 16348
rect 3102 16292 3106 16348
rect 3042 16288 3106 16292
rect 3122 16348 3186 16352
rect 3122 16292 3126 16348
rect 3126 16292 3182 16348
rect 3182 16292 3186 16348
rect 3122 16288 3186 16292
rect 4813 16348 4877 16352
rect 4813 16292 4817 16348
rect 4817 16292 4873 16348
rect 4873 16292 4877 16348
rect 4813 16288 4877 16292
rect 4893 16348 4957 16352
rect 4893 16292 4897 16348
rect 4897 16292 4953 16348
rect 4953 16292 4957 16348
rect 4893 16288 4957 16292
rect 4973 16348 5037 16352
rect 4973 16292 4977 16348
rect 4977 16292 5033 16348
rect 5033 16292 5037 16348
rect 4973 16288 5037 16292
rect 5053 16348 5117 16352
rect 5053 16292 5057 16348
rect 5057 16292 5113 16348
rect 5113 16292 5117 16348
rect 5053 16288 5117 16292
rect 1917 15804 1981 15808
rect 1917 15748 1921 15804
rect 1921 15748 1977 15804
rect 1977 15748 1981 15804
rect 1917 15744 1981 15748
rect 1997 15804 2061 15808
rect 1997 15748 2001 15804
rect 2001 15748 2057 15804
rect 2057 15748 2061 15804
rect 1997 15744 2061 15748
rect 2077 15804 2141 15808
rect 2077 15748 2081 15804
rect 2081 15748 2137 15804
rect 2137 15748 2141 15804
rect 2077 15744 2141 15748
rect 2157 15804 2221 15808
rect 2157 15748 2161 15804
rect 2161 15748 2217 15804
rect 2217 15748 2221 15804
rect 2157 15744 2221 15748
rect 3848 15804 3912 15808
rect 3848 15748 3852 15804
rect 3852 15748 3908 15804
rect 3908 15748 3912 15804
rect 3848 15744 3912 15748
rect 3928 15804 3992 15808
rect 3928 15748 3932 15804
rect 3932 15748 3988 15804
rect 3988 15748 3992 15804
rect 3928 15744 3992 15748
rect 4008 15804 4072 15808
rect 4008 15748 4012 15804
rect 4012 15748 4068 15804
rect 4068 15748 4072 15804
rect 4008 15744 4072 15748
rect 4088 15804 4152 15808
rect 4088 15748 4092 15804
rect 4092 15748 4148 15804
rect 4148 15748 4152 15804
rect 4088 15744 4152 15748
rect 5778 15804 5842 15808
rect 5778 15748 5782 15804
rect 5782 15748 5838 15804
rect 5838 15748 5842 15804
rect 5778 15744 5842 15748
rect 5858 15804 5922 15808
rect 5858 15748 5862 15804
rect 5862 15748 5918 15804
rect 5918 15748 5922 15804
rect 5858 15744 5922 15748
rect 5938 15804 6002 15808
rect 5938 15748 5942 15804
rect 5942 15748 5998 15804
rect 5998 15748 6002 15804
rect 5938 15744 6002 15748
rect 6018 15804 6082 15808
rect 6018 15748 6022 15804
rect 6022 15748 6078 15804
rect 6078 15748 6082 15804
rect 6018 15744 6082 15748
rect 2882 15260 2946 15264
rect 2882 15204 2886 15260
rect 2886 15204 2942 15260
rect 2942 15204 2946 15260
rect 2882 15200 2946 15204
rect 2962 15260 3026 15264
rect 2962 15204 2966 15260
rect 2966 15204 3022 15260
rect 3022 15204 3026 15260
rect 2962 15200 3026 15204
rect 3042 15260 3106 15264
rect 3042 15204 3046 15260
rect 3046 15204 3102 15260
rect 3102 15204 3106 15260
rect 3042 15200 3106 15204
rect 3122 15260 3186 15264
rect 3122 15204 3126 15260
rect 3126 15204 3182 15260
rect 3182 15204 3186 15260
rect 3122 15200 3186 15204
rect 4813 15260 4877 15264
rect 4813 15204 4817 15260
rect 4817 15204 4873 15260
rect 4873 15204 4877 15260
rect 4813 15200 4877 15204
rect 4893 15260 4957 15264
rect 4893 15204 4897 15260
rect 4897 15204 4953 15260
rect 4953 15204 4957 15260
rect 4893 15200 4957 15204
rect 4973 15260 5037 15264
rect 4973 15204 4977 15260
rect 4977 15204 5033 15260
rect 5033 15204 5037 15260
rect 4973 15200 5037 15204
rect 5053 15260 5117 15264
rect 5053 15204 5057 15260
rect 5057 15204 5113 15260
rect 5113 15204 5117 15260
rect 5053 15200 5117 15204
rect 1917 14716 1981 14720
rect 1917 14660 1921 14716
rect 1921 14660 1977 14716
rect 1977 14660 1981 14716
rect 1917 14656 1981 14660
rect 1997 14716 2061 14720
rect 1997 14660 2001 14716
rect 2001 14660 2057 14716
rect 2057 14660 2061 14716
rect 1997 14656 2061 14660
rect 2077 14716 2141 14720
rect 2077 14660 2081 14716
rect 2081 14660 2137 14716
rect 2137 14660 2141 14716
rect 2077 14656 2141 14660
rect 2157 14716 2221 14720
rect 2157 14660 2161 14716
rect 2161 14660 2217 14716
rect 2217 14660 2221 14716
rect 2157 14656 2221 14660
rect 3848 14716 3912 14720
rect 3848 14660 3852 14716
rect 3852 14660 3908 14716
rect 3908 14660 3912 14716
rect 3848 14656 3912 14660
rect 3928 14716 3992 14720
rect 3928 14660 3932 14716
rect 3932 14660 3988 14716
rect 3988 14660 3992 14716
rect 3928 14656 3992 14660
rect 4008 14716 4072 14720
rect 4008 14660 4012 14716
rect 4012 14660 4068 14716
rect 4068 14660 4072 14716
rect 4008 14656 4072 14660
rect 4088 14716 4152 14720
rect 4088 14660 4092 14716
rect 4092 14660 4148 14716
rect 4148 14660 4152 14716
rect 4088 14656 4152 14660
rect 5778 14716 5842 14720
rect 5778 14660 5782 14716
rect 5782 14660 5838 14716
rect 5838 14660 5842 14716
rect 5778 14656 5842 14660
rect 5858 14716 5922 14720
rect 5858 14660 5862 14716
rect 5862 14660 5918 14716
rect 5918 14660 5922 14716
rect 5858 14656 5922 14660
rect 5938 14716 6002 14720
rect 5938 14660 5942 14716
rect 5942 14660 5998 14716
rect 5998 14660 6002 14716
rect 5938 14656 6002 14660
rect 6018 14716 6082 14720
rect 6018 14660 6022 14716
rect 6022 14660 6078 14716
rect 6078 14660 6082 14716
rect 6018 14656 6082 14660
rect 2882 14172 2946 14176
rect 2882 14116 2886 14172
rect 2886 14116 2942 14172
rect 2942 14116 2946 14172
rect 2882 14112 2946 14116
rect 2962 14172 3026 14176
rect 2962 14116 2966 14172
rect 2966 14116 3022 14172
rect 3022 14116 3026 14172
rect 2962 14112 3026 14116
rect 3042 14172 3106 14176
rect 3042 14116 3046 14172
rect 3046 14116 3102 14172
rect 3102 14116 3106 14172
rect 3042 14112 3106 14116
rect 3122 14172 3186 14176
rect 3122 14116 3126 14172
rect 3126 14116 3182 14172
rect 3182 14116 3186 14172
rect 3122 14112 3186 14116
rect 4813 14172 4877 14176
rect 4813 14116 4817 14172
rect 4817 14116 4873 14172
rect 4873 14116 4877 14172
rect 4813 14112 4877 14116
rect 4893 14172 4957 14176
rect 4893 14116 4897 14172
rect 4897 14116 4953 14172
rect 4953 14116 4957 14172
rect 4893 14112 4957 14116
rect 4973 14172 5037 14176
rect 4973 14116 4977 14172
rect 4977 14116 5033 14172
rect 5033 14116 5037 14172
rect 4973 14112 5037 14116
rect 5053 14172 5117 14176
rect 5053 14116 5057 14172
rect 5057 14116 5113 14172
rect 5113 14116 5117 14172
rect 5053 14112 5117 14116
rect 1917 13628 1981 13632
rect 1917 13572 1921 13628
rect 1921 13572 1977 13628
rect 1977 13572 1981 13628
rect 1917 13568 1981 13572
rect 1997 13628 2061 13632
rect 1997 13572 2001 13628
rect 2001 13572 2057 13628
rect 2057 13572 2061 13628
rect 1997 13568 2061 13572
rect 2077 13628 2141 13632
rect 2077 13572 2081 13628
rect 2081 13572 2137 13628
rect 2137 13572 2141 13628
rect 2077 13568 2141 13572
rect 2157 13628 2221 13632
rect 2157 13572 2161 13628
rect 2161 13572 2217 13628
rect 2217 13572 2221 13628
rect 2157 13568 2221 13572
rect 3848 13628 3912 13632
rect 3848 13572 3852 13628
rect 3852 13572 3908 13628
rect 3908 13572 3912 13628
rect 3848 13568 3912 13572
rect 3928 13628 3992 13632
rect 3928 13572 3932 13628
rect 3932 13572 3988 13628
rect 3988 13572 3992 13628
rect 3928 13568 3992 13572
rect 4008 13628 4072 13632
rect 4008 13572 4012 13628
rect 4012 13572 4068 13628
rect 4068 13572 4072 13628
rect 4008 13568 4072 13572
rect 4088 13628 4152 13632
rect 4088 13572 4092 13628
rect 4092 13572 4148 13628
rect 4148 13572 4152 13628
rect 4088 13568 4152 13572
rect 5778 13628 5842 13632
rect 5778 13572 5782 13628
rect 5782 13572 5838 13628
rect 5838 13572 5842 13628
rect 5778 13568 5842 13572
rect 5858 13628 5922 13632
rect 5858 13572 5862 13628
rect 5862 13572 5918 13628
rect 5918 13572 5922 13628
rect 5858 13568 5922 13572
rect 5938 13628 6002 13632
rect 5938 13572 5942 13628
rect 5942 13572 5998 13628
rect 5998 13572 6002 13628
rect 5938 13568 6002 13572
rect 6018 13628 6082 13632
rect 6018 13572 6022 13628
rect 6022 13572 6078 13628
rect 6078 13572 6082 13628
rect 6018 13568 6082 13572
rect 2882 13084 2946 13088
rect 2882 13028 2886 13084
rect 2886 13028 2942 13084
rect 2942 13028 2946 13084
rect 2882 13024 2946 13028
rect 2962 13084 3026 13088
rect 2962 13028 2966 13084
rect 2966 13028 3022 13084
rect 3022 13028 3026 13084
rect 2962 13024 3026 13028
rect 3042 13084 3106 13088
rect 3042 13028 3046 13084
rect 3046 13028 3102 13084
rect 3102 13028 3106 13084
rect 3042 13024 3106 13028
rect 3122 13084 3186 13088
rect 3122 13028 3126 13084
rect 3126 13028 3182 13084
rect 3182 13028 3186 13084
rect 3122 13024 3186 13028
rect 4813 13084 4877 13088
rect 4813 13028 4817 13084
rect 4817 13028 4873 13084
rect 4873 13028 4877 13084
rect 4813 13024 4877 13028
rect 4893 13084 4957 13088
rect 4893 13028 4897 13084
rect 4897 13028 4953 13084
rect 4953 13028 4957 13084
rect 4893 13024 4957 13028
rect 4973 13084 5037 13088
rect 4973 13028 4977 13084
rect 4977 13028 5033 13084
rect 5033 13028 5037 13084
rect 4973 13024 5037 13028
rect 5053 13084 5117 13088
rect 5053 13028 5057 13084
rect 5057 13028 5113 13084
rect 5113 13028 5117 13084
rect 5053 13024 5117 13028
rect 1917 12540 1981 12544
rect 1917 12484 1921 12540
rect 1921 12484 1977 12540
rect 1977 12484 1981 12540
rect 1917 12480 1981 12484
rect 1997 12540 2061 12544
rect 1997 12484 2001 12540
rect 2001 12484 2057 12540
rect 2057 12484 2061 12540
rect 1997 12480 2061 12484
rect 2077 12540 2141 12544
rect 2077 12484 2081 12540
rect 2081 12484 2137 12540
rect 2137 12484 2141 12540
rect 2077 12480 2141 12484
rect 2157 12540 2221 12544
rect 2157 12484 2161 12540
rect 2161 12484 2217 12540
rect 2217 12484 2221 12540
rect 2157 12480 2221 12484
rect 3848 12540 3912 12544
rect 3848 12484 3852 12540
rect 3852 12484 3908 12540
rect 3908 12484 3912 12540
rect 3848 12480 3912 12484
rect 3928 12540 3992 12544
rect 3928 12484 3932 12540
rect 3932 12484 3988 12540
rect 3988 12484 3992 12540
rect 3928 12480 3992 12484
rect 4008 12540 4072 12544
rect 4008 12484 4012 12540
rect 4012 12484 4068 12540
rect 4068 12484 4072 12540
rect 4008 12480 4072 12484
rect 4088 12540 4152 12544
rect 4088 12484 4092 12540
rect 4092 12484 4148 12540
rect 4148 12484 4152 12540
rect 4088 12480 4152 12484
rect 5778 12540 5842 12544
rect 5778 12484 5782 12540
rect 5782 12484 5838 12540
rect 5838 12484 5842 12540
rect 5778 12480 5842 12484
rect 5858 12540 5922 12544
rect 5858 12484 5862 12540
rect 5862 12484 5918 12540
rect 5918 12484 5922 12540
rect 5858 12480 5922 12484
rect 5938 12540 6002 12544
rect 5938 12484 5942 12540
rect 5942 12484 5998 12540
rect 5998 12484 6002 12540
rect 5938 12480 6002 12484
rect 6018 12540 6082 12544
rect 6018 12484 6022 12540
rect 6022 12484 6078 12540
rect 6078 12484 6082 12540
rect 6018 12480 6082 12484
rect 2882 11996 2946 12000
rect 2882 11940 2886 11996
rect 2886 11940 2942 11996
rect 2942 11940 2946 11996
rect 2882 11936 2946 11940
rect 2962 11996 3026 12000
rect 2962 11940 2966 11996
rect 2966 11940 3022 11996
rect 3022 11940 3026 11996
rect 2962 11936 3026 11940
rect 3042 11996 3106 12000
rect 3042 11940 3046 11996
rect 3046 11940 3102 11996
rect 3102 11940 3106 11996
rect 3042 11936 3106 11940
rect 3122 11996 3186 12000
rect 3122 11940 3126 11996
rect 3126 11940 3182 11996
rect 3182 11940 3186 11996
rect 3122 11936 3186 11940
rect 4813 11996 4877 12000
rect 4813 11940 4817 11996
rect 4817 11940 4873 11996
rect 4873 11940 4877 11996
rect 4813 11936 4877 11940
rect 4893 11996 4957 12000
rect 4893 11940 4897 11996
rect 4897 11940 4953 11996
rect 4953 11940 4957 11996
rect 4893 11936 4957 11940
rect 4973 11996 5037 12000
rect 4973 11940 4977 11996
rect 4977 11940 5033 11996
rect 5033 11940 5037 11996
rect 4973 11936 5037 11940
rect 5053 11996 5117 12000
rect 5053 11940 5057 11996
rect 5057 11940 5113 11996
rect 5113 11940 5117 11996
rect 5053 11936 5117 11940
rect 1917 11452 1981 11456
rect 1917 11396 1921 11452
rect 1921 11396 1977 11452
rect 1977 11396 1981 11452
rect 1917 11392 1981 11396
rect 1997 11452 2061 11456
rect 1997 11396 2001 11452
rect 2001 11396 2057 11452
rect 2057 11396 2061 11452
rect 1997 11392 2061 11396
rect 2077 11452 2141 11456
rect 2077 11396 2081 11452
rect 2081 11396 2137 11452
rect 2137 11396 2141 11452
rect 2077 11392 2141 11396
rect 2157 11452 2221 11456
rect 2157 11396 2161 11452
rect 2161 11396 2217 11452
rect 2217 11396 2221 11452
rect 2157 11392 2221 11396
rect 3848 11452 3912 11456
rect 3848 11396 3852 11452
rect 3852 11396 3908 11452
rect 3908 11396 3912 11452
rect 3848 11392 3912 11396
rect 3928 11452 3992 11456
rect 3928 11396 3932 11452
rect 3932 11396 3988 11452
rect 3988 11396 3992 11452
rect 3928 11392 3992 11396
rect 4008 11452 4072 11456
rect 4008 11396 4012 11452
rect 4012 11396 4068 11452
rect 4068 11396 4072 11452
rect 4008 11392 4072 11396
rect 4088 11452 4152 11456
rect 4088 11396 4092 11452
rect 4092 11396 4148 11452
rect 4148 11396 4152 11452
rect 4088 11392 4152 11396
rect 5778 11452 5842 11456
rect 5778 11396 5782 11452
rect 5782 11396 5838 11452
rect 5838 11396 5842 11452
rect 5778 11392 5842 11396
rect 5858 11452 5922 11456
rect 5858 11396 5862 11452
rect 5862 11396 5918 11452
rect 5918 11396 5922 11452
rect 5858 11392 5922 11396
rect 5938 11452 6002 11456
rect 5938 11396 5942 11452
rect 5942 11396 5998 11452
rect 5998 11396 6002 11452
rect 5938 11392 6002 11396
rect 6018 11452 6082 11456
rect 6018 11396 6022 11452
rect 6022 11396 6078 11452
rect 6078 11396 6082 11452
rect 6018 11392 6082 11396
rect 2882 10908 2946 10912
rect 2882 10852 2886 10908
rect 2886 10852 2942 10908
rect 2942 10852 2946 10908
rect 2882 10848 2946 10852
rect 2962 10908 3026 10912
rect 2962 10852 2966 10908
rect 2966 10852 3022 10908
rect 3022 10852 3026 10908
rect 2962 10848 3026 10852
rect 3042 10908 3106 10912
rect 3042 10852 3046 10908
rect 3046 10852 3102 10908
rect 3102 10852 3106 10908
rect 3042 10848 3106 10852
rect 3122 10908 3186 10912
rect 3122 10852 3126 10908
rect 3126 10852 3182 10908
rect 3182 10852 3186 10908
rect 3122 10848 3186 10852
rect 4813 10908 4877 10912
rect 4813 10852 4817 10908
rect 4817 10852 4873 10908
rect 4873 10852 4877 10908
rect 4813 10848 4877 10852
rect 4893 10908 4957 10912
rect 4893 10852 4897 10908
rect 4897 10852 4953 10908
rect 4953 10852 4957 10908
rect 4893 10848 4957 10852
rect 4973 10908 5037 10912
rect 4973 10852 4977 10908
rect 4977 10852 5033 10908
rect 5033 10852 5037 10908
rect 4973 10848 5037 10852
rect 5053 10908 5117 10912
rect 5053 10852 5057 10908
rect 5057 10852 5113 10908
rect 5113 10852 5117 10908
rect 5053 10848 5117 10852
rect 1917 10364 1981 10368
rect 1917 10308 1921 10364
rect 1921 10308 1977 10364
rect 1977 10308 1981 10364
rect 1917 10304 1981 10308
rect 1997 10364 2061 10368
rect 1997 10308 2001 10364
rect 2001 10308 2057 10364
rect 2057 10308 2061 10364
rect 1997 10304 2061 10308
rect 2077 10364 2141 10368
rect 2077 10308 2081 10364
rect 2081 10308 2137 10364
rect 2137 10308 2141 10364
rect 2077 10304 2141 10308
rect 2157 10364 2221 10368
rect 2157 10308 2161 10364
rect 2161 10308 2217 10364
rect 2217 10308 2221 10364
rect 2157 10304 2221 10308
rect 3848 10364 3912 10368
rect 3848 10308 3852 10364
rect 3852 10308 3908 10364
rect 3908 10308 3912 10364
rect 3848 10304 3912 10308
rect 3928 10364 3992 10368
rect 3928 10308 3932 10364
rect 3932 10308 3988 10364
rect 3988 10308 3992 10364
rect 3928 10304 3992 10308
rect 4008 10364 4072 10368
rect 4008 10308 4012 10364
rect 4012 10308 4068 10364
rect 4068 10308 4072 10364
rect 4008 10304 4072 10308
rect 4088 10364 4152 10368
rect 4088 10308 4092 10364
rect 4092 10308 4148 10364
rect 4148 10308 4152 10364
rect 4088 10304 4152 10308
rect 5778 10364 5842 10368
rect 5778 10308 5782 10364
rect 5782 10308 5838 10364
rect 5838 10308 5842 10364
rect 5778 10304 5842 10308
rect 5858 10364 5922 10368
rect 5858 10308 5862 10364
rect 5862 10308 5918 10364
rect 5918 10308 5922 10364
rect 5858 10304 5922 10308
rect 5938 10364 6002 10368
rect 5938 10308 5942 10364
rect 5942 10308 5998 10364
rect 5998 10308 6002 10364
rect 5938 10304 6002 10308
rect 6018 10364 6082 10368
rect 6018 10308 6022 10364
rect 6022 10308 6078 10364
rect 6078 10308 6082 10364
rect 6018 10304 6082 10308
rect 2882 9820 2946 9824
rect 2882 9764 2886 9820
rect 2886 9764 2942 9820
rect 2942 9764 2946 9820
rect 2882 9760 2946 9764
rect 2962 9820 3026 9824
rect 2962 9764 2966 9820
rect 2966 9764 3022 9820
rect 3022 9764 3026 9820
rect 2962 9760 3026 9764
rect 3042 9820 3106 9824
rect 3042 9764 3046 9820
rect 3046 9764 3102 9820
rect 3102 9764 3106 9820
rect 3042 9760 3106 9764
rect 3122 9820 3186 9824
rect 3122 9764 3126 9820
rect 3126 9764 3182 9820
rect 3182 9764 3186 9820
rect 3122 9760 3186 9764
rect 4813 9820 4877 9824
rect 4813 9764 4817 9820
rect 4817 9764 4873 9820
rect 4873 9764 4877 9820
rect 4813 9760 4877 9764
rect 4893 9820 4957 9824
rect 4893 9764 4897 9820
rect 4897 9764 4953 9820
rect 4953 9764 4957 9820
rect 4893 9760 4957 9764
rect 4973 9820 5037 9824
rect 4973 9764 4977 9820
rect 4977 9764 5033 9820
rect 5033 9764 5037 9820
rect 4973 9760 5037 9764
rect 5053 9820 5117 9824
rect 5053 9764 5057 9820
rect 5057 9764 5113 9820
rect 5113 9764 5117 9820
rect 5053 9760 5117 9764
rect 1917 9276 1981 9280
rect 1917 9220 1921 9276
rect 1921 9220 1977 9276
rect 1977 9220 1981 9276
rect 1917 9216 1981 9220
rect 1997 9276 2061 9280
rect 1997 9220 2001 9276
rect 2001 9220 2057 9276
rect 2057 9220 2061 9276
rect 1997 9216 2061 9220
rect 2077 9276 2141 9280
rect 2077 9220 2081 9276
rect 2081 9220 2137 9276
rect 2137 9220 2141 9276
rect 2077 9216 2141 9220
rect 2157 9276 2221 9280
rect 2157 9220 2161 9276
rect 2161 9220 2217 9276
rect 2217 9220 2221 9276
rect 2157 9216 2221 9220
rect 3848 9276 3912 9280
rect 3848 9220 3852 9276
rect 3852 9220 3908 9276
rect 3908 9220 3912 9276
rect 3848 9216 3912 9220
rect 3928 9276 3992 9280
rect 3928 9220 3932 9276
rect 3932 9220 3988 9276
rect 3988 9220 3992 9276
rect 3928 9216 3992 9220
rect 4008 9276 4072 9280
rect 4008 9220 4012 9276
rect 4012 9220 4068 9276
rect 4068 9220 4072 9276
rect 4008 9216 4072 9220
rect 4088 9276 4152 9280
rect 4088 9220 4092 9276
rect 4092 9220 4148 9276
rect 4148 9220 4152 9276
rect 4088 9216 4152 9220
rect 5778 9276 5842 9280
rect 5778 9220 5782 9276
rect 5782 9220 5838 9276
rect 5838 9220 5842 9276
rect 5778 9216 5842 9220
rect 5858 9276 5922 9280
rect 5858 9220 5862 9276
rect 5862 9220 5918 9276
rect 5918 9220 5922 9276
rect 5858 9216 5922 9220
rect 5938 9276 6002 9280
rect 5938 9220 5942 9276
rect 5942 9220 5998 9276
rect 5998 9220 6002 9276
rect 5938 9216 6002 9220
rect 6018 9276 6082 9280
rect 6018 9220 6022 9276
rect 6022 9220 6078 9276
rect 6078 9220 6082 9276
rect 6018 9216 6082 9220
rect 2882 8732 2946 8736
rect 2882 8676 2886 8732
rect 2886 8676 2942 8732
rect 2942 8676 2946 8732
rect 2882 8672 2946 8676
rect 2962 8732 3026 8736
rect 2962 8676 2966 8732
rect 2966 8676 3022 8732
rect 3022 8676 3026 8732
rect 2962 8672 3026 8676
rect 3042 8732 3106 8736
rect 3042 8676 3046 8732
rect 3046 8676 3102 8732
rect 3102 8676 3106 8732
rect 3042 8672 3106 8676
rect 3122 8732 3186 8736
rect 3122 8676 3126 8732
rect 3126 8676 3182 8732
rect 3182 8676 3186 8732
rect 3122 8672 3186 8676
rect 4813 8732 4877 8736
rect 4813 8676 4817 8732
rect 4817 8676 4873 8732
rect 4873 8676 4877 8732
rect 4813 8672 4877 8676
rect 4893 8732 4957 8736
rect 4893 8676 4897 8732
rect 4897 8676 4953 8732
rect 4953 8676 4957 8732
rect 4893 8672 4957 8676
rect 4973 8732 5037 8736
rect 4973 8676 4977 8732
rect 4977 8676 5033 8732
rect 5033 8676 5037 8732
rect 4973 8672 5037 8676
rect 5053 8732 5117 8736
rect 5053 8676 5057 8732
rect 5057 8676 5113 8732
rect 5113 8676 5117 8732
rect 5053 8672 5117 8676
rect 1917 8188 1981 8192
rect 1917 8132 1921 8188
rect 1921 8132 1977 8188
rect 1977 8132 1981 8188
rect 1917 8128 1981 8132
rect 1997 8188 2061 8192
rect 1997 8132 2001 8188
rect 2001 8132 2057 8188
rect 2057 8132 2061 8188
rect 1997 8128 2061 8132
rect 2077 8188 2141 8192
rect 2077 8132 2081 8188
rect 2081 8132 2137 8188
rect 2137 8132 2141 8188
rect 2077 8128 2141 8132
rect 2157 8188 2221 8192
rect 2157 8132 2161 8188
rect 2161 8132 2217 8188
rect 2217 8132 2221 8188
rect 2157 8128 2221 8132
rect 3848 8188 3912 8192
rect 3848 8132 3852 8188
rect 3852 8132 3908 8188
rect 3908 8132 3912 8188
rect 3848 8128 3912 8132
rect 3928 8188 3992 8192
rect 3928 8132 3932 8188
rect 3932 8132 3988 8188
rect 3988 8132 3992 8188
rect 3928 8128 3992 8132
rect 4008 8188 4072 8192
rect 4008 8132 4012 8188
rect 4012 8132 4068 8188
rect 4068 8132 4072 8188
rect 4008 8128 4072 8132
rect 4088 8188 4152 8192
rect 4088 8132 4092 8188
rect 4092 8132 4148 8188
rect 4148 8132 4152 8188
rect 4088 8128 4152 8132
rect 5778 8188 5842 8192
rect 5778 8132 5782 8188
rect 5782 8132 5838 8188
rect 5838 8132 5842 8188
rect 5778 8128 5842 8132
rect 5858 8188 5922 8192
rect 5858 8132 5862 8188
rect 5862 8132 5918 8188
rect 5918 8132 5922 8188
rect 5858 8128 5922 8132
rect 5938 8188 6002 8192
rect 5938 8132 5942 8188
rect 5942 8132 5998 8188
rect 5998 8132 6002 8188
rect 5938 8128 6002 8132
rect 6018 8188 6082 8192
rect 6018 8132 6022 8188
rect 6022 8132 6078 8188
rect 6078 8132 6082 8188
rect 6018 8128 6082 8132
rect 2882 7644 2946 7648
rect 2882 7588 2886 7644
rect 2886 7588 2942 7644
rect 2942 7588 2946 7644
rect 2882 7584 2946 7588
rect 2962 7644 3026 7648
rect 2962 7588 2966 7644
rect 2966 7588 3022 7644
rect 3022 7588 3026 7644
rect 2962 7584 3026 7588
rect 3042 7644 3106 7648
rect 3042 7588 3046 7644
rect 3046 7588 3102 7644
rect 3102 7588 3106 7644
rect 3042 7584 3106 7588
rect 3122 7644 3186 7648
rect 3122 7588 3126 7644
rect 3126 7588 3182 7644
rect 3182 7588 3186 7644
rect 3122 7584 3186 7588
rect 4813 7644 4877 7648
rect 4813 7588 4817 7644
rect 4817 7588 4873 7644
rect 4873 7588 4877 7644
rect 4813 7584 4877 7588
rect 4893 7644 4957 7648
rect 4893 7588 4897 7644
rect 4897 7588 4953 7644
rect 4953 7588 4957 7644
rect 4893 7584 4957 7588
rect 4973 7644 5037 7648
rect 4973 7588 4977 7644
rect 4977 7588 5033 7644
rect 5033 7588 5037 7644
rect 4973 7584 5037 7588
rect 5053 7644 5117 7648
rect 5053 7588 5057 7644
rect 5057 7588 5113 7644
rect 5113 7588 5117 7644
rect 5053 7584 5117 7588
rect 1917 7100 1981 7104
rect 1917 7044 1921 7100
rect 1921 7044 1977 7100
rect 1977 7044 1981 7100
rect 1917 7040 1981 7044
rect 1997 7100 2061 7104
rect 1997 7044 2001 7100
rect 2001 7044 2057 7100
rect 2057 7044 2061 7100
rect 1997 7040 2061 7044
rect 2077 7100 2141 7104
rect 2077 7044 2081 7100
rect 2081 7044 2137 7100
rect 2137 7044 2141 7100
rect 2077 7040 2141 7044
rect 2157 7100 2221 7104
rect 2157 7044 2161 7100
rect 2161 7044 2217 7100
rect 2217 7044 2221 7100
rect 2157 7040 2221 7044
rect 3848 7100 3912 7104
rect 3848 7044 3852 7100
rect 3852 7044 3908 7100
rect 3908 7044 3912 7100
rect 3848 7040 3912 7044
rect 3928 7100 3992 7104
rect 3928 7044 3932 7100
rect 3932 7044 3988 7100
rect 3988 7044 3992 7100
rect 3928 7040 3992 7044
rect 4008 7100 4072 7104
rect 4008 7044 4012 7100
rect 4012 7044 4068 7100
rect 4068 7044 4072 7100
rect 4008 7040 4072 7044
rect 4088 7100 4152 7104
rect 4088 7044 4092 7100
rect 4092 7044 4148 7100
rect 4148 7044 4152 7100
rect 4088 7040 4152 7044
rect 5778 7100 5842 7104
rect 5778 7044 5782 7100
rect 5782 7044 5838 7100
rect 5838 7044 5842 7100
rect 5778 7040 5842 7044
rect 5858 7100 5922 7104
rect 5858 7044 5862 7100
rect 5862 7044 5918 7100
rect 5918 7044 5922 7100
rect 5858 7040 5922 7044
rect 5938 7100 6002 7104
rect 5938 7044 5942 7100
rect 5942 7044 5998 7100
rect 5998 7044 6002 7100
rect 5938 7040 6002 7044
rect 6018 7100 6082 7104
rect 6018 7044 6022 7100
rect 6022 7044 6078 7100
rect 6078 7044 6082 7100
rect 6018 7040 6082 7044
rect 2882 6556 2946 6560
rect 2882 6500 2886 6556
rect 2886 6500 2942 6556
rect 2942 6500 2946 6556
rect 2882 6496 2946 6500
rect 2962 6556 3026 6560
rect 2962 6500 2966 6556
rect 2966 6500 3022 6556
rect 3022 6500 3026 6556
rect 2962 6496 3026 6500
rect 3042 6556 3106 6560
rect 3042 6500 3046 6556
rect 3046 6500 3102 6556
rect 3102 6500 3106 6556
rect 3042 6496 3106 6500
rect 3122 6556 3186 6560
rect 3122 6500 3126 6556
rect 3126 6500 3182 6556
rect 3182 6500 3186 6556
rect 3122 6496 3186 6500
rect 4813 6556 4877 6560
rect 4813 6500 4817 6556
rect 4817 6500 4873 6556
rect 4873 6500 4877 6556
rect 4813 6496 4877 6500
rect 4893 6556 4957 6560
rect 4893 6500 4897 6556
rect 4897 6500 4953 6556
rect 4953 6500 4957 6556
rect 4893 6496 4957 6500
rect 4973 6556 5037 6560
rect 4973 6500 4977 6556
rect 4977 6500 5033 6556
rect 5033 6500 5037 6556
rect 4973 6496 5037 6500
rect 5053 6556 5117 6560
rect 5053 6500 5057 6556
rect 5057 6500 5113 6556
rect 5113 6500 5117 6556
rect 5053 6496 5117 6500
rect 1917 6012 1981 6016
rect 1917 5956 1921 6012
rect 1921 5956 1977 6012
rect 1977 5956 1981 6012
rect 1917 5952 1981 5956
rect 1997 6012 2061 6016
rect 1997 5956 2001 6012
rect 2001 5956 2057 6012
rect 2057 5956 2061 6012
rect 1997 5952 2061 5956
rect 2077 6012 2141 6016
rect 2077 5956 2081 6012
rect 2081 5956 2137 6012
rect 2137 5956 2141 6012
rect 2077 5952 2141 5956
rect 2157 6012 2221 6016
rect 2157 5956 2161 6012
rect 2161 5956 2217 6012
rect 2217 5956 2221 6012
rect 2157 5952 2221 5956
rect 3848 6012 3912 6016
rect 3848 5956 3852 6012
rect 3852 5956 3908 6012
rect 3908 5956 3912 6012
rect 3848 5952 3912 5956
rect 3928 6012 3992 6016
rect 3928 5956 3932 6012
rect 3932 5956 3988 6012
rect 3988 5956 3992 6012
rect 3928 5952 3992 5956
rect 4008 6012 4072 6016
rect 4008 5956 4012 6012
rect 4012 5956 4068 6012
rect 4068 5956 4072 6012
rect 4008 5952 4072 5956
rect 4088 6012 4152 6016
rect 4088 5956 4092 6012
rect 4092 5956 4148 6012
rect 4148 5956 4152 6012
rect 4088 5952 4152 5956
rect 5778 6012 5842 6016
rect 5778 5956 5782 6012
rect 5782 5956 5838 6012
rect 5838 5956 5842 6012
rect 5778 5952 5842 5956
rect 5858 6012 5922 6016
rect 5858 5956 5862 6012
rect 5862 5956 5918 6012
rect 5918 5956 5922 6012
rect 5858 5952 5922 5956
rect 5938 6012 6002 6016
rect 5938 5956 5942 6012
rect 5942 5956 5998 6012
rect 5998 5956 6002 6012
rect 5938 5952 6002 5956
rect 6018 6012 6082 6016
rect 6018 5956 6022 6012
rect 6022 5956 6078 6012
rect 6078 5956 6082 6012
rect 6018 5952 6082 5956
rect 2882 5468 2946 5472
rect 2882 5412 2886 5468
rect 2886 5412 2942 5468
rect 2942 5412 2946 5468
rect 2882 5408 2946 5412
rect 2962 5468 3026 5472
rect 2962 5412 2966 5468
rect 2966 5412 3022 5468
rect 3022 5412 3026 5468
rect 2962 5408 3026 5412
rect 3042 5468 3106 5472
rect 3042 5412 3046 5468
rect 3046 5412 3102 5468
rect 3102 5412 3106 5468
rect 3042 5408 3106 5412
rect 3122 5468 3186 5472
rect 3122 5412 3126 5468
rect 3126 5412 3182 5468
rect 3182 5412 3186 5468
rect 3122 5408 3186 5412
rect 4813 5468 4877 5472
rect 4813 5412 4817 5468
rect 4817 5412 4873 5468
rect 4873 5412 4877 5468
rect 4813 5408 4877 5412
rect 4893 5468 4957 5472
rect 4893 5412 4897 5468
rect 4897 5412 4953 5468
rect 4953 5412 4957 5468
rect 4893 5408 4957 5412
rect 4973 5468 5037 5472
rect 4973 5412 4977 5468
rect 4977 5412 5033 5468
rect 5033 5412 5037 5468
rect 4973 5408 5037 5412
rect 5053 5468 5117 5472
rect 5053 5412 5057 5468
rect 5057 5412 5113 5468
rect 5113 5412 5117 5468
rect 5053 5408 5117 5412
rect 1917 4924 1981 4928
rect 1917 4868 1921 4924
rect 1921 4868 1977 4924
rect 1977 4868 1981 4924
rect 1917 4864 1981 4868
rect 1997 4924 2061 4928
rect 1997 4868 2001 4924
rect 2001 4868 2057 4924
rect 2057 4868 2061 4924
rect 1997 4864 2061 4868
rect 2077 4924 2141 4928
rect 2077 4868 2081 4924
rect 2081 4868 2137 4924
rect 2137 4868 2141 4924
rect 2077 4864 2141 4868
rect 2157 4924 2221 4928
rect 2157 4868 2161 4924
rect 2161 4868 2217 4924
rect 2217 4868 2221 4924
rect 2157 4864 2221 4868
rect 3848 4924 3912 4928
rect 3848 4868 3852 4924
rect 3852 4868 3908 4924
rect 3908 4868 3912 4924
rect 3848 4864 3912 4868
rect 3928 4924 3992 4928
rect 3928 4868 3932 4924
rect 3932 4868 3988 4924
rect 3988 4868 3992 4924
rect 3928 4864 3992 4868
rect 4008 4924 4072 4928
rect 4008 4868 4012 4924
rect 4012 4868 4068 4924
rect 4068 4868 4072 4924
rect 4008 4864 4072 4868
rect 4088 4924 4152 4928
rect 4088 4868 4092 4924
rect 4092 4868 4148 4924
rect 4148 4868 4152 4924
rect 4088 4864 4152 4868
rect 5778 4924 5842 4928
rect 5778 4868 5782 4924
rect 5782 4868 5838 4924
rect 5838 4868 5842 4924
rect 5778 4864 5842 4868
rect 5858 4924 5922 4928
rect 5858 4868 5862 4924
rect 5862 4868 5918 4924
rect 5918 4868 5922 4924
rect 5858 4864 5922 4868
rect 5938 4924 6002 4928
rect 5938 4868 5942 4924
rect 5942 4868 5998 4924
rect 5998 4868 6002 4924
rect 5938 4864 6002 4868
rect 6018 4924 6082 4928
rect 6018 4868 6022 4924
rect 6022 4868 6078 4924
rect 6078 4868 6082 4924
rect 6018 4864 6082 4868
rect 2882 4380 2946 4384
rect 2882 4324 2886 4380
rect 2886 4324 2942 4380
rect 2942 4324 2946 4380
rect 2882 4320 2946 4324
rect 2962 4380 3026 4384
rect 2962 4324 2966 4380
rect 2966 4324 3022 4380
rect 3022 4324 3026 4380
rect 2962 4320 3026 4324
rect 3042 4380 3106 4384
rect 3042 4324 3046 4380
rect 3046 4324 3102 4380
rect 3102 4324 3106 4380
rect 3042 4320 3106 4324
rect 3122 4380 3186 4384
rect 3122 4324 3126 4380
rect 3126 4324 3182 4380
rect 3182 4324 3186 4380
rect 3122 4320 3186 4324
rect 4813 4380 4877 4384
rect 4813 4324 4817 4380
rect 4817 4324 4873 4380
rect 4873 4324 4877 4380
rect 4813 4320 4877 4324
rect 4893 4380 4957 4384
rect 4893 4324 4897 4380
rect 4897 4324 4953 4380
rect 4953 4324 4957 4380
rect 4893 4320 4957 4324
rect 4973 4380 5037 4384
rect 4973 4324 4977 4380
rect 4977 4324 5033 4380
rect 5033 4324 5037 4380
rect 4973 4320 5037 4324
rect 5053 4380 5117 4384
rect 5053 4324 5057 4380
rect 5057 4324 5113 4380
rect 5113 4324 5117 4380
rect 5053 4320 5117 4324
rect 1917 3836 1981 3840
rect 1917 3780 1921 3836
rect 1921 3780 1977 3836
rect 1977 3780 1981 3836
rect 1917 3776 1981 3780
rect 1997 3836 2061 3840
rect 1997 3780 2001 3836
rect 2001 3780 2057 3836
rect 2057 3780 2061 3836
rect 1997 3776 2061 3780
rect 2077 3836 2141 3840
rect 2077 3780 2081 3836
rect 2081 3780 2137 3836
rect 2137 3780 2141 3836
rect 2077 3776 2141 3780
rect 2157 3836 2221 3840
rect 2157 3780 2161 3836
rect 2161 3780 2217 3836
rect 2217 3780 2221 3836
rect 2157 3776 2221 3780
rect 3848 3836 3912 3840
rect 3848 3780 3852 3836
rect 3852 3780 3908 3836
rect 3908 3780 3912 3836
rect 3848 3776 3912 3780
rect 3928 3836 3992 3840
rect 3928 3780 3932 3836
rect 3932 3780 3988 3836
rect 3988 3780 3992 3836
rect 3928 3776 3992 3780
rect 4008 3836 4072 3840
rect 4008 3780 4012 3836
rect 4012 3780 4068 3836
rect 4068 3780 4072 3836
rect 4008 3776 4072 3780
rect 4088 3836 4152 3840
rect 4088 3780 4092 3836
rect 4092 3780 4148 3836
rect 4148 3780 4152 3836
rect 4088 3776 4152 3780
rect 5778 3836 5842 3840
rect 5778 3780 5782 3836
rect 5782 3780 5838 3836
rect 5838 3780 5842 3836
rect 5778 3776 5842 3780
rect 5858 3836 5922 3840
rect 5858 3780 5862 3836
rect 5862 3780 5918 3836
rect 5918 3780 5922 3836
rect 5858 3776 5922 3780
rect 5938 3836 6002 3840
rect 5938 3780 5942 3836
rect 5942 3780 5998 3836
rect 5998 3780 6002 3836
rect 5938 3776 6002 3780
rect 6018 3836 6082 3840
rect 6018 3780 6022 3836
rect 6022 3780 6078 3836
rect 6078 3780 6082 3836
rect 6018 3776 6082 3780
rect 2882 3292 2946 3296
rect 2882 3236 2886 3292
rect 2886 3236 2942 3292
rect 2942 3236 2946 3292
rect 2882 3232 2946 3236
rect 2962 3292 3026 3296
rect 2962 3236 2966 3292
rect 2966 3236 3022 3292
rect 3022 3236 3026 3292
rect 2962 3232 3026 3236
rect 3042 3292 3106 3296
rect 3042 3236 3046 3292
rect 3046 3236 3102 3292
rect 3102 3236 3106 3292
rect 3042 3232 3106 3236
rect 3122 3292 3186 3296
rect 3122 3236 3126 3292
rect 3126 3236 3182 3292
rect 3182 3236 3186 3292
rect 3122 3232 3186 3236
rect 4813 3292 4877 3296
rect 4813 3236 4817 3292
rect 4817 3236 4873 3292
rect 4873 3236 4877 3292
rect 4813 3232 4877 3236
rect 4893 3292 4957 3296
rect 4893 3236 4897 3292
rect 4897 3236 4953 3292
rect 4953 3236 4957 3292
rect 4893 3232 4957 3236
rect 4973 3292 5037 3296
rect 4973 3236 4977 3292
rect 4977 3236 5033 3292
rect 5033 3236 5037 3292
rect 4973 3232 5037 3236
rect 5053 3292 5117 3296
rect 5053 3236 5057 3292
rect 5057 3236 5113 3292
rect 5113 3236 5117 3292
rect 5053 3232 5117 3236
rect 1917 2748 1981 2752
rect 1917 2692 1921 2748
rect 1921 2692 1977 2748
rect 1977 2692 1981 2748
rect 1917 2688 1981 2692
rect 1997 2748 2061 2752
rect 1997 2692 2001 2748
rect 2001 2692 2057 2748
rect 2057 2692 2061 2748
rect 1997 2688 2061 2692
rect 2077 2748 2141 2752
rect 2077 2692 2081 2748
rect 2081 2692 2137 2748
rect 2137 2692 2141 2748
rect 2077 2688 2141 2692
rect 2157 2748 2221 2752
rect 2157 2692 2161 2748
rect 2161 2692 2217 2748
rect 2217 2692 2221 2748
rect 2157 2688 2221 2692
rect 3848 2748 3912 2752
rect 3848 2692 3852 2748
rect 3852 2692 3908 2748
rect 3908 2692 3912 2748
rect 3848 2688 3912 2692
rect 3928 2748 3992 2752
rect 3928 2692 3932 2748
rect 3932 2692 3988 2748
rect 3988 2692 3992 2748
rect 3928 2688 3992 2692
rect 4008 2748 4072 2752
rect 4008 2692 4012 2748
rect 4012 2692 4068 2748
rect 4068 2692 4072 2748
rect 4008 2688 4072 2692
rect 4088 2748 4152 2752
rect 4088 2692 4092 2748
rect 4092 2692 4148 2748
rect 4148 2692 4152 2748
rect 4088 2688 4152 2692
rect 5778 2748 5842 2752
rect 5778 2692 5782 2748
rect 5782 2692 5838 2748
rect 5838 2692 5842 2748
rect 5778 2688 5842 2692
rect 5858 2748 5922 2752
rect 5858 2692 5862 2748
rect 5862 2692 5918 2748
rect 5918 2692 5922 2748
rect 5858 2688 5922 2692
rect 5938 2748 6002 2752
rect 5938 2692 5942 2748
rect 5942 2692 5998 2748
rect 5998 2692 6002 2748
rect 5938 2688 6002 2692
rect 6018 2748 6082 2752
rect 6018 2692 6022 2748
rect 6022 2692 6078 2748
rect 6078 2692 6082 2748
rect 6018 2688 6082 2692
rect 2882 2204 2946 2208
rect 2882 2148 2886 2204
rect 2886 2148 2942 2204
rect 2942 2148 2946 2204
rect 2882 2144 2946 2148
rect 2962 2204 3026 2208
rect 2962 2148 2966 2204
rect 2966 2148 3022 2204
rect 3022 2148 3026 2204
rect 2962 2144 3026 2148
rect 3042 2204 3106 2208
rect 3042 2148 3046 2204
rect 3046 2148 3102 2204
rect 3102 2148 3106 2204
rect 3042 2144 3106 2148
rect 3122 2204 3186 2208
rect 3122 2148 3126 2204
rect 3126 2148 3182 2204
rect 3182 2148 3186 2204
rect 3122 2144 3186 2148
rect 4813 2204 4877 2208
rect 4813 2148 4817 2204
rect 4817 2148 4873 2204
rect 4873 2148 4877 2204
rect 4813 2144 4877 2148
rect 4893 2204 4957 2208
rect 4893 2148 4897 2204
rect 4897 2148 4953 2204
rect 4953 2148 4957 2204
rect 4893 2144 4957 2148
rect 4973 2204 5037 2208
rect 4973 2148 4977 2204
rect 4977 2148 5033 2204
rect 5033 2148 5037 2204
rect 4973 2144 5037 2148
rect 5053 2204 5117 2208
rect 5053 2148 5057 2204
rect 5057 2148 5113 2204
rect 5113 2148 5117 2204
rect 5053 2144 5117 2148
<< metal4 >>
rect 1909 57152 2229 57712
rect 1909 57088 1917 57152
rect 1981 57088 1997 57152
rect 2061 57088 2077 57152
rect 2141 57088 2157 57152
rect 2221 57088 2229 57152
rect 1909 56064 2229 57088
rect 1909 56000 1917 56064
rect 1981 56000 1997 56064
rect 2061 56000 2077 56064
rect 2141 56000 2157 56064
rect 2221 56000 2229 56064
rect 1909 54976 2229 56000
rect 1909 54912 1917 54976
rect 1981 54912 1997 54976
rect 2061 54912 2077 54976
rect 2141 54912 2157 54976
rect 2221 54912 2229 54976
rect 1909 53888 2229 54912
rect 1909 53824 1917 53888
rect 1981 53824 1997 53888
rect 2061 53824 2077 53888
rect 2141 53824 2157 53888
rect 2221 53824 2229 53888
rect 1909 52800 2229 53824
rect 1909 52736 1917 52800
rect 1981 52736 1997 52800
rect 2061 52736 2077 52800
rect 2141 52736 2157 52800
rect 2221 52736 2229 52800
rect 1909 51712 2229 52736
rect 1909 51648 1917 51712
rect 1981 51648 1997 51712
rect 2061 51648 2077 51712
rect 2141 51648 2157 51712
rect 2221 51648 2229 51712
rect 1909 50624 2229 51648
rect 1909 50560 1917 50624
rect 1981 50560 1997 50624
rect 2061 50560 2077 50624
rect 2141 50560 2157 50624
rect 2221 50560 2229 50624
rect 1909 49536 2229 50560
rect 1909 49472 1917 49536
rect 1981 49472 1997 49536
rect 2061 49472 2077 49536
rect 2141 49472 2157 49536
rect 2221 49472 2229 49536
rect 1909 48448 2229 49472
rect 1909 48384 1917 48448
rect 1981 48384 1997 48448
rect 2061 48384 2077 48448
rect 2141 48384 2157 48448
rect 2221 48384 2229 48448
rect 1909 47360 2229 48384
rect 2874 57696 3194 57712
rect 2874 57632 2882 57696
rect 2946 57632 2962 57696
rect 3026 57632 3042 57696
rect 3106 57632 3122 57696
rect 3186 57632 3194 57696
rect 2874 56608 3194 57632
rect 2874 56544 2882 56608
rect 2946 56544 2962 56608
rect 3026 56544 3042 56608
rect 3106 56544 3122 56608
rect 3186 56544 3194 56608
rect 2874 55520 3194 56544
rect 2874 55456 2882 55520
rect 2946 55456 2962 55520
rect 3026 55456 3042 55520
rect 3106 55456 3122 55520
rect 3186 55456 3194 55520
rect 2874 54432 3194 55456
rect 2874 54368 2882 54432
rect 2946 54368 2962 54432
rect 3026 54368 3042 54432
rect 3106 54368 3122 54432
rect 3186 54368 3194 54432
rect 2874 53344 3194 54368
rect 2874 53280 2882 53344
rect 2946 53280 2962 53344
rect 3026 53280 3042 53344
rect 3106 53280 3122 53344
rect 3186 53280 3194 53344
rect 2874 52256 3194 53280
rect 2874 52192 2882 52256
rect 2946 52192 2962 52256
rect 3026 52192 3042 52256
rect 3106 52192 3122 52256
rect 3186 52192 3194 52256
rect 2874 51168 3194 52192
rect 2874 51104 2882 51168
rect 2946 51104 2962 51168
rect 3026 51104 3042 51168
rect 3106 51104 3122 51168
rect 3186 51104 3194 51168
rect 2874 50080 3194 51104
rect 2874 50016 2882 50080
rect 2946 50016 2962 50080
rect 3026 50016 3042 50080
rect 3106 50016 3122 50080
rect 3186 50016 3194 50080
rect 2874 48992 3194 50016
rect 2874 48928 2882 48992
rect 2946 48928 2962 48992
rect 3026 48928 3042 48992
rect 3106 48928 3122 48992
rect 3186 48928 3194 48992
rect 2635 48108 2701 48109
rect 2635 48044 2636 48108
rect 2700 48044 2701 48108
rect 2635 48043 2701 48044
rect 1909 47296 1917 47360
rect 1981 47296 1997 47360
rect 2061 47296 2077 47360
rect 2141 47296 2157 47360
rect 2221 47296 2229 47360
rect 1909 46272 2229 47296
rect 1909 46208 1917 46272
rect 1981 46208 1997 46272
rect 2061 46208 2077 46272
rect 2141 46208 2157 46272
rect 2221 46208 2229 46272
rect 1909 45184 2229 46208
rect 1909 45120 1917 45184
rect 1981 45120 1997 45184
rect 2061 45120 2077 45184
rect 2141 45120 2157 45184
rect 2221 45120 2229 45184
rect 1909 44096 2229 45120
rect 1909 44032 1917 44096
rect 1981 44032 1997 44096
rect 2061 44032 2077 44096
rect 2141 44032 2157 44096
rect 2221 44032 2229 44096
rect 1909 43008 2229 44032
rect 1909 42944 1917 43008
rect 1981 42944 1997 43008
rect 2061 42944 2077 43008
rect 2141 42944 2157 43008
rect 2221 42944 2229 43008
rect 1909 41920 2229 42944
rect 1909 41856 1917 41920
rect 1981 41856 1997 41920
rect 2061 41856 2077 41920
rect 2141 41856 2157 41920
rect 2221 41856 2229 41920
rect 1715 41580 1781 41581
rect 1715 41516 1716 41580
rect 1780 41516 1781 41580
rect 1715 41515 1781 41516
rect 1718 37909 1778 41515
rect 1909 40832 2229 41856
rect 1909 40768 1917 40832
rect 1981 40768 1997 40832
rect 2061 40768 2077 40832
rect 2141 40768 2157 40832
rect 2221 40768 2229 40832
rect 1909 39744 2229 40768
rect 1909 39680 1917 39744
rect 1981 39680 1997 39744
rect 2061 39680 2077 39744
rect 2141 39680 2157 39744
rect 2221 39680 2229 39744
rect 1909 38656 2229 39680
rect 2638 38997 2698 48043
rect 2874 47904 3194 48928
rect 2874 47840 2882 47904
rect 2946 47840 2962 47904
rect 3026 47840 3042 47904
rect 3106 47840 3122 47904
rect 3186 47840 3194 47904
rect 2874 46816 3194 47840
rect 2874 46752 2882 46816
rect 2946 46752 2962 46816
rect 3026 46752 3042 46816
rect 3106 46752 3122 46816
rect 3186 46752 3194 46816
rect 2874 45728 3194 46752
rect 2874 45664 2882 45728
rect 2946 45664 2962 45728
rect 3026 45664 3042 45728
rect 3106 45664 3122 45728
rect 3186 45664 3194 45728
rect 2874 44640 3194 45664
rect 2874 44576 2882 44640
rect 2946 44576 2962 44640
rect 3026 44576 3042 44640
rect 3106 44576 3122 44640
rect 3186 44576 3194 44640
rect 2874 43552 3194 44576
rect 3839 57152 4160 57712
rect 3839 57088 3848 57152
rect 3912 57088 3928 57152
rect 3992 57088 4008 57152
rect 4072 57088 4088 57152
rect 4152 57088 4160 57152
rect 3839 56064 4160 57088
rect 3839 56000 3848 56064
rect 3912 56000 3928 56064
rect 3992 56000 4008 56064
rect 4072 56000 4088 56064
rect 4152 56000 4160 56064
rect 3839 54976 4160 56000
rect 4805 57696 5125 57712
rect 4805 57632 4813 57696
rect 4877 57632 4893 57696
rect 4957 57632 4973 57696
rect 5037 57632 5053 57696
rect 5117 57632 5125 57696
rect 4805 56608 5125 57632
rect 4805 56544 4813 56608
rect 4877 56544 4893 56608
rect 4957 56544 4973 56608
rect 5037 56544 5053 56608
rect 5117 56544 5125 56608
rect 4805 55520 5125 56544
rect 4805 55456 4813 55520
rect 4877 55456 4893 55520
rect 4957 55456 4973 55520
rect 5037 55456 5053 55520
rect 5117 55456 5125 55520
rect 4291 55316 4357 55317
rect 4291 55252 4292 55316
rect 4356 55252 4357 55316
rect 4291 55251 4357 55252
rect 3839 54912 3848 54976
rect 3912 54912 3928 54976
rect 3992 54912 4008 54976
rect 4072 54912 4088 54976
rect 4152 54912 4160 54976
rect 3839 53888 4160 54912
rect 3839 53824 3848 53888
rect 3912 53824 3928 53888
rect 3992 53824 4008 53888
rect 4072 53824 4088 53888
rect 4152 53824 4160 53888
rect 3839 52800 4160 53824
rect 3839 52736 3848 52800
rect 3912 52736 3928 52800
rect 3992 52736 4008 52800
rect 4072 52736 4088 52800
rect 4152 52736 4160 52800
rect 3839 51712 4160 52736
rect 3839 51648 3848 51712
rect 3912 51648 3928 51712
rect 3992 51648 4008 51712
rect 4072 51648 4088 51712
rect 4152 51648 4160 51712
rect 3839 50624 4160 51648
rect 3839 50560 3848 50624
rect 3912 50560 3928 50624
rect 3992 50560 4008 50624
rect 4072 50560 4088 50624
rect 4152 50560 4160 50624
rect 3839 49536 4160 50560
rect 3839 49472 3848 49536
rect 3912 49472 3928 49536
rect 3992 49472 4008 49536
rect 4072 49472 4088 49536
rect 4152 49472 4160 49536
rect 3839 48448 4160 49472
rect 3839 48384 3848 48448
rect 3912 48384 3928 48448
rect 3992 48384 4008 48448
rect 4072 48384 4088 48448
rect 4152 48384 4160 48448
rect 3839 47360 4160 48384
rect 3839 47296 3848 47360
rect 3912 47296 3928 47360
rect 3992 47296 4008 47360
rect 4072 47296 4088 47360
rect 4152 47296 4160 47360
rect 3839 46272 4160 47296
rect 3839 46208 3848 46272
rect 3912 46208 3928 46272
rect 3992 46208 4008 46272
rect 4072 46208 4088 46272
rect 4152 46208 4160 46272
rect 3839 45184 4160 46208
rect 3839 45120 3848 45184
rect 3912 45120 3928 45184
rect 3992 45120 4008 45184
rect 4072 45120 4088 45184
rect 4152 45120 4160 45184
rect 3839 44096 4160 45120
rect 3839 44032 3848 44096
rect 3912 44032 3928 44096
rect 3992 44032 4008 44096
rect 4072 44032 4088 44096
rect 4152 44032 4160 44096
rect 3371 43756 3437 43757
rect 3371 43692 3372 43756
rect 3436 43692 3437 43756
rect 3371 43691 3437 43692
rect 2874 43488 2882 43552
rect 2946 43488 2962 43552
rect 3026 43488 3042 43552
rect 3106 43488 3122 43552
rect 3186 43488 3194 43552
rect 2874 42464 3194 43488
rect 2874 42400 2882 42464
rect 2946 42400 2962 42464
rect 3026 42400 3042 42464
rect 3106 42400 3122 42464
rect 3186 42400 3194 42464
rect 2874 41376 3194 42400
rect 2874 41312 2882 41376
rect 2946 41312 2962 41376
rect 3026 41312 3042 41376
rect 3106 41312 3122 41376
rect 3186 41312 3194 41376
rect 2874 40288 3194 41312
rect 3374 41173 3434 43691
rect 3839 43008 4160 44032
rect 3839 42944 3848 43008
rect 3912 42944 3928 43008
rect 3992 42944 4008 43008
rect 4072 42944 4088 43008
rect 4152 42944 4160 43008
rect 3555 42124 3621 42125
rect 3555 42060 3556 42124
rect 3620 42060 3621 42124
rect 3555 42059 3621 42060
rect 3371 41172 3437 41173
rect 3371 41108 3372 41172
rect 3436 41108 3437 41172
rect 3371 41107 3437 41108
rect 2874 40224 2882 40288
rect 2946 40224 2962 40288
rect 3026 40224 3042 40288
rect 3106 40224 3122 40288
rect 3186 40224 3194 40288
rect 2874 39200 3194 40224
rect 2874 39136 2882 39200
rect 2946 39136 2962 39200
rect 3026 39136 3042 39200
rect 3106 39136 3122 39200
rect 3186 39136 3194 39200
rect 2635 38996 2701 38997
rect 2635 38932 2636 38996
rect 2700 38932 2701 38996
rect 2635 38931 2701 38932
rect 2635 38724 2701 38725
rect 2635 38660 2636 38724
rect 2700 38660 2701 38724
rect 2635 38659 2701 38660
rect 1909 38592 1917 38656
rect 1981 38592 1997 38656
rect 2061 38592 2077 38656
rect 2141 38592 2157 38656
rect 2221 38592 2229 38656
rect 1715 37908 1781 37909
rect 1715 37844 1716 37908
rect 1780 37844 1781 37908
rect 1715 37843 1781 37844
rect 1909 37568 2229 38592
rect 2451 38588 2517 38589
rect 2451 38524 2452 38588
rect 2516 38524 2517 38588
rect 2451 38523 2517 38524
rect 1909 37504 1917 37568
rect 1981 37504 1997 37568
rect 2061 37504 2077 37568
rect 2141 37504 2157 37568
rect 2221 37504 2229 37568
rect 1909 36480 2229 37504
rect 1909 36416 1917 36480
rect 1981 36416 1997 36480
rect 2061 36416 2077 36480
rect 2141 36416 2157 36480
rect 2221 36416 2229 36480
rect 1909 35392 2229 36416
rect 1909 35328 1917 35392
rect 1981 35328 1997 35392
rect 2061 35328 2077 35392
rect 2141 35328 2157 35392
rect 2221 35328 2229 35392
rect 1909 34304 2229 35328
rect 1909 34240 1917 34304
rect 1981 34240 1997 34304
rect 2061 34240 2077 34304
rect 2141 34240 2157 34304
rect 2221 34240 2229 34304
rect 1909 33216 2229 34240
rect 1909 33152 1917 33216
rect 1981 33152 1997 33216
rect 2061 33152 2077 33216
rect 2141 33152 2157 33216
rect 2221 33152 2229 33216
rect 1909 32128 2229 33152
rect 1909 32064 1917 32128
rect 1981 32064 1997 32128
rect 2061 32064 2077 32128
rect 2141 32064 2157 32128
rect 2221 32064 2229 32128
rect 1909 31040 2229 32064
rect 2454 31245 2514 38523
rect 2638 36957 2698 38659
rect 2874 38112 3194 39136
rect 3371 38316 3437 38317
rect 3371 38252 3372 38316
rect 3436 38252 3437 38316
rect 3371 38251 3437 38252
rect 2874 38048 2882 38112
rect 2946 38048 2962 38112
rect 3026 38048 3042 38112
rect 3106 38048 3122 38112
rect 3186 38048 3194 38112
rect 2874 37024 3194 38048
rect 2874 36960 2882 37024
rect 2946 36960 2962 37024
rect 3026 36960 3042 37024
rect 3106 36960 3122 37024
rect 3186 36960 3194 37024
rect 2635 36956 2701 36957
rect 2635 36892 2636 36956
rect 2700 36892 2701 36956
rect 2635 36891 2701 36892
rect 2874 35936 3194 36960
rect 2874 35872 2882 35936
rect 2946 35872 2962 35936
rect 3026 35872 3042 35936
rect 3106 35872 3122 35936
rect 3186 35872 3194 35936
rect 2874 34848 3194 35872
rect 2874 34784 2882 34848
rect 2946 34784 2962 34848
rect 3026 34784 3042 34848
rect 3106 34784 3122 34848
rect 3186 34784 3194 34848
rect 2874 33760 3194 34784
rect 2874 33696 2882 33760
rect 2946 33696 2962 33760
rect 3026 33696 3042 33760
rect 3106 33696 3122 33760
rect 3186 33696 3194 33760
rect 2874 32672 3194 33696
rect 2874 32608 2882 32672
rect 2946 32608 2962 32672
rect 3026 32608 3042 32672
rect 3106 32608 3122 32672
rect 3186 32608 3194 32672
rect 2874 31584 3194 32608
rect 2874 31520 2882 31584
rect 2946 31520 2962 31584
rect 3026 31520 3042 31584
rect 3106 31520 3122 31584
rect 3186 31520 3194 31584
rect 2451 31244 2517 31245
rect 2451 31180 2452 31244
rect 2516 31180 2517 31244
rect 2451 31179 2517 31180
rect 1909 30976 1917 31040
rect 1981 30976 1997 31040
rect 2061 30976 2077 31040
rect 2141 30976 2157 31040
rect 2221 30976 2229 31040
rect 1909 29952 2229 30976
rect 1909 29888 1917 29952
rect 1981 29888 1997 29952
rect 2061 29888 2077 29952
rect 2141 29888 2157 29952
rect 2221 29888 2229 29952
rect 1909 28864 2229 29888
rect 1909 28800 1917 28864
rect 1981 28800 1997 28864
rect 2061 28800 2077 28864
rect 2141 28800 2157 28864
rect 2221 28800 2229 28864
rect 1909 27776 2229 28800
rect 1909 27712 1917 27776
rect 1981 27712 1997 27776
rect 2061 27712 2077 27776
rect 2141 27712 2157 27776
rect 2221 27712 2229 27776
rect 1909 26688 2229 27712
rect 1909 26624 1917 26688
rect 1981 26624 1997 26688
rect 2061 26624 2077 26688
rect 2141 26624 2157 26688
rect 2221 26624 2229 26688
rect 1909 25600 2229 26624
rect 1909 25536 1917 25600
rect 1981 25536 1997 25600
rect 2061 25536 2077 25600
rect 2141 25536 2157 25600
rect 2221 25536 2229 25600
rect 1909 24512 2229 25536
rect 1909 24448 1917 24512
rect 1981 24448 1997 24512
rect 2061 24448 2077 24512
rect 2141 24448 2157 24512
rect 2221 24448 2229 24512
rect 1909 23424 2229 24448
rect 1909 23360 1917 23424
rect 1981 23360 1997 23424
rect 2061 23360 2077 23424
rect 2141 23360 2157 23424
rect 2221 23360 2229 23424
rect 1909 22336 2229 23360
rect 1909 22272 1917 22336
rect 1981 22272 1997 22336
rect 2061 22272 2077 22336
rect 2141 22272 2157 22336
rect 2221 22272 2229 22336
rect 1909 21248 2229 22272
rect 1909 21184 1917 21248
rect 1981 21184 1997 21248
rect 2061 21184 2077 21248
rect 2141 21184 2157 21248
rect 2221 21184 2229 21248
rect 1909 20160 2229 21184
rect 1909 20096 1917 20160
rect 1981 20096 1997 20160
rect 2061 20096 2077 20160
rect 2141 20096 2157 20160
rect 2221 20096 2229 20160
rect 1909 19072 2229 20096
rect 1909 19008 1917 19072
rect 1981 19008 1997 19072
rect 2061 19008 2077 19072
rect 2141 19008 2157 19072
rect 2221 19008 2229 19072
rect 1909 17984 2229 19008
rect 1909 17920 1917 17984
rect 1981 17920 1997 17984
rect 2061 17920 2077 17984
rect 2141 17920 2157 17984
rect 2221 17920 2229 17984
rect 1909 16896 2229 17920
rect 1909 16832 1917 16896
rect 1981 16832 1997 16896
rect 2061 16832 2077 16896
rect 2141 16832 2157 16896
rect 2221 16832 2229 16896
rect 1909 15808 2229 16832
rect 1909 15744 1917 15808
rect 1981 15744 1997 15808
rect 2061 15744 2077 15808
rect 2141 15744 2157 15808
rect 2221 15744 2229 15808
rect 1909 14720 2229 15744
rect 1909 14656 1917 14720
rect 1981 14656 1997 14720
rect 2061 14656 2077 14720
rect 2141 14656 2157 14720
rect 2221 14656 2229 14720
rect 1909 13632 2229 14656
rect 1909 13568 1917 13632
rect 1981 13568 1997 13632
rect 2061 13568 2077 13632
rect 2141 13568 2157 13632
rect 2221 13568 2229 13632
rect 1909 12544 2229 13568
rect 1909 12480 1917 12544
rect 1981 12480 1997 12544
rect 2061 12480 2077 12544
rect 2141 12480 2157 12544
rect 2221 12480 2229 12544
rect 1909 11456 2229 12480
rect 1909 11392 1917 11456
rect 1981 11392 1997 11456
rect 2061 11392 2077 11456
rect 2141 11392 2157 11456
rect 2221 11392 2229 11456
rect 1909 10368 2229 11392
rect 1909 10304 1917 10368
rect 1981 10304 1997 10368
rect 2061 10304 2077 10368
rect 2141 10304 2157 10368
rect 2221 10304 2229 10368
rect 1909 9280 2229 10304
rect 1909 9216 1917 9280
rect 1981 9216 1997 9280
rect 2061 9216 2077 9280
rect 2141 9216 2157 9280
rect 2221 9216 2229 9280
rect 1909 8192 2229 9216
rect 1909 8128 1917 8192
rect 1981 8128 1997 8192
rect 2061 8128 2077 8192
rect 2141 8128 2157 8192
rect 2221 8128 2229 8192
rect 1909 7104 2229 8128
rect 1909 7040 1917 7104
rect 1981 7040 1997 7104
rect 2061 7040 2077 7104
rect 2141 7040 2157 7104
rect 2221 7040 2229 7104
rect 1909 6016 2229 7040
rect 1909 5952 1917 6016
rect 1981 5952 1997 6016
rect 2061 5952 2077 6016
rect 2141 5952 2157 6016
rect 2221 5952 2229 6016
rect 1909 4928 2229 5952
rect 1909 4864 1917 4928
rect 1981 4864 1997 4928
rect 2061 4864 2077 4928
rect 2141 4864 2157 4928
rect 2221 4864 2229 4928
rect 1909 3840 2229 4864
rect 1909 3776 1917 3840
rect 1981 3776 1997 3840
rect 2061 3776 2077 3840
rect 2141 3776 2157 3840
rect 2221 3776 2229 3840
rect 1909 2752 2229 3776
rect 1909 2688 1917 2752
rect 1981 2688 1997 2752
rect 2061 2688 2077 2752
rect 2141 2688 2157 2752
rect 2221 2688 2229 2752
rect 1909 2128 2229 2688
rect 2874 30496 3194 31520
rect 2874 30432 2882 30496
rect 2946 30432 2962 30496
rect 3026 30432 3042 30496
rect 3106 30432 3122 30496
rect 3186 30432 3194 30496
rect 2874 29408 3194 30432
rect 3374 29885 3434 38251
rect 3558 31789 3618 42059
rect 3839 41920 4160 42944
rect 3839 41856 3848 41920
rect 3912 41856 3928 41920
rect 3992 41856 4008 41920
rect 4072 41856 4088 41920
rect 4152 41856 4160 41920
rect 3839 40832 4160 41856
rect 3839 40768 3848 40832
rect 3912 40768 3928 40832
rect 3992 40768 4008 40832
rect 4072 40768 4088 40832
rect 4152 40768 4160 40832
rect 3839 39744 4160 40768
rect 3839 39680 3848 39744
rect 3912 39680 3928 39744
rect 3992 39680 4008 39744
rect 4072 39680 4088 39744
rect 4152 39680 4160 39744
rect 3839 38656 4160 39680
rect 3839 38592 3848 38656
rect 3912 38592 3928 38656
rect 3992 38592 4008 38656
rect 4072 38592 4088 38656
rect 4152 38592 4160 38656
rect 3839 37568 4160 38592
rect 3839 37504 3848 37568
rect 3912 37504 3928 37568
rect 3992 37504 4008 37568
rect 4072 37504 4088 37568
rect 4152 37504 4160 37568
rect 3839 36480 4160 37504
rect 3839 36416 3848 36480
rect 3912 36416 3928 36480
rect 3992 36416 4008 36480
rect 4072 36416 4088 36480
rect 4152 36416 4160 36480
rect 3839 35392 4160 36416
rect 3839 35328 3848 35392
rect 3912 35328 3928 35392
rect 3992 35328 4008 35392
rect 4072 35328 4088 35392
rect 4152 35328 4160 35392
rect 3839 34304 4160 35328
rect 3839 34240 3848 34304
rect 3912 34240 3928 34304
rect 3992 34240 4008 34304
rect 4072 34240 4088 34304
rect 4152 34240 4160 34304
rect 3839 33216 4160 34240
rect 3839 33152 3848 33216
rect 3912 33152 3928 33216
rect 3992 33152 4008 33216
rect 4072 33152 4088 33216
rect 4152 33152 4160 33216
rect 3839 32128 4160 33152
rect 4294 32877 4354 55251
rect 4805 54432 5125 55456
rect 4805 54368 4813 54432
rect 4877 54368 4893 54432
rect 4957 54368 4973 54432
rect 5037 54368 5053 54432
rect 5117 54368 5125 54432
rect 4805 53344 5125 54368
rect 4805 53280 4813 53344
rect 4877 53280 4893 53344
rect 4957 53280 4973 53344
rect 5037 53280 5053 53344
rect 5117 53280 5125 53344
rect 4805 52256 5125 53280
rect 4805 52192 4813 52256
rect 4877 52192 4893 52256
rect 4957 52192 4973 52256
rect 5037 52192 5053 52256
rect 5117 52192 5125 52256
rect 4805 51168 5125 52192
rect 4805 51104 4813 51168
rect 4877 51104 4893 51168
rect 4957 51104 4973 51168
rect 5037 51104 5053 51168
rect 5117 51104 5125 51168
rect 4805 50080 5125 51104
rect 4805 50016 4813 50080
rect 4877 50016 4893 50080
rect 4957 50016 4973 50080
rect 5037 50016 5053 50080
rect 5117 50016 5125 50080
rect 4805 48992 5125 50016
rect 4805 48928 4813 48992
rect 4877 48928 4893 48992
rect 4957 48928 4973 48992
rect 5037 48928 5053 48992
rect 5117 48928 5125 48992
rect 4805 47904 5125 48928
rect 5770 57152 6090 57712
rect 5770 57088 5778 57152
rect 5842 57088 5858 57152
rect 5922 57088 5938 57152
rect 6002 57088 6018 57152
rect 6082 57088 6090 57152
rect 5770 56064 6090 57088
rect 5770 56000 5778 56064
rect 5842 56000 5858 56064
rect 5922 56000 5938 56064
rect 6002 56000 6018 56064
rect 6082 56000 6090 56064
rect 5770 54976 6090 56000
rect 5770 54912 5778 54976
rect 5842 54912 5858 54976
rect 5922 54912 5938 54976
rect 6002 54912 6018 54976
rect 6082 54912 6090 54976
rect 5770 53888 6090 54912
rect 5770 53824 5778 53888
rect 5842 53824 5858 53888
rect 5922 53824 5938 53888
rect 6002 53824 6018 53888
rect 6082 53824 6090 53888
rect 5770 52800 6090 53824
rect 5770 52736 5778 52800
rect 5842 52736 5858 52800
rect 5922 52736 5938 52800
rect 6002 52736 6018 52800
rect 6082 52736 6090 52800
rect 5770 51712 6090 52736
rect 5770 51648 5778 51712
rect 5842 51648 5858 51712
rect 5922 51648 5938 51712
rect 6002 51648 6018 51712
rect 6082 51648 6090 51712
rect 5770 50624 6090 51648
rect 5770 50560 5778 50624
rect 5842 50560 5858 50624
rect 5922 50560 5938 50624
rect 6002 50560 6018 50624
rect 6082 50560 6090 50624
rect 5770 49536 6090 50560
rect 5770 49472 5778 49536
rect 5842 49472 5858 49536
rect 5922 49472 5938 49536
rect 6002 49472 6018 49536
rect 6082 49472 6090 49536
rect 5770 48448 6090 49472
rect 5770 48384 5778 48448
rect 5842 48384 5858 48448
rect 5922 48384 5938 48448
rect 6002 48384 6018 48448
rect 6082 48384 6090 48448
rect 5395 48108 5461 48109
rect 5395 48044 5396 48108
rect 5460 48044 5461 48108
rect 5395 48043 5461 48044
rect 4805 47840 4813 47904
rect 4877 47840 4893 47904
rect 4957 47840 4973 47904
rect 5037 47840 5053 47904
rect 5117 47840 5125 47904
rect 4659 47836 4725 47837
rect 4659 47772 4660 47836
rect 4724 47772 4725 47836
rect 4659 47771 4725 47772
rect 4662 42261 4722 47771
rect 4805 46816 5125 47840
rect 4805 46752 4813 46816
rect 4877 46752 4893 46816
rect 4957 46752 4973 46816
rect 5037 46752 5053 46816
rect 5117 46752 5125 46816
rect 4805 45728 5125 46752
rect 4805 45664 4813 45728
rect 4877 45664 4893 45728
rect 4957 45664 4973 45728
rect 5037 45664 5053 45728
rect 5117 45664 5125 45728
rect 4805 44640 5125 45664
rect 5211 45388 5277 45389
rect 5211 45324 5212 45388
rect 5276 45324 5277 45388
rect 5211 45323 5277 45324
rect 4805 44576 4813 44640
rect 4877 44576 4893 44640
rect 4957 44576 4973 44640
rect 5037 44576 5053 44640
rect 5117 44576 5125 44640
rect 4805 43552 5125 44576
rect 4805 43488 4813 43552
rect 4877 43488 4893 43552
rect 4957 43488 4973 43552
rect 5037 43488 5053 43552
rect 5117 43488 5125 43552
rect 4805 42464 5125 43488
rect 4805 42400 4813 42464
rect 4877 42400 4893 42464
rect 4957 42400 4973 42464
rect 5037 42400 5053 42464
rect 5117 42400 5125 42464
rect 4659 42260 4725 42261
rect 4659 42196 4660 42260
rect 4724 42196 4725 42260
rect 4659 42195 4725 42196
rect 4659 41988 4725 41989
rect 4659 41924 4660 41988
rect 4724 41924 4725 41988
rect 4659 41923 4725 41924
rect 4475 41852 4541 41853
rect 4475 41788 4476 41852
rect 4540 41788 4541 41852
rect 4475 41787 4541 41788
rect 4478 41170 4538 41787
rect 4662 41309 4722 41923
rect 4805 41376 5125 42400
rect 4805 41312 4813 41376
rect 4877 41312 4893 41376
rect 4957 41312 4973 41376
rect 5037 41312 5053 41376
rect 5117 41312 5125 41376
rect 4659 41308 4725 41309
rect 4659 41244 4660 41308
rect 4724 41244 4725 41308
rect 4659 41243 4725 41244
rect 4478 41110 4722 41170
rect 4475 41036 4541 41037
rect 4475 40972 4476 41036
rect 4540 40972 4541 41036
rect 4475 40971 4541 40972
rect 4478 34509 4538 40971
rect 4475 34508 4541 34509
rect 4475 34444 4476 34508
rect 4540 34444 4541 34508
rect 4475 34443 4541 34444
rect 4291 32876 4357 32877
rect 4291 32812 4292 32876
rect 4356 32812 4357 32876
rect 4291 32811 4357 32812
rect 4662 32333 4722 41110
rect 4805 40288 5125 41312
rect 5214 40901 5274 45323
rect 5398 41717 5458 48043
rect 5770 47360 6090 48384
rect 5770 47296 5778 47360
rect 5842 47296 5858 47360
rect 5922 47296 5938 47360
rect 6002 47296 6018 47360
rect 6082 47296 6090 47360
rect 5770 46272 6090 47296
rect 5770 46208 5778 46272
rect 5842 46208 5858 46272
rect 5922 46208 5938 46272
rect 6002 46208 6018 46272
rect 6082 46208 6090 46272
rect 5770 45184 6090 46208
rect 5770 45120 5778 45184
rect 5842 45120 5858 45184
rect 5922 45120 5938 45184
rect 6002 45120 6018 45184
rect 6082 45120 6090 45184
rect 5770 44096 6090 45120
rect 5770 44032 5778 44096
rect 5842 44032 5858 44096
rect 5922 44032 5938 44096
rect 6002 44032 6018 44096
rect 6082 44032 6090 44096
rect 5579 43348 5645 43349
rect 5579 43284 5580 43348
rect 5644 43284 5645 43348
rect 5579 43283 5645 43284
rect 5395 41716 5461 41717
rect 5395 41652 5396 41716
rect 5460 41652 5461 41716
rect 5395 41651 5461 41652
rect 5211 40900 5277 40901
rect 5211 40836 5212 40900
rect 5276 40836 5277 40900
rect 5211 40835 5277 40836
rect 4805 40224 4813 40288
rect 4877 40224 4893 40288
rect 4957 40224 4973 40288
rect 5037 40224 5053 40288
rect 5117 40224 5125 40288
rect 4805 39200 5125 40224
rect 4805 39136 4813 39200
rect 4877 39136 4893 39200
rect 4957 39136 4973 39200
rect 5037 39136 5053 39200
rect 5117 39136 5125 39200
rect 4805 38112 5125 39136
rect 5582 38997 5642 43283
rect 5770 43008 6090 44032
rect 5770 42944 5778 43008
rect 5842 42944 5858 43008
rect 5922 42944 5938 43008
rect 6002 42944 6018 43008
rect 6082 42944 6090 43008
rect 5770 41920 6090 42944
rect 5770 41856 5778 41920
rect 5842 41856 5858 41920
rect 5922 41856 5938 41920
rect 6002 41856 6018 41920
rect 6082 41856 6090 41920
rect 5770 40832 6090 41856
rect 5770 40768 5778 40832
rect 5842 40768 5858 40832
rect 5922 40768 5938 40832
rect 6002 40768 6018 40832
rect 6082 40768 6090 40832
rect 5770 39744 6090 40768
rect 5770 39680 5778 39744
rect 5842 39680 5858 39744
rect 5922 39680 5938 39744
rect 6002 39680 6018 39744
rect 6082 39680 6090 39744
rect 5579 38996 5645 38997
rect 5579 38932 5580 38996
rect 5644 38932 5645 38996
rect 5579 38931 5645 38932
rect 4805 38048 4813 38112
rect 4877 38048 4893 38112
rect 4957 38048 4973 38112
rect 5037 38048 5053 38112
rect 5117 38048 5125 38112
rect 4805 37024 5125 38048
rect 4805 36960 4813 37024
rect 4877 36960 4893 37024
rect 4957 36960 4973 37024
rect 5037 36960 5053 37024
rect 5117 36960 5125 37024
rect 4805 35936 5125 36960
rect 4805 35872 4813 35936
rect 4877 35872 4893 35936
rect 4957 35872 4973 35936
rect 5037 35872 5053 35936
rect 5117 35872 5125 35936
rect 4805 34848 5125 35872
rect 4805 34784 4813 34848
rect 4877 34784 4893 34848
rect 4957 34784 4973 34848
rect 5037 34784 5053 34848
rect 5117 34784 5125 34848
rect 4805 33760 5125 34784
rect 4805 33696 4813 33760
rect 4877 33696 4893 33760
rect 4957 33696 4973 33760
rect 5037 33696 5053 33760
rect 5117 33696 5125 33760
rect 4805 32672 5125 33696
rect 4805 32608 4813 32672
rect 4877 32608 4893 32672
rect 4957 32608 4973 32672
rect 5037 32608 5053 32672
rect 5117 32608 5125 32672
rect 4659 32332 4725 32333
rect 4659 32268 4660 32332
rect 4724 32268 4725 32332
rect 4659 32267 4725 32268
rect 3839 32064 3848 32128
rect 3912 32064 3928 32128
rect 3992 32064 4008 32128
rect 4072 32064 4088 32128
rect 4152 32064 4160 32128
rect 3555 31788 3621 31789
rect 3555 31724 3556 31788
rect 3620 31724 3621 31788
rect 3555 31723 3621 31724
rect 3839 31040 4160 32064
rect 3839 30976 3848 31040
rect 3912 30976 3928 31040
rect 3992 30976 4008 31040
rect 4072 30976 4088 31040
rect 4152 30976 4160 31040
rect 3839 29952 4160 30976
rect 3839 29888 3848 29952
rect 3912 29888 3928 29952
rect 3992 29888 4008 29952
rect 4072 29888 4088 29952
rect 4152 29888 4160 29952
rect 3371 29884 3437 29885
rect 3371 29820 3372 29884
rect 3436 29820 3437 29884
rect 3371 29819 3437 29820
rect 2874 29344 2882 29408
rect 2946 29344 2962 29408
rect 3026 29344 3042 29408
rect 3106 29344 3122 29408
rect 3186 29344 3194 29408
rect 2874 28320 3194 29344
rect 2874 28256 2882 28320
rect 2946 28256 2962 28320
rect 3026 28256 3042 28320
rect 3106 28256 3122 28320
rect 3186 28256 3194 28320
rect 2874 27232 3194 28256
rect 2874 27168 2882 27232
rect 2946 27168 2962 27232
rect 3026 27168 3042 27232
rect 3106 27168 3122 27232
rect 3186 27168 3194 27232
rect 2874 26144 3194 27168
rect 2874 26080 2882 26144
rect 2946 26080 2962 26144
rect 3026 26080 3042 26144
rect 3106 26080 3122 26144
rect 3186 26080 3194 26144
rect 2874 25056 3194 26080
rect 2874 24992 2882 25056
rect 2946 24992 2962 25056
rect 3026 24992 3042 25056
rect 3106 24992 3122 25056
rect 3186 24992 3194 25056
rect 2874 23968 3194 24992
rect 2874 23904 2882 23968
rect 2946 23904 2962 23968
rect 3026 23904 3042 23968
rect 3106 23904 3122 23968
rect 3186 23904 3194 23968
rect 2874 22880 3194 23904
rect 2874 22816 2882 22880
rect 2946 22816 2962 22880
rect 3026 22816 3042 22880
rect 3106 22816 3122 22880
rect 3186 22816 3194 22880
rect 2874 21792 3194 22816
rect 2874 21728 2882 21792
rect 2946 21728 2962 21792
rect 3026 21728 3042 21792
rect 3106 21728 3122 21792
rect 3186 21728 3194 21792
rect 2874 20704 3194 21728
rect 2874 20640 2882 20704
rect 2946 20640 2962 20704
rect 3026 20640 3042 20704
rect 3106 20640 3122 20704
rect 3186 20640 3194 20704
rect 2874 19616 3194 20640
rect 2874 19552 2882 19616
rect 2946 19552 2962 19616
rect 3026 19552 3042 19616
rect 3106 19552 3122 19616
rect 3186 19552 3194 19616
rect 2874 18528 3194 19552
rect 2874 18464 2882 18528
rect 2946 18464 2962 18528
rect 3026 18464 3042 18528
rect 3106 18464 3122 18528
rect 3186 18464 3194 18528
rect 2874 17440 3194 18464
rect 2874 17376 2882 17440
rect 2946 17376 2962 17440
rect 3026 17376 3042 17440
rect 3106 17376 3122 17440
rect 3186 17376 3194 17440
rect 2874 16352 3194 17376
rect 2874 16288 2882 16352
rect 2946 16288 2962 16352
rect 3026 16288 3042 16352
rect 3106 16288 3122 16352
rect 3186 16288 3194 16352
rect 2874 15264 3194 16288
rect 2874 15200 2882 15264
rect 2946 15200 2962 15264
rect 3026 15200 3042 15264
rect 3106 15200 3122 15264
rect 3186 15200 3194 15264
rect 2874 14176 3194 15200
rect 2874 14112 2882 14176
rect 2946 14112 2962 14176
rect 3026 14112 3042 14176
rect 3106 14112 3122 14176
rect 3186 14112 3194 14176
rect 2874 13088 3194 14112
rect 2874 13024 2882 13088
rect 2946 13024 2962 13088
rect 3026 13024 3042 13088
rect 3106 13024 3122 13088
rect 3186 13024 3194 13088
rect 2874 12000 3194 13024
rect 2874 11936 2882 12000
rect 2946 11936 2962 12000
rect 3026 11936 3042 12000
rect 3106 11936 3122 12000
rect 3186 11936 3194 12000
rect 2874 10912 3194 11936
rect 2874 10848 2882 10912
rect 2946 10848 2962 10912
rect 3026 10848 3042 10912
rect 3106 10848 3122 10912
rect 3186 10848 3194 10912
rect 2874 9824 3194 10848
rect 2874 9760 2882 9824
rect 2946 9760 2962 9824
rect 3026 9760 3042 9824
rect 3106 9760 3122 9824
rect 3186 9760 3194 9824
rect 2874 8736 3194 9760
rect 2874 8672 2882 8736
rect 2946 8672 2962 8736
rect 3026 8672 3042 8736
rect 3106 8672 3122 8736
rect 3186 8672 3194 8736
rect 2874 7648 3194 8672
rect 2874 7584 2882 7648
rect 2946 7584 2962 7648
rect 3026 7584 3042 7648
rect 3106 7584 3122 7648
rect 3186 7584 3194 7648
rect 2874 6560 3194 7584
rect 2874 6496 2882 6560
rect 2946 6496 2962 6560
rect 3026 6496 3042 6560
rect 3106 6496 3122 6560
rect 3186 6496 3194 6560
rect 2874 5472 3194 6496
rect 2874 5408 2882 5472
rect 2946 5408 2962 5472
rect 3026 5408 3042 5472
rect 3106 5408 3122 5472
rect 3186 5408 3194 5472
rect 2874 4384 3194 5408
rect 2874 4320 2882 4384
rect 2946 4320 2962 4384
rect 3026 4320 3042 4384
rect 3106 4320 3122 4384
rect 3186 4320 3194 4384
rect 2874 3296 3194 4320
rect 2874 3232 2882 3296
rect 2946 3232 2962 3296
rect 3026 3232 3042 3296
rect 3106 3232 3122 3296
rect 3186 3232 3194 3296
rect 2874 2208 3194 3232
rect 2874 2144 2882 2208
rect 2946 2144 2962 2208
rect 3026 2144 3042 2208
rect 3106 2144 3122 2208
rect 3186 2144 3194 2208
rect 2874 2128 3194 2144
rect 3839 28864 4160 29888
rect 3839 28800 3848 28864
rect 3912 28800 3928 28864
rect 3992 28800 4008 28864
rect 4072 28800 4088 28864
rect 4152 28800 4160 28864
rect 3839 27776 4160 28800
rect 3839 27712 3848 27776
rect 3912 27712 3928 27776
rect 3992 27712 4008 27776
rect 4072 27712 4088 27776
rect 4152 27712 4160 27776
rect 3839 26688 4160 27712
rect 3839 26624 3848 26688
rect 3912 26624 3928 26688
rect 3992 26624 4008 26688
rect 4072 26624 4088 26688
rect 4152 26624 4160 26688
rect 3839 25600 4160 26624
rect 3839 25536 3848 25600
rect 3912 25536 3928 25600
rect 3992 25536 4008 25600
rect 4072 25536 4088 25600
rect 4152 25536 4160 25600
rect 3839 24512 4160 25536
rect 3839 24448 3848 24512
rect 3912 24448 3928 24512
rect 3992 24448 4008 24512
rect 4072 24448 4088 24512
rect 4152 24448 4160 24512
rect 3839 23424 4160 24448
rect 3839 23360 3848 23424
rect 3912 23360 3928 23424
rect 3992 23360 4008 23424
rect 4072 23360 4088 23424
rect 4152 23360 4160 23424
rect 3839 22336 4160 23360
rect 3839 22272 3848 22336
rect 3912 22272 3928 22336
rect 3992 22272 4008 22336
rect 4072 22272 4088 22336
rect 4152 22272 4160 22336
rect 3839 21248 4160 22272
rect 3839 21184 3848 21248
rect 3912 21184 3928 21248
rect 3992 21184 4008 21248
rect 4072 21184 4088 21248
rect 4152 21184 4160 21248
rect 3839 20160 4160 21184
rect 3839 20096 3848 20160
rect 3912 20096 3928 20160
rect 3992 20096 4008 20160
rect 4072 20096 4088 20160
rect 4152 20096 4160 20160
rect 3839 19072 4160 20096
rect 3839 19008 3848 19072
rect 3912 19008 3928 19072
rect 3992 19008 4008 19072
rect 4072 19008 4088 19072
rect 4152 19008 4160 19072
rect 3839 17984 4160 19008
rect 3839 17920 3848 17984
rect 3912 17920 3928 17984
rect 3992 17920 4008 17984
rect 4072 17920 4088 17984
rect 4152 17920 4160 17984
rect 3839 16896 4160 17920
rect 3839 16832 3848 16896
rect 3912 16832 3928 16896
rect 3992 16832 4008 16896
rect 4072 16832 4088 16896
rect 4152 16832 4160 16896
rect 3839 15808 4160 16832
rect 3839 15744 3848 15808
rect 3912 15744 3928 15808
rect 3992 15744 4008 15808
rect 4072 15744 4088 15808
rect 4152 15744 4160 15808
rect 3839 14720 4160 15744
rect 3839 14656 3848 14720
rect 3912 14656 3928 14720
rect 3992 14656 4008 14720
rect 4072 14656 4088 14720
rect 4152 14656 4160 14720
rect 3839 13632 4160 14656
rect 3839 13568 3848 13632
rect 3912 13568 3928 13632
rect 3992 13568 4008 13632
rect 4072 13568 4088 13632
rect 4152 13568 4160 13632
rect 3839 12544 4160 13568
rect 3839 12480 3848 12544
rect 3912 12480 3928 12544
rect 3992 12480 4008 12544
rect 4072 12480 4088 12544
rect 4152 12480 4160 12544
rect 3839 11456 4160 12480
rect 3839 11392 3848 11456
rect 3912 11392 3928 11456
rect 3992 11392 4008 11456
rect 4072 11392 4088 11456
rect 4152 11392 4160 11456
rect 3839 10368 4160 11392
rect 3839 10304 3848 10368
rect 3912 10304 3928 10368
rect 3992 10304 4008 10368
rect 4072 10304 4088 10368
rect 4152 10304 4160 10368
rect 3839 9280 4160 10304
rect 3839 9216 3848 9280
rect 3912 9216 3928 9280
rect 3992 9216 4008 9280
rect 4072 9216 4088 9280
rect 4152 9216 4160 9280
rect 3839 8192 4160 9216
rect 3839 8128 3848 8192
rect 3912 8128 3928 8192
rect 3992 8128 4008 8192
rect 4072 8128 4088 8192
rect 4152 8128 4160 8192
rect 3839 7104 4160 8128
rect 3839 7040 3848 7104
rect 3912 7040 3928 7104
rect 3992 7040 4008 7104
rect 4072 7040 4088 7104
rect 4152 7040 4160 7104
rect 3839 6016 4160 7040
rect 3839 5952 3848 6016
rect 3912 5952 3928 6016
rect 3992 5952 4008 6016
rect 4072 5952 4088 6016
rect 4152 5952 4160 6016
rect 3839 4928 4160 5952
rect 3839 4864 3848 4928
rect 3912 4864 3928 4928
rect 3992 4864 4008 4928
rect 4072 4864 4088 4928
rect 4152 4864 4160 4928
rect 3839 3840 4160 4864
rect 3839 3776 3848 3840
rect 3912 3776 3928 3840
rect 3992 3776 4008 3840
rect 4072 3776 4088 3840
rect 4152 3776 4160 3840
rect 3839 2752 4160 3776
rect 3839 2688 3848 2752
rect 3912 2688 3928 2752
rect 3992 2688 4008 2752
rect 4072 2688 4088 2752
rect 4152 2688 4160 2752
rect 3839 2128 4160 2688
rect 4805 31584 5125 32608
rect 4805 31520 4813 31584
rect 4877 31520 4893 31584
rect 4957 31520 4973 31584
rect 5037 31520 5053 31584
rect 5117 31520 5125 31584
rect 4805 30496 5125 31520
rect 4805 30432 4813 30496
rect 4877 30432 4893 30496
rect 4957 30432 4973 30496
rect 5037 30432 5053 30496
rect 5117 30432 5125 30496
rect 4805 29408 5125 30432
rect 4805 29344 4813 29408
rect 4877 29344 4893 29408
rect 4957 29344 4973 29408
rect 5037 29344 5053 29408
rect 5117 29344 5125 29408
rect 4805 28320 5125 29344
rect 4805 28256 4813 28320
rect 4877 28256 4893 28320
rect 4957 28256 4973 28320
rect 5037 28256 5053 28320
rect 5117 28256 5125 28320
rect 4805 27232 5125 28256
rect 4805 27168 4813 27232
rect 4877 27168 4893 27232
rect 4957 27168 4973 27232
rect 5037 27168 5053 27232
rect 5117 27168 5125 27232
rect 4805 26144 5125 27168
rect 4805 26080 4813 26144
rect 4877 26080 4893 26144
rect 4957 26080 4973 26144
rect 5037 26080 5053 26144
rect 5117 26080 5125 26144
rect 4805 25056 5125 26080
rect 4805 24992 4813 25056
rect 4877 24992 4893 25056
rect 4957 24992 4973 25056
rect 5037 24992 5053 25056
rect 5117 24992 5125 25056
rect 4805 23968 5125 24992
rect 4805 23904 4813 23968
rect 4877 23904 4893 23968
rect 4957 23904 4973 23968
rect 5037 23904 5053 23968
rect 5117 23904 5125 23968
rect 4805 22880 5125 23904
rect 4805 22816 4813 22880
rect 4877 22816 4893 22880
rect 4957 22816 4973 22880
rect 5037 22816 5053 22880
rect 5117 22816 5125 22880
rect 4805 21792 5125 22816
rect 4805 21728 4813 21792
rect 4877 21728 4893 21792
rect 4957 21728 4973 21792
rect 5037 21728 5053 21792
rect 5117 21728 5125 21792
rect 4805 20704 5125 21728
rect 4805 20640 4813 20704
rect 4877 20640 4893 20704
rect 4957 20640 4973 20704
rect 5037 20640 5053 20704
rect 5117 20640 5125 20704
rect 4805 19616 5125 20640
rect 4805 19552 4813 19616
rect 4877 19552 4893 19616
rect 4957 19552 4973 19616
rect 5037 19552 5053 19616
rect 5117 19552 5125 19616
rect 4805 18528 5125 19552
rect 4805 18464 4813 18528
rect 4877 18464 4893 18528
rect 4957 18464 4973 18528
rect 5037 18464 5053 18528
rect 5117 18464 5125 18528
rect 4805 17440 5125 18464
rect 4805 17376 4813 17440
rect 4877 17376 4893 17440
rect 4957 17376 4973 17440
rect 5037 17376 5053 17440
rect 5117 17376 5125 17440
rect 4805 16352 5125 17376
rect 4805 16288 4813 16352
rect 4877 16288 4893 16352
rect 4957 16288 4973 16352
rect 5037 16288 5053 16352
rect 5117 16288 5125 16352
rect 4805 15264 5125 16288
rect 4805 15200 4813 15264
rect 4877 15200 4893 15264
rect 4957 15200 4973 15264
rect 5037 15200 5053 15264
rect 5117 15200 5125 15264
rect 4805 14176 5125 15200
rect 4805 14112 4813 14176
rect 4877 14112 4893 14176
rect 4957 14112 4973 14176
rect 5037 14112 5053 14176
rect 5117 14112 5125 14176
rect 4805 13088 5125 14112
rect 4805 13024 4813 13088
rect 4877 13024 4893 13088
rect 4957 13024 4973 13088
rect 5037 13024 5053 13088
rect 5117 13024 5125 13088
rect 4805 12000 5125 13024
rect 4805 11936 4813 12000
rect 4877 11936 4893 12000
rect 4957 11936 4973 12000
rect 5037 11936 5053 12000
rect 5117 11936 5125 12000
rect 4805 10912 5125 11936
rect 4805 10848 4813 10912
rect 4877 10848 4893 10912
rect 4957 10848 4973 10912
rect 5037 10848 5053 10912
rect 5117 10848 5125 10912
rect 4805 9824 5125 10848
rect 4805 9760 4813 9824
rect 4877 9760 4893 9824
rect 4957 9760 4973 9824
rect 5037 9760 5053 9824
rect 5117 9760 5125 9824
rect 4805 8736 5125 9760
rect 4805 8672 4813 8736
rect 4877 8672 4893 8736
rect 4957 8672 4973 8736
rect 5037 8672 5053 8736
rect 5117 8672 5125 8736
rect 4805 7648 5125 8672
rect 4805 7584 4813 7648
rect 4877 7584 4893 7648
rect 4957 7584 4973 7648
rect 5037 7584 5053 7648
rect 5117 7584 5125 7648
rect 4805 6560 5125 7584
rect 4805 6496 4813 6560
rect 4877 6496 4893 6560
rect 4957 6496 4973 6560
rect 5037 6496 5053 6560
rect 5117 6496 5125 6560
rect 4805 5472 5125 6496
rect 4805 5408 4813 5472
rect 4877 5408 4893 5472
rect 4957 5408 4973 5472
rect 5037 5408 5053 5472
rect 5117 5408 5125 5472
rect 4805 4384 5125 5408
rect 4805 4320 4813 4384
rect 4877 4320 4893 4384
rect 4957 4320 4973 4384
rect 5037 4320 5053 4384
rect 5117 4320 5125 4384
rect 4805 3296 5125 4320
rect 4805 3232 4813 3296
rect 4877 3232 4893 3296
rect 4957 3232 4973 3296
rect 5037 3232 5053 3296
rect 5117 3232 5125 3296
rect 4805 2208 5125 3232
rect 4805 2144 4813 2208
rect 4877 2144 4893 2208
rect 4957 2144 4973 2208
rect 5037 2144 5053 2208
rect 5117 2144 5125 2208
rect 4805 2128 5125 2144
rect 5770 38656 6090 39680
rect 5770 38592 5778 38656
rect 5842 38592 5858 38656
rect 5922 38592 5938 38656
rect 6002 38592 6018 38656
rect 6082 38592 6090 38656
rect 5770 37568 6090 38592
rect 5770 37504 5778 37568
rect 5842 37504 5858 37568
rect 5922 37504 5938 37568
rect 6002 37504 6018 37568
rect 6082 37504 6090 37568
rect 5770 36480 6090 37504
rect 5770 36416 5778 36480
rect 5842 36416 5858 36480
rect 5922 36416 5938 36480
rect 6002 36416 6018 36480
rect 6082 36416 6090 36480
rect 5770 35392 6090 36416
rect 5770 35328 5778 35392
rect 5842 35328 5858 35392
rect 5922 35328 5938 35392
rect 6002 35328 6018 35392
rect 6082 35328 6090 35392
rect 5770 34304 6090 35328
rect 5770 34240 5778 34304
rect 5842 34240 5858 34304
rect 5922 34240 5938 34304
rect 6002 34240 6018 34304
rect 6082 34240 6090 34304
rect 5770 33216 6090 34240
rect 5770 33152 5778 33216
rect 5842 33152 5858 33216
rect 5922 33152 5938 33216
rect 6002 33152 6018 33216
rect 6082 33152 6090 33216
rect 5770 32128 6090 33152
rect 5770 32064 5778 32128
rect 5842 32064 5858 32128
rect 5922 32064 5938 32128
rect 6002 32064 6018 32128
rect 6082 32064 6090 32128
rect 5770 31040 6090 32064
rect 5770 30976 5778 31040
rect 5842 30976 5858 31040
rect 5922 30976 5938 31040
rect 6002 30976 6018 31040
rect 6082 30976 6090 31040
rect 5770 29952 6090 30976
rect 5770 29888 5778 29952
rect 5842 29888 5858 29952
rect 5922 29888 5938 29952
rect 6002 29888 6018 29952
rect 6082 29888 6090 29952
rect 5770 28864 6090 29888
rect 5770 28800 5778 28864
rect 5842 28800 5858 28864
rect 5922 28800 5938 28864
rect 6002 28800 6018 28864
rect 6082 28800 6090 28864
rect 5770 27776 6090 28800
rect 5770 27712 5778 27776
rect 5842 27712 5858 27776
rect 5922 27712 5938 27776
rect 6002 27712 6018 27776
rect 6082 27712 6090 27776
rect 5770 26688 6090 27712
rect 5770 26624 5778 26688
rect 5842 26624 5858 26688
rect 5922 26624 5938 26688
rect 6002 26624 6018 26688
rect 6082 26624 6090 26688
rect 5770 25600 6090 26624
rect 5770 25536 5778 25600
rect 5842 25536 5858 25600
rect 5922 25536 5938 25600
rect 6002 25536 6018 25600
rect 6082 25536 6090 25600
rect 5770 24512 6090 25536
rect 5770 24448 5778 24512
rect 5842 24448 5858 24512
rect 5922 24448 5938 24512
rect 6002 24448 6018 24512
rect 6082 24448 6090 24512
rect 5770 23424 6090 24448
rect 5770 23360 5778 23424
rect 5842 23360 5858 23424
rect 5922 23360 5938 23424
rect 6002 23360 6018 23424
rect 6082 23360 6090 23424
rect 5770 22336 6090 23360
rect 5770 22272 5778 22336
rect 5842 22272 5858 22336
rect 5922 22272 5938 22336
rect 6002 22272 6018 22336
rect 6082 22272 6090 22336
rect 5770 21248 6090 22272
rect 5770 21184 5778 21248
rect 5842 21184 5858 21248
rect 5922 21184 5938 21248
rect 6002 21184 6018 21248
rect 6082 21184 6090 21248
rect 5770 20160 6090 21184
rect 5770 20096 5778 20160
rect 5842 20096 5858 20160
rect 5922 20096 5938 20160
rect 6002 20096 6018 20160
rect 6082 20096 6090 20160
rect 5770 19072 6090 20096
rect 5770 19008 5778 19072
rect 5842 19008 5858 19072
rect 5922 19008 5938 19072
rect 6002 19008 6018 19072
rect 6082 19008 6090 19072
rect 5770 17984 6090 19008
rect 5770 17920 5778 17984
rect 5842 17920 5858 17984
rect 5922 17920 5938 17984
rect 6002 17920 6018 17984
rect 6082 17920 6090 17984
rect 5770 16896 6090 17920
rect 5770 16832 5778 16896
rect 5842 16832 5858 16896
rect 5922 16832 5938 16896
rect 6002 16832 6018 16896
rect 6082 16832 6090 16896
rect 5770 15808 6090 16832
rect 5770 15744 5778 15808
rect 5842 15744 5858 15808
rect 5922 15744 5938 15808
rect 6002 15744 6018 15808
rect 6082 15744 6090 15808
rect 5770 14720 6090 15744
rect 5770 14656 5778 14720
rect 5842 14656 5858 14720
rect 5922 14656 5938 14720
rect 6002 14656 6018 14720
rect 6082 14656 6090 14720
rect 5770 13632 6090 14656
rect 5770 13568 5778 13632
rect 5842 13568 5858 13632
rect 5922 13568 5938 13632
rect 6002 13568 6018 13632
rect 6082 13568 6090 13632
rect 5770 12544 6090 13568
rect 5770 12480 5778 12544
rect 5842 12480 5858 12544
rect 5922 12480 5938 12544
rect 6002 12480 6018 12544
rect 6082 12480 6090 12544
rect 5770 11456 6090 12480
rect 5770 11392 5778 11456
rect 5842 11392 5858 11456
rect 5922 11392 5938 11456
rect 6002 11392 6018 11456
rect 6082 11392 6090 11456
rect 5770 10368 6090 11392
rect 5770 10304 5778 10368
rect 5842 10304 5858 10368
rect 5922 10304 5938 10368
rect 6002 10304 6018 10368
rect 6082 10304 6090 10368
rect 5770 9280 6090 10304
rect 5770 9216 5778 9280
rect 5842 9216 5858 9280
rect 5922 9216 5938 9280
rect 6002 9216 6018 9280
rect 6082 9216 6090 9280
rect 5770 8192 6090 9216
rect 5770 8128 5778 8192
rect 5842 8128 5858 8192
rect 5922 8128 5938 8192
rect 6002 8128 6018 8192
rect 6082 8128 6090 8192
rect 5770 7104 6090 8128
rect 5770 7040 5778 7104
rect 5842 7040 5858 7104
rect 5922 7040 5938 7104
rect 6002 7040 6018 7104
rect 6082 7040 6090 7104
rect 5770 6016 6090 7040
rect 5770 5952 5778 6016
rect 5842 5952 5858 6016
rect 5922 5952 5938 6016
rect 6002 5952 6018 6016
rect 6082 5952 6090 6016
rect 5770 4928 6090 5952
rect 5770 4864 5778 4928
rect 5842 4864 5858 4928
rect 5922 4864 5938 4928
rect 6002 4864 6018 4928
rect 6082 4864 6090 4928
rect 5770 3840 6090 4864
rect 5770 3776 5778 3840
rect 5842 3776 5858 3840
rect 5922 3776 5938 3840
rect 6002 3776 6018 3840
rect 6082 3776 6090 3840
rect 5770 2752 6090 3776
rect 5770 2688 5778 2752
rect 5842 2688 5858 2752
rect 5922 2688 5938 2752
rect 6002 2688 6018 2752
rect 6082 2688 6090 2752
rect 5770 2128 6090 2688
use sky130_fd_sc_hd__decap_12  FILLER_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1635330089
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_7
timestamp 1635330089
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635330089
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output114 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1635330089
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1635330089
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23
timestamp 1635330089
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_28
timestamp 1635330089
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1635330089
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1635330089
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1635330089
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1635330089
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1635330089
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635330089
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1635330089
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1635330089
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1635330089
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1635330089
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1635330089
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635330089
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635330089
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1635330089
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1635330089
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_7
timestamp 1635330089
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635330089
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1635330089
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1635330089
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1635330089
transform 1 0 4600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1635330089
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1635330089
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_45
timestamp 1635330089
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1635330089
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635330089
transform -1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1635330089
transform 1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1635330089
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1635330089
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1635330089
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635330089
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1635330089
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1635330089
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1635330089
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1635330089
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1635330089
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1635330089
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1635330089
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_42
timestamp 1635330089
transform 1 0 4968 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp 1635330089
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1635330089
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1635330089
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635330089
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1635330089
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp 1635330089
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1635330089
transform 1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 1635330089
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1635330089
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635330089
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _030_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _041_
timestamp 1635330089
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1635330089
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1635330089
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_35
timestamp 1635330089
transform 1 0 4324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1635330089
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _027_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1635330089
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1635330089
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_55
timestamp 1635330089
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635330089
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _019_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 5336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_14
timestamp 1635330089
transform 1 0 2392 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1635330089
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635330089
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1635330089
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1635330089
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_22
timestamp 1635330089
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_28
timestamp 1635330089
transform 1 0 3680 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 4416 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1635330089
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1635330089
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1635330089
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635330089
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1635330089
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_19
timestamp 1635330089
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1635330089
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1635330089
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1635330089
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635330089
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635330089
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1635330089
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1635330089
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1635330089
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1635330089
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1635330089
transform 1 0 3864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_22
timestamp 1635330089
transform 1 0 3128 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1635330089
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1635330089
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _025__1
timestamp 1635330089
transform 1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1635330089
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1635330089
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 4140 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp 1635330089
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1635330089
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1635330089
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635330089
transform -1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635330089
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1635330089
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1635330089
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1635330089
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_7
timestamp 1635330089
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635330089
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1635330089
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635330089
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1635330089
transform 1 0 4048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1635330089
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1635330089
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1635330089
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_44
timestamp 1635330089
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1635330089
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_58
timestamp 1635330089
transform 1 0 6440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635330089
transform -1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _028_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 5520 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_19
timestamp 1635330089
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_7
timestamp 1635330089
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635330089
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1635330089
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 1635330089
transform 1 0 3404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1635330089
transform 1 0 4048 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_39
timestamp 1635330089
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _032_
timestamp 1635330089
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1635330089
transform 1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  net99_2
timestamp 1635330089
transform 1 0 3772 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 1635330089
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1635330089
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1635330089
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635330089
transform -1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1635330089
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _026_
timestamp 1635330089
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1635330089
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1635330089
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635330089
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1635330089
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1635330089
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1635330089
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_37
timestamp 1635330089
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1635330089
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1635330089
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1635330089
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1635330089
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1635330089
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635330089
transform -1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _024_
timestamp 1635330089
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1635330089
transform 1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1635330089
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1635330089
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635330089
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_30
timestamp 1635330089
transform 1 0 3864 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1635330089
transform 1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _111_
timestamp 1635330089
transform 1 0 4416 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1635330089
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1635330089
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635330089
transform -1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1635330089
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_14
timestamp 1635330089
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1635330089
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635330089
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1635330089
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1635330089
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1635330089
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1635330089
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1635330089
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1635330089
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1635330089
transform 1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1635330089
transform 1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635330089
transform -1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1635330089
transform 1 0 5888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1635330089
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_19
timestamp 1635330089
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_7
timestamp 1635330089
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1635330089
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1635330089
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635330089
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635330089
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1635330089
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_31
timestamp 1635330089
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1635330089
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1635330089
transform 1 0 4048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_40
timestamp 1635330089
transform 1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1635330089
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp 1635330089
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1635330089
transform 1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1635330089
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1635330089
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_45
timestamp 1635330089
transform 1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_48
timestamp 1635330089
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_43
timestamp 1635330089
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1635330089
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635330089
transform -1 0 6808 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635330089
transform -1 0 6808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1635330089
transform 1 0 6440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_52
timestamp 1635330089
transform 1 0 5888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1635330089
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_19
timestamp 1635330089
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_7
timestamp 1635330089
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635330089
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1635330089
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_31
timestamp 1635330089
transform 1 0 3956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_37
timestamp 1635330089
transform 1 0 4508 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1635330089
transform 1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1635330089
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1635330089
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635330089
transform -1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1635330089
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1635330089
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1635330089
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1635330089
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635330089
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1635330089
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1635330089
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1635330089
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1635330089
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1635330089
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1635330089
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1635330089
transform 1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_48
timestamp 1635330089
transform 1 0 5520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1635330089
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635330089
transform -1 0 6808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1635330089
transform 1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635330089
transform 1 0 5244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_18
timestamp 1635330089
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_6
timestamp 1635330089
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635330089
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1635330089
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_30
timestamp 1635330089
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_42
timestamp 1635330089
transform 1 0 4968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1635330089
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1635330089
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635330089
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1635330089
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _018_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 5336 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1635330089
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1635330089
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635330089
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635330089
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1635330089
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 1635330089
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1635330089
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_49
timestamp 1635330089
transform 1 0 5612 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1635330089
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635330089
transform -1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635330089
transform 1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_18
timestamp 1635330089
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_6
timestamp 1635330089
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1635330089
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_6
timestamp 1635330089
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635330089
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635330089
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635330089
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1635330089
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_30
timestamp 1635330089
transform 1 0 3864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_38
timestamp 1635330089
transform 1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1635330089
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1635330089
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_37
timestamp 1635330089
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1635330089
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _078_
timestamp 1635330089
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1635330089
transform 1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_45
timestamp 1635330089
transform 1 0 5244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1635330089
transform 1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_49
timestamp 1635330089
transform 1 0 5612 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1635330089
transform 1 0 5888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1635330089
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1635330089
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1635330089
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635330089
transform -1 0 6808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635330089
transform -1 0 6808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1635330089
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_15
timestamp 1635330089
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1635330089
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635330089
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_25
timestamp 1635330089
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_37
timestamp 1635330089
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1635330089
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1635330089
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1635330089
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635330089
transform -1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1635330089
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635330089
transform 1 0 5612 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1635330089
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_6
timestamp 1635330089
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635330089
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1635330089
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1635330089
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1635330089
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1635330089
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1635330089
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_55
timestamp 1635330089
transform 1 0 6164 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635330089
transform -1 0 6808 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _021_
timestamp 1635330089
transform 1 0 5612 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_18
timestamp 1635330089
transform 1 0 2760 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_6
timestamp 1635330089
transform 1 0 1656 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635330089
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1635330089
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_30
timestamp 1635330089
transform 1 0 3864 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1635330089
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1635330089
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1635330089
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635330089
transform -1 0 6808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1635330089
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _022_
timestamp 1635330089
transform 1 0 5336 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1635330089
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_6
timestamp 1635330089
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635330089
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1635330089
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1635330089
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1635330089
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1635330089
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1635330089
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_48
timestamp 1635330089
transform 1 0 5520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1635330089
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635330089
transform -1 0 6808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635330089
transform 1 0 5888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635330089
transform 1 0 5244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1635330089
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1635330089
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635330089
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1635330089
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1635330089
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_43
timestamp 1635330089
transform 1 0 5060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1635330089
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1635330089
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635330089
transform -1 0 6808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1635330089
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635330089
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1635330089
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_6
timestamp 1635330089
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_18
timestamp 1635330089
transform 1 0 2760 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_6
timestamp 1635330089
transform 1 0 1656 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635330089
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635330089
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635330089
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635330089
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1635330089
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1635330089
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_37
timestamp 1635330089
transform 1 0 4508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_30
timestamp 1635330089
transform 1 0 3864 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_38
timestamp 1635330089
transform 1 0 4600 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1635330089
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1635330089
transform 1 0 4140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _084_
timestamp 1635330089
transform 1 0 4232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1635330089
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_46
timestamp 1635330089
transform 1 0 5336 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1635330089
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1635330089
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635330089
transform -1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635330089
transform -1 0 6808 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1635330089
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _020_
timestamp 1635330089
transform 1 0 5612 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635330089
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1635330089
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1635330089
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635330089
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1635330089
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1635330089
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_35
timestamp 1635330089
transform 1 0 4324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1635330089
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1635330089
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1635330089
transform 1 0 4416 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_44
timestamp 1635330089
transform 1 0 5152 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_48
timestamp 1635330089
transform 1 0 5520 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_55
timestamp 1635330089
transform 1 0 6164 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635330089
transform -1 0 6808 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1635330089
transform 1 0 5888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1635330089
transform 1 0 5244 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_18
timestamp 1635330089
transform 1 0 2760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_6
timestamp 1635330089
transform 1 0 1656 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635330089
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1635330089
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1635330089
transform 1 0 3864 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_42
timestamp 1635330089
transform 1 0 4968 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_48
timestamp 1635330089
transform 1 0 5520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1635330089
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1635330089
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635330089
transform -1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1635330089
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635330089
transform 1 0 5612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_18
timestamp 1635330089
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_6
timestamp 1635330089
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635330089
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1635330089
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1635330089
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1635330089
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1635330089
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1635330089
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_49
timestamp 1635330089
transform 1 0 5612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_55
timestamp 1635330089
transform 1 0 6164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635330089
transform -1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635330089
transform 1 0 5888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1635330089
transform 1 0 2760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_6
timestamp 1635330089
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635330089
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635330089
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_22
timestamp 1635330089
transform 1 0 3128 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1635330089
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_39
timestamp 1635330089
transform 1 0 4692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1635330089
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_47
timestamp 1635330089
transform 1 0 5428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1635330089
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1635330089
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635330089
transform -1 0 6808 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1635330089
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635330089
transform 1 0 5612 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1635330089
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1635330089
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635330089
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _085_
timestamp 1635330089
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1635330089
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1635330089
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1635330089
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_41
timestamp 1635330089
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1635330089
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_49
timestamp 1635330089
transform 1 0 5612 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_55
timestamp 1635330089
transform 1 0 6164 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635330089
transform -1 0 6808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635330089
transform 1 0 5888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_18
timestamp 1635330089
transform 1 0 2760 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_6
timestamp 1635330089
transform 1 0 1656 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_18
timestamp 1635330089
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_6
timestamp 1635330089
transform 1 0 1656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635330089
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635330089
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635330089
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635330089
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_30
timestamp 1635330089
transform 1 0 3864 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1635330089
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1635330089
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_41
timestamp 1635330089
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1635330089
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_48
timestamp 1635330089
transform 1 0 5520 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_42
timestamp 1635330089
transform 1 0 4968 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635330089
transform 1 0 5888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635330089
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_55
timestamp 1635330089
transform 1 0 6164 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_49
timestamp 1635330089
transform 1 0 5612 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1635330089
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1635330089
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635330089
transform -1 0 6808 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635330089
transform -1 0 6808 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1635330089
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1635330089
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1635330089
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635330089
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1635330089
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_39
timestamp 1635330089
transform 1 0 4692 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_47
timestamp 1635330089
transform 1 0 5428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1635330089
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1635330089
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635330089
transform -1 0 6808 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1635330089
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635330089
transform 1 0 5612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_18
timestamp 1635330089
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_6
timestamp 1635330089
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635330089
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635330089
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1635330089
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1635330089
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_35
timestamp 1635330089
transform 1 0 4324 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_40
timestamp 1635330089
transform 1 0 4784 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1635330089
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1635330089
transform 1 0 4416 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_48
timestamp 1635330089
transform 1 0 5520 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_55
timestamp 1635330089
transform 1 0 6164 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635330089
transform -1 0 6808 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _016_
timestamp 1635330089
transform 1 0 5612 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_18
timestamp 1635330089
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_6
timestamp 1635330089
transform 1 0 1656 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635330089
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635330089
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_30
timestamp 1635330089
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_45
timestamp 1635330089
transform 1 0 5244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1635330089
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1635330089
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635330089
transform -1 0 6808 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1635330089
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635330089
transform 1 0 5612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635330089
transform 1 0 4968 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_18
timestamp 1635330089
transform 1 0 2760 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_6
timestamp 1635330089
transform 1 0 1656 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635330089
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _087_
timestamp 1635330089
transform 1 0 2944 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635330089
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1635330089
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1635330089
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_37
timestamp 1635330089
transform 1 0 4508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1635330089
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _086_
timestamp 1635330089
transform 1 0 4140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1635330089
transform 1 0 4876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_44
timestamp 1635330089
transform 1 0 5152 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_55
timestamp 1635330089
transform 1 0 6164 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635330089
transform -1 0 6808 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _023_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 5520 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_39_18
timestamp 1635330089
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_6
timestamp 1635330089
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1635330089
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1635330089
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1635330089
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635330089
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635330089
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1635330089
transform 1 0 1472 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635330089
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_30
timestamp 1635330089
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1635330089
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1635330089
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_37
timestamp 1635330089
transform 1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1635330089
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1635330089
transform 1 0 4140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1635330089
transform 1 0 5244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _015_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 5152 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_48
timestamp 1635330089
transform 1 0 5520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_42
timestamp 1635330089
transform 1 0 4968 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635330089
transform 1 0 5888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1635330089
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635330089
transform -1 0 6808 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635330089
transform -1 0 6808 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_55
timestamp 1635330089
transform 1 0 6164 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1635330089
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1635330089
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_18
timestamp 1635330089
transform 1 0 2760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_6
timestamp 1635330089
transform 1 0 1656 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635330089
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635330089
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_30
timestamp 1635330089
transform 1 0 3864 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_42
timestamp 1635330089
transform 1 0 4968 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_48
timestamp 1635330089
transform 1 0 5520 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1635330089
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1635330089
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635330089
transform -1 0 6808 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1635330089
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635330089
transform 1 0 5612 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1635330089
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1635330089
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635330089
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1635330089
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635330089
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_41
timestamp 1635330089
transform 1 0 4876 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1635330089
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_47
timestamp 1635330089
transform 1 0 5428 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_51
timestamp 1635330089
transform 1 0 5796 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_55
timestamp 1635330089
transform 1 0 6164 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635330089
transform -1 0 6808 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _094_
timestamp 1635330089
transform 1 0 5060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1635330089
transform 1 0 5888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_18
timestamp 1635330089
transform 1 0 2760 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_6
timestamp 1635330089
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635330089
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635330089
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_30
timestamp 1635330089
transform 1 0 3864 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_36
timestamp 1635330089
transform 1 0 4416 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_41
timestamp 1635330089
transform 1 0 4876 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _092_
timestamp 1635330089
transform 1 0 4508 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_49
timestamp 1635330089
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1635330089
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1635330089
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635330089
transform -1 0 6808 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1635330089
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _093_
timestamp 1635330089
transform 1 0 5244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_18
timestamp 1635330089
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_6
timestamp 1635330089
transform 1 0 1656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635330089
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635330089
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1635330089
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1635330089
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_41
timestamp 1635330089
transform 1 0 4876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1635330089
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_48
timestamp 1635330089
transform 1 0 5520 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_55
timestamp 1635330089
transform 1 0 6164 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635330089
transform -1 0 6808 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1635330089
transform 1 0 5888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1635330089
transform 1 0 5244 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_18
timestamp 1635330089
transform 1 0 2760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_6
timestamp 1635330089
transform 1 0 1656 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635330089
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635330089
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_25
timestamp 1635330089
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_37
timestamp 1635330089
transform 1 0 4508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _048_
timestamp 1635330089
transform 1 0 3036 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1635330089
transform 1 0 4876 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_44
timestamp 1635330089
transform 1 0 5152 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1635330089
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1635330089
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635330089
transform -1 0 6808 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1635330089
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _095_
timestamp 1635330089
transform 1 0 5520 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _096_
timestamp 1635330089
transform 1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1635330089
transform 1 0 1564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635330089
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635330089
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_8
timestamp 1635330089
transform 1 0 1840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1635330089
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1635330089
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635330089
transform 1 0 2208 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1635330089
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_11
timestamp 1635330089
transform 1 0 2116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1635330089
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1635330089
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1635330089
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_37
timestamp 1635330089
transform 1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1635330089
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_39
timestamp 1635330089
transform 1 0 4692 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1635330089
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1635330089
transform 1 0 4140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1635330089
transform 1 0 5612 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _017_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 5520 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_47_47
timestamp 1635330089
transform 1 0 5428 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_45
timestamp 1635330089
transform 1 0 5244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1635330089
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1635330089
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1635330089
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_55
timestamp 1635330089
transform 1 0 6164 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635330089
transform -1 0 6808 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635330089
transform -1 0 6808 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_10
timestamp 1635330089
transform 1 0 2024 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1635330089
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635330089
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1635330089
transform 1 0 1748 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_22
timestamp 1635330089
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1635330089
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_41
timestamp 1635330089
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1635330089
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_46
timestamp 1635330089
transform 1 0 5336 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_55
timestamp 1635330089
transform 1 0 6164 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635330089
transform -1 0 6808 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1635330089
transform 1 0 4968 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1635330089
transform 1 0 5888 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_14
timestamp 1635330089
transform 1 0 2392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_6
timestamp 1635330089
transform 1 0 1656 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635330089
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1635330089
transform 1 0 2024 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1635330089
transform 1 0 2760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635330089
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_22
timestamp 1635330089
transform 1 0 3128 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_34
timestamp 1635330089
transform 1 0 4232 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1635330089
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1635330089
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635330089
transform -1 0 6808 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1635330089
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 4968 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_50_14
timestamp 1635330089
transform 1 0 2392 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1635330089
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_6
timestamp 1635330089
transform 1 0 1656 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635330089
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1635330089
transform 1 0 2576 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635330089
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1635330089
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_41
timestamp 1635330089
transform 1 0 4876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1635330089
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_55
timestamp 1635330089
transform 1 0 6164 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635330089
transform -1 0 6808 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input98
timestamp 1635330089
transform 1 0 5244 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_51_11
timestamp 1635330089
transform 1 0 2116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_18
timestamp 1635330089
transform 1 0 2760 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1635330089
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635330089
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1635330089
transform 1 0 2484 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1635330089
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1635330089
transform 1 0 3864 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_42
timestamp 1635330089
transform 1 0 4968 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1635330089
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1635330089
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1635330089
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635330089
transform -1 0 6808 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1635330089
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _100_
timestamp 1635330089
transform 1 0 5244 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_13
timestamp 1635330089
transform 1 0 2300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1635330089
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1635330089
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635330089
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635330089
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1635330089
transform 1 0 1380 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_52_25
timestamp 1635330089
transform 1 0 3404 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1635330089
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_41
timestamp 1635330089
transform 1 0 4876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_27
timestamp 1635330089
transform 1 0 3588 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_35
timestamp 1635330089
transform 1 0 4324 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_41
timestamp 1635330089
transform 1 0 4876 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1635330089
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _054_
timestamp 1635330089
transform 1 0 4508 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1635330089
transform 1 0 5244 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1635330089
transform 1 0 5612 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_48
timestamp 1635330089
transform 1 0 5520 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1635330089
transform 1 0 5888 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1635330089
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1635330089
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_55
timestamp 1635330089
transform 1 0 6164 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635330089
transform -1 0 6808 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635330089
transform -1 0 6808 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1635330089
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_11
timestamp 1635330089
transform 1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_18
timestamp 1635330089
transform 1 0 2760 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1635330089
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635330089
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1635330089
transform 1 0 2484 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1635330089
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1635330089
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1635330089
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_41
timestamp 1635330089
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1635330089
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_49
timestamp 1635330089
transform 1 0 5612 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_55
timestamp 1635330089
transform 1 0 6164 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635330089
transform -1 0 6808 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1635330089
transform 1 0 5888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_11
timestamp 1635330089
transform 1 0 2116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1635330089
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635330089
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1635330089
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_23
timestamp 1635330089
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_35
timestamp 1635330089
transform 1 0 4324 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_41
timestamp 1635330089
transform 1 0 4876 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1635330089
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1635330089
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635330089
transform -1 0 6808 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1635330089
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1635330089
transform 1 0 4968 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1635330089
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1635330089
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635330089
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1635330089
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1635330089
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_41
timestamp 1635330089
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1635330089
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_55
timestamp 1635330089
transform 1 0 6164 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635330089
transform -1 0 6808 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1635330089
transform 1 0 5244 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_57_11
timestamp 1635330089
transform 1 0 2116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1635330089
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635330089
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1635330089
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_23
timestamp 1635330089
transform 1 0 3220 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_35
timestamp 1635330089
transform 1 0 4324 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_41
timestamp 1635330089
transform 1 0 4876 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1635330089
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1635330089
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635330089
transform -1 0 6808 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1635330089
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1635330089
transform 1 0 4968 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_58_11
timestamp 1635330089
transform 1 0 2116 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_19
timestamp 1635330089
transform 1 0 2852 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_3
timestamp 1635330089
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635330089
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1635330089
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1635330089
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1635330089
transform 1 0 4048 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1635330089
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1635330089
transform 1 0 3036 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp 1635330089
transform 1 0 3772 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_44
timestamp 1635330089
transform 1 0 5152 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_55
timestamp 1635330089
transform 1 0 6164 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635330089
transform -1 0 6808 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1635330089
transform 1 0 5244 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_59_11
timestamp 1635330089
transform 1 0 2116 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_18
timestamp 1635330089
transform 1 0 2760 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1635330089
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1635330089
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1635330089
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635330089
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635330089
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1635330089
transform 1 0 2484 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1635330089
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1635330089
transform 1 0 3864 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1635330089
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1635330089
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_41
timestamp 1635330089
transform 1 0 4876 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1635330089
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1635330089
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1635330089
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_55
timestamp 1635330089
transform 1 0 6164 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635330089
transform -1 0 6808 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635330089
transform -1 0 6808 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1635330089
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1635330089
transform 1 0 4968 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1635330089
transform 1 0 5244 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_61_11
timestamp 1635330089
transform 1 0 2116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1635330089
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635330089
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1635330089
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_23
timestamp 1635330089
transform 1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_38
timestamp 1635330089
transform 1 0 4600 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1635330089
transform 1 0 4324 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1635330089
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1635330089
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635330089
transform -1 0 6808 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1635330089
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1635330089
transform 1 0 4968 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1635330089
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1635330089
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635330089
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1635330089
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1635330089
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1635330089
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_41
timestamp 1635330089
transform 1 0 4876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1635330089
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_55
timestamp 1635330089
transform 1 0 6164 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635330089
transform -1 0 6808 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1635330089
transform 1 0 5244 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_63_19
timestamp 1635330089
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_7
timestamp 1635330089
transform 1 0 1748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635330089
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1635330089
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_31
timestamp 1635330089
transform 1 0 3956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_39
timestamp 1635330089
transform 1 0 4692 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1635330089
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1635330089
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635330089
transform -1 0 6808 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1635330089
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1635330089
transform 1 0 4968 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1635330089
transform 1 0 2116 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1635330089
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1635330089
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635330089
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1635330089
transform 1 0 1840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1635330089
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1635330089
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1635330089
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1635330089
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1635330089
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_55
timestamp 1635330089
transform 1 0 6164 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635330089
transform -1 0 6808 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1635330089
transform 1 0 5244 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_65_19
timestamp 1635330089
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_7
timestamp 1635330089
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635330089
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1635330089
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_31
timestamp 1635330089
transform 1 0 3956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_39
timestamp 1635330089
transform 1 0 4692 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_52
timestamp 1635330089
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1635330089
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635330089
transform -1 0 6808 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1635330089
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1635330089
transform 1 0 4968 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1635330089
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_7
timestamp 1635330089
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1635330089
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1635330089
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635330089
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635330089
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1635330089
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1635330089
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_29
timestamp 1635330089
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_37
timestamp 1635330089
transform 1 0 4508 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_27
timestamp 1635330089
transform 1 0 3588 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_34
timestamp 1635330089
transform 1 0 4232 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1635330089
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _067_
timestamp 1635330089
transform 1 0 4140 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _068_
timestamp 1635330089
transform 1 0 3864 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_46
timestamp 1635330089
transform 1 0 5336 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1635330089
transform 1 0 5612 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_49
timestamp 1635330089
transform 1 0 5612 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1635330089
transform 1 0 5888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1635330089
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 1635330089
transform 1 0 5888 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_55
timestamp 1635330089
transform 1 0 6164 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635330089
transform -1 0 6808 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635330089
transform -1 0 6808 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 1635330089
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_19
timestamp 1635330089
transform 1 0 2852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_7
timestamp 1635330089
transform 1 0 1748 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635330089
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1635330089
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1635330089
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1635330089
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_41
timestamp 1635330089
transform 1 0 4876 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1635330089
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_49
timestamp 1635330089
transform 1 0 5612 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_55
timestamp 1635330089
transform 1 0 6164 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635330089
transform -1 0 6808 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1635330089
transform 1 0 5888 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_11
timestamp 1635330089
transform 1 0 2116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1635330089
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635330089
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _069_
timestamp 1635330089
transform 1 0 1748 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_23
timestamp 1635330089
transform 1 0 3220 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_35
timestamp 1635330089
transform 1 0 4324 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_47
timestamp 1635330089
transform 1 0 5428 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1635330089
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_57
timestamp 1635330089
transform 1 0 6348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635330089
transform -1 0 6808 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1635330089
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1635330089
transform 1 0 5612 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1635330089
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1635330089
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635330089
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1635330089
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1635330089
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1635330089
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_41
timestamp 1635330089
transform 1 0 4876 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1635330089
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_55
timestamp 1635330089
transform 1 0 6164 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635330089
transform -1 0 6808 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1635330089
transform 1 0 5244 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_71_19
timestamp 1635330089
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_7
timestamp 1635330089
transform 1 0 1748 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635330089
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1635330089
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_31
timestamp 1635330089
transform 1 0 3956 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_39
timestamp 1635330089
transform 1 0 4692 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_52
timestamp 1635330089
transform 1 0 5888 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_57
timestamp 1635330089
transform 1 0 6348 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635330089
transform -1 0 6808 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1635330089
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1635330089
transform 1 0 4968 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_72_19
timestamp 1635330089
transform 1 0 2852 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_7
timestamp 1635330089
transform 1 0 1748 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_14
timestamp 1635330089
transform 1 0 2392 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_7
timestamp 1635330089
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635330089
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635330089
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp 1635330089
transform 1 0 2116 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1635330089
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1635330089
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1635330089
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_29
timestamp 1635330089
transform 1 0 3772 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_37
timestamp 1635330089
transform 1 0 4508 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_26
timestamp 1635330089
transform 1 0 3496 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_38
timestamp 1635330089
transform 1 0 4600 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1635330089
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp 1635330089
transform 1 0 3036 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _070_
timestamp 1635330089
transform 1 0 4140 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635330089
transform 1 0 5336 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_55
timestamp 1635330089
transform 1 0 6164 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_52
timestamp 1635330089
transform 1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_57
timestamp 1635330089
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635330089
transform -1 0 6808 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635330089
transform -1 0 6808 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1635330089
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input91
timestamp 1635330089
transform 1 0 5244 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1635330089
transform 1 0 5520 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1635330089
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1635330089
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635330089
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1635330089
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1635330089
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1635330089
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635330089
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_53
timestamp 1635330089
transform 1 0 5980 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635330089
transform -1 0 6808 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_19
timestamp 1635330089
transform 1 0 2852 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_7
timestamp 1635330089
transform 1 0 1748 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635330089
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1635330089
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_31
timestamp 1635330089
transform 1 0 3956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_43
timestamp 1635330089
transform 1 0 5060 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_47
timestamp 1635330089
transform 1 0 5428 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_52
timestamp 1635330089
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_57
timestamp 1635330089
transform 1 0 6348 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635330089
transform -1 0 6808 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635330089
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1635330089
transform 1 0 5520 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_19
timestamp 1635330089
transform 1 0 2852 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_7
timestamp 1635330089
transform 1 0 1748 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635330089
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1635330089
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1635330089
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1635330089
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_41
timestamp 1635330089
transform 1 0 4876 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635330089
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_49
timestamp 1635330089
transform 1 0 5612 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_55
timestamp 1635330089
transform 1 0 6164 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635330089
transform -1 0 6808 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1635330089
transform 1 0 5796 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_19
timestamp 1635330089
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_7
timestamp 1635330089
transform 1 0 1748 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635330089
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1635330089
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_31
timestamp 1635330089
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_43
timestamp 1635330089
transform 1 0 5060 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_47
timestamp 1635330089
transform 1 0 5428 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_52
timestamp 1635330089
transform 1 0 5888 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1635330089
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635330089
transform -1 0 6808 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635330089
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1635330089
transform 1 0 5520 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_11
timestamp 1635330089
transform 1 0 2116 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_16
timestamp 1635330089
transform 1 0 2576 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1635330089
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635330089
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1635330089
transform 1 0 2300 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1635330089
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_41
timestamp 1635330089
transform 1 0 4876 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635330089
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_49
timestamp 1635330089
transform 1 0 5612 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_55
timestamp 1635330089
transform 1 0 6164 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635330089
transform -1 0 6808 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1635330089
transform 1 0 5796 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_19
timestamp 1635330089
transform 1 0 2852 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_7
timestamp 1635330089
transform 1 0 1748 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_19
timestamp 1635330089
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_7
timestamp 1635330089
transform 1 0 1748 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635330089
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1635330089
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1635330089
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1635330089
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_31
timestamp 1635330089
transform 1 0 3956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1635330089
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1635330089
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_41
timestamp 1635330089
transform 1 0 4876 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635330089
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_43
timestamp 1635330089
transform 1 0 5060 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1635330089
transform 1 0 5336 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1635330089
transform 1 0 5796 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1635330089
transform 1 0 5520 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_49
timestamp 1635330089
transform 1 0 5612 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635330089
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_55
timestamp 1635330089
transform 1 0 6164 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1635330089
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1635330089
transform -1 0 6808 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635330089
transform -1 0 6808 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_57
timestamp 1635330089
transform 1 0 6348 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_15
timestamp 1635330089
transform 1 0 2484 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1635330089
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1635330089
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1635330089
transform 1 0 2760 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_21
timestamp 1635330089
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_36
timestamp 1635330089
transform 1 0 4416 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1635330089
transform 1 0 4140 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1635330089
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_57
timestamp 1635330089
transform 1 0 6348 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1635330089
transform -1 0 6808 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635330089
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1635330089
transform 1 0 5520 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_19
timestamp 1635330089
transform 1 0 2852 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_7
timestamp 1635330089
transform 1 0 1748 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1635330089
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1635330089
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1635330089
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1635330089
transform 1 0 4048 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635330089
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1635330089
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1635330089
transform 1 0 5612 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_44
timestamp 1635330089
transform 1 0 5152 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_48
timestamp 1635330089
transform 1 0 5520 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_55
timestamp 1635330089
transform 1 0 6164 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1635330089
transform -1 0 6808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1635330089
transform 1 0 5796 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_19
timestamp 1635330089
transform 1 0 2852 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_7
timestamp 1635330089
transform 1 0 1748 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1635330089
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1635330089
transform 1 0 1380 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_31
timestamp 1635330089
transform 1 0 3956 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1635330089
transform 1 0 5336 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_83_43
timestamp 1635330089
transform 1 0 5060 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_52
timestamp 1635330089
transform 1 0 5888 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_57
timestamp 1635330089
transform 1 0 6348 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1635330089
transform -1 0 6808 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635330089
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1635330089
transform 1 0 5520 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_19
timestamp 1635330089
transform 1 0 2852 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_7
timestamp 1635330089
transform 1 0 1748 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1635330089
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1635330089
transform 1 0 1380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_24
timestamp 1635330089
transform 1 0 3312 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_32
timestamp 1635330089
transform 1 0 4048 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635330089
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1635330089
transform 1 0 3772 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1635330089
transform 1 0 3036 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_84_44
timestamp 1635330089
transform 1 0 5152 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_50
timestamp 1635330089
transform 1 0 5704 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_55
timestamp 1635330089
transform 1 0 6164 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1635330089
transform -1 0 6808 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1635330089
transform 1 0 5796 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1635330089
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1635330089
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_19
timestamp 1635330089
transform 1 0 2852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_7
timestamp 1635330089
transform 1 0 1748 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1635330089
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1635330089
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1635330089
transform 1 0 1380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1635330089
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_39
timestamp 1635330089
transform 1 0 4692 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1635330089
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1635330089
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_41
timestamp 1635330089
transform 1 0 4876 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635330089
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_45
timestamp 1635330089
transform 1 0 5244 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1635330089
transform 1 0 5336 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1635330089
transform 1 0 5796 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1635330089
transform 1 0 5520 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_49
timestamp 1635330089
transform 1 0 5612 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635330089
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_55
timestamp 1635330089
transform 1 0 6164 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_52
timestamp 1635330089
transform 1 0 5888 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1635330089
transform -1 0 6808 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1635330089
transform -1 0 6808 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_57
timestamp 1635330089
transform 1 0 6348 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_14
timestamp 1635330089
transform 1 0 2392 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_7
timestamp 1635330089
transform 1 0 1748 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1635330089
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1635330089
transform 1 0 2116 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1635330089
transform 1 0 1380 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_26
timestamp 1635330089
transform 1 0 3496 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_38
timestamp 1635330089
transform 1 0 4600 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1635330089
transform 1 0 5336 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_52
timestamp 1635330089
transform 1 0 5888 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_57
timestamp 1635330089
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1635330089
transform -1 0 6808 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635330089
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1635330089
transform 1 0 5520 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_20
timestamp 1635330089
transform 1 0 2944 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1635330089
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_8
timestamp 1635330089
transform 1 0 1840 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1635330089
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1635330089
transform 1 0 1564 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1635330089
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_41
timestamp 1635330089
transform 1 0 4876 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635330089
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_49
timestamp 1635330089
transform 1 0 5612 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_55
timestamp 1635330089
transform 1 0 6164 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1635330089
transform -1 0 6808 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1635330089
transform 1 0 5796 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_14
timestamp 1635330089
transform 1 0 2392 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_7
timestamp 1635330089
transform 1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1635330089
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1635330089
transform 1 0 2116 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1635330089
transform 1 0 2760 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1635330089
transform 1 0 1380 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_21
timestamp 1635330089
transform 1 0 3036 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_33
timestamp 1635330089
transform 1 0 4140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_89_45
timestamp 1635330089
transform 1 0 5244 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_52
timestamp 1635330089
transform 1 0 5888 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_57
timestamp 1635330089
transform 1 0 6348 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1635330089
transform -1 0 6808 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635330089
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1635330089
transform 1 0 5520 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_19
timestamp 1635330089
transform 1 0 2852 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_7
timestamp 1635330089
transform 1 0 1748 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1635330089
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1635330089
transform 1 0 1380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1635330089
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1635330089
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_41
timestamp 1635330089
transform 1 0 4876 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635330089
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1635330089
transform 1 0 5612 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_55
timestamp 1635330089
transform 1 0 6164 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1635330089
transform -1 0 6808 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1635330089
transform 1 0 5796 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_19
timestamp 1635330089
transform 1 0 2852 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_91_7
timestamp 1635330089
transform 1 0 1748 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1635330089
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1635330089
transform 1 0 1380 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_25
timestamp 1635330089
transform 1 0 3404 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_29
timestamp 1635330089
transform 1 0 3772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_41
timestamp 1635330089
transform 1 0 4876 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1635330089
transform 1 0 3496 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_91_47
timestamp 1635330089
transform 1 0 5428 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_52
timestamp 1635330089
transform 1 0 5888 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_57
timestamp 1635330089
transform 1 0 6348 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1635330089
transform -1 0 6808 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635330089
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1635330089
transform 1 0 5520 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_15
timestamp 1635330089
transform 1 0 2484 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1635330089
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_19
timestamp 1635330089
transform 1 0 2852 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_7
timestamp 1635330089
transform 1 0 1748 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1635330089
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1635330089
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1635330089
transform 1 0 1380 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_24
timestamp 1635330089
transform 1 0 3312 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1635330089
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_41
timestamp 1635330089
transform 1 0 4876 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_28
timestamp 1635330089
transform 1 0 3680 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_40
timestamp 1635330089
transform 1 0 4784 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635330089
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1635330089
transform 1 0 3404 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1635330089
transform 1 0 3036 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1635330089
transform 1 0 5336 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1635330089
transform 1 0 5520 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1635330089
transform 1 0 5796 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_49
timestamp 1635330089
transform 1 0 5612 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635330089
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_52
timestamp 1635330089
transform 1 0 5888 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_55
timestamp 1635330089
transform 1 0 6164 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1635330089
transform -1 0 6808 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1635330089
transform -1 0 6808 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1635330089
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_19
timestamp 1635330089
transform 1 0 2852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_7
timestamp 1635330089
transform 1 0 1748 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1635330089
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1635330089
transform 1 0 1380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1635330089
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1635330089
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_41
timestamp 1635330089
transform 1 0 4876 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635330089
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1635330089
transform 1 0 5612 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_55
timestamp 1635330089
transform 1 0 6164 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1635330089
transform -1 0 6808 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1635330089
transform 1 0 5796 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_15
timestamp 1635330089
transform 1 0 2484 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1635330089
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1635330089
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_26
timestamp 1635330089
transform 1 0 3496 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_38
timestamp 1635330089
transform 1 0 4600 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1635330089
transform 1 0 3220 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1635330089
transform 1 0 4876 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_44
timestamp 1635330089
transform 1 0 5152 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_52
timestamp 1635330089
transform 1 0 5888 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_57
timestamp 1635330089
transform 1 0 6348 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1635330089
transform -1 0 6808 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635330089
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1635330089
transform 1 0 5520 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_14
timestamp 1635330089
transform 1 0 2392 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_7
timestamp 1635330089
transform 1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1635330089
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1635330089
transform 1 0 2116 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1635330089
transform 1 0 1380 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_26
timestamp 1635330089
transform 1 0 3496 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_32
timestamp 1635330089
transform 1 0 4048 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635330089
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1635330089
transform 1 0 3772 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_96_44
timestamp 1635330089
transform 1 0 5152 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_50
timestamp 1635330089
transform 1 0 5704 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_55
timestamp 1635330089
transform 1 0 6164 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1635330089
transform -1 0 6808 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1635330089
transform 1 0 5796 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_14
timestamp 1635330089
transform 1 0 2392 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_97_7
timestamp 1635330089
transform 1 0 1748 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1635330089
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1635330089
transform 1 0 2944 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1635330089
transform 1 0 2116 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1635330089
transform 1 0 1380 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_23
timestamp 1635330089
transform 1 0 3220 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_31
timestamp 1635330089
transform 1 0 3956 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_35
timestamp 1635330089
transform 1 0 4324 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1635330089
transform 1 0 4692 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1635330089
transform 1 0 4048 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1635330089
transform 1 0 5336 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_42
timestamp 1635330089
transform 1 0 4968 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_52
timestamp 1635330089
transform 1 0 5888 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_57
timestamp 1635330089
transform 1 0 6348 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1635330089
transform -1 0 6808 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635330089
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1635330089
transform 1 0 5520 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_19
timestamp 1635330089
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_7
timestamp 1635330089
transform 1 0 1748 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1635330089
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1635330089
transform 1 0 1380 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1635330089
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_29
timestamp 1635330089
transform 1 0 3772 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_33
timestamp 1635330089
transform 1 0 4140 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_37
timestamp 1635330089
transform 1 0 4508 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635330089
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1635330089
transform 1 0 4232 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_49
timestamp 1635330089
transform 1 0 5612 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_55
timestamp 1635330089
transform 1 0 6164 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1635330089
transform -1 0 6808 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1635330089
transform 1 0 5796 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_19
timestamp 1635330089
transform 1 0 2852 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_7
timestamp 1635330089
transform 1 0 1748 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_19
timestamp 1635330089
transform 1 0 2852 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_7
timestamp 1635330089
transform 1 0 1748 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1635330089
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1635330089
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1635330089
transform 1 0 1380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1635330089
transform 1 0 1380 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1635330089
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_29
timestamp 1635330089
transform 1 0 3772 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_39
timestamp 1635330089
transform 1 0 4692 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_31
timestamp 1635330089
transform 1 0 3956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635330089
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1635330089
transform 1 0 4324 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1635330089
transform 1 0 5060 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_43
timestamp 1635330089
transform 1 0 5060 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1635330089
transform 1 0 5796 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1635330089
transform 1 0 5520 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_47
timestamp 1635330089
transform 1 0 5428 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_47
timestamp 1635330089
transform 1 0 5428 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635330089
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_52
timestamp 1635330089
transform 1 0 5888 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_55
timestamp 1635330089
transform 1 0 6164 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1635330089
transform -1 0 6808 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1635330089
transform -1 0 6808 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_57
timestamp 1635330089
transform 1 0 6348 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_15
timestamp 1635330089
transform 1 0 2484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_7
timestamp 1635330089
transform 1 0 1748 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1635330089
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1635330089
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1635330089
transform 1 0 2116 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1635330089
transform 1 0 2852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_23
timestamp 1635330089
transform 1 0 3220 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1635330089
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_29
timestamp 1635330089
transform 1 0 3772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_36
timestamp 1635330089
transform 1 0 4416 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635330089
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1635330089
transform 1 0 4784 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1635330089
transform 1 0 4048 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_44
timestamp 1635330089
transform 1 0 5152 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_52
timestamp 1635330089
transform 1 0 5888 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1635330089
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1635330089
transform -1 0 6808 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635330089
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1635330089
transform 1 0 5520 0 -1 57664
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 5584 800 5704 6 ram_addr0[0]
port 0 nsew signal tristate
rlabel metal3 s 0 6264 800 6384 6 ram_addr0[1]
port 1 nsew signal tristate
rlabel metal3 s 0 7080 800 7200 6 ram_addr0[2]
port 2 nsew signal tristate
rlabel metal3 s 0 7760 800 7880 6 ram_addr0[3]
port 3 nsew signal tristate
rlabel metal3 s 0 8576 800 8696 6 ram_addr0[4]
port 4 nsew signal tristate
rlabel metal3 s 0 9256 800 9376 6 ram_addr0[5]
port 5 nsew signal tristate
rlabel metal3 s 0 10072 800 10192 6 ram_addr0[6]
port 6 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 ram_addr0[7]
port 7 nsew signal tristate
rlabel metal3 s 0 280 800 400 6 ram_clk0
port 8 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 ram_csb0
port 9 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 ram_din0[0]
port 10 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 ram_din0[10]
port 11 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 ram_din0[11]
port 12 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 ram_din0[12]
port 13 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 ram_din0[13]
port 14 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 ram_din0[14]
port 15 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 ram_din0[15]
port 16 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 ram_din0[16]
port 17 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 ram_din0[17]
port 18 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 ram_din0[18]
port 19 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 ram_din0[19]
port 20 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 ram_din0[1]
port 21 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 ram_din0[20]
port 22 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 ram_din0[21]
port 23 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 ram_din0[22]
port 24 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 ram_din0[23]
port 25 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 ram_din0[24]
port 26 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 ram_din0[25]
port 27 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 ram_din0[26]
port 28 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 ram_din0[27]
port 29 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 ram_din0[28]
port 30 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 ram_din0[29]
port 31 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 ram_din0[2]
port 32 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 ram_din0[30]
port 33 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 ram_din0[31]
port 34 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 ram_din0[3]
port 35 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 ram_din0[4]
port 36 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 ram_din0[5]
port 37 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 ram_din0[6]
port 38 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 ram_din0[7]
port 39 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 ram_din0[8]
port 40 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 ram_din0[9]
port 41 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 ram_dout0[0]
port 42 nsew signal tristate
rlabel metal3 s 0 43528 800 43648 6 ram_dout0[10]
port 43 nsew signal tristate
rlabel metal3 s 0 44208 800 44328 6 ram_dout0[11]
port 44 nsew signal tristate
rlabel metal3 s 0 45024 800 45144 6 ram_dout0[12]
port 45 nsew signal tristate
rlabel metal3 s 0 45704 800 45824 6 ram_dout0[13]
port 46 nsew signal tristate
rlabel metal3 s 0 46520 800 46640 6 ram_dout0[14]
port 47 nsew signal tristate
rlabel metal3 s 0 47336 800 47456 6 ram_dout0[15]
port 48 nsew signal tristate
rlabel metal3 s 0 48016 800 48136 6 ram_dout0[16]
port 49 nsew signal tristate
rlabel metal3 s 0 48832 800 48952 6 ram_dout0[17]
port 50 nsew signal tristate
rlabel metal3 s 0 49512 800 49632 6 ram_dout0[18]
port 51 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 ram_dout0[19]
port 52 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 ram_dout0[1]
port 53 nsew signal tristate
rlabel metal3 s 0 51144 800 51264 6 ram_dout0[20]
port 54 nsew signal tristate
rlabel metal3 s 0 51824 800 51944 6 ram_dout0[21]
port 55 nsew signal tristate
rlabel metal3 s 0 52640 800 52760 6 ram_dout0[22]
port 56 nsew signal tristate
rlabel metal3 s 0 53320 800 53440 6 ram_dout0[23]
port 57 nsew signal tristate
rlabel metal3 s 0 54136 800 54256 6 ram_dout0[24]
port 58 nsew signal tristate
rlabel metal3 s 0 54816 800 54936 6 ram_dout0[25]
port 59 nsew signal tristate
rlabel metal3 s 0 55632 800 55752 6 ram_dout0[26]
port 60 nsew signal tristate
rlabel metal3 s 0 56448 800 56568 6 ram_dout0[27]
port 61 nsew signal tristate
rlabel metal3 s 0 57128 800 57248 6 ram_dout0[28]
port 62 nsew signal tristate
rlabel metal3 s 0 57944 800 58064 6 ram_dout0[29]
port 63 nsew signal tristate
rlabel metal3 s 0 37408 800 37528 6 ram_dout0[2]
port 64 nsew signal tristate
rlabel metal3 s 0 58624 800 58744 6 ram_dout0[30]
port 65 nsew signal tristate
rlabel metal3 s 0 59440 800 59560 6 ram_dout0[31]
port 66 nsew signal tristate
rlabel metal3 s 0 38224 800 38344 6 ram_dout0[3]
port 67 nsew signal tristate
rlabel metal3 s 0 38904 800 39024 6 ram_dout0[4]
port 68 nsew signal tristate
rlabel metal3 s 0 39720 800 39840 6 ram_dout0[5]
port 69 nsew signal tristate
rlabel metal3 s 0 40400 800 40520 6 ram_dout0[6]
port 70 nsew signal tristate
rlabel metal3 s 0 41216 800 41336 6 ram_dout0[7]
port 71 nsew signal tristate
rlabel metal3 s 0 42032 800 42152 6 ram_dout0[8]
port 72 nsew signal tristate
rlabel metal3 s 0 42712 800 42832 6 ram_dout0[9]
port 73 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 ram_web0
port 74 nsew signal tristate
rlabel metal3 s 0 2456 800 2576 6 ram_wmask0[0]
port 75 nsew signal tristate
rlabel metal3 s 0 3272 800 3392 6 ram_wmask0[1]
port 76 nsew signal tristate
rlabel metal3 s 0 3952 800 4072 6 ram_wmask0[2]
port 77 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 ram_wmask0[3]
port 78 nsew signal tristate
rlabel metal4 s 1909 2128 2229 57712 6 vccd1
port 79 nsew power input
rlabel metal4 s 3839 2128 4159 57712 6 vccd1
port 79 nsew power input
rlabel metal4 s 5770 2128 6090 57712 6 vccd1
port 79 nsew power input
rlabel metal4 s 2874 2128 3194 57712 6 vssd1
port 80 nsew ground input
rlabel metal4 s 4805 2128 5125 57712 6 vssd1
port 80 nsew ground input
rlabel metal3 s 7200 280 8000 400 6 wb_clk_i
port 81 nsew signal input
rlabel metal3 s 7200 824 8000 944 6 wb_rst_i
port 82 nsew signal input
rlabel metal3 s 7200 3000 8000 3120 6 wbs_ack_o
port 83 nsew signal tristate
rlabel metal3 s 7200 5856 8000 5976 6 wbs_adr_i[0]
port 84 nsew signal input
rlabel metal3 s 7200 11568 8000 11688 6 wbs_adr_i[10]
port 85 nsew signal input
rlabel metal3 s 7200 12112 8000 12232 6 wbs_adr_i[11]
port 86 nsew signal input
rlabel metal3 s 7200 12656 8000 12776 6 wbs_adr_i[12]
port 87 nsew signal input
rlabel metal3 s 7200 13200 8000 13320 6 wbs_adr_i[13]
port 88 nsew signal input
rlabel metal3 s 7200 13744 8000 13864 6 wbs_adr_i[14]
port 89 nsew signal input
rlabel metal3 s 7200 14424 8000 14544 6 wbs_adr_i[15]
port 90 nsew signal input
rlabel metal3 s 7200 14968 8000 15088 6 wbs_adr_i[16]
port 91 nsew signal input
rlabel metal3 s 7200 15512 8000 15632 6 wbs_adr_i[17]
port 92 nsew signal input
rlabel metal3 s 7200 16056 8000 16176 6 wbs_adr_i[18]
port 93 nsew signal input
rlabel metal3 s 7200 16600 8000 16720 6 wbs_adr_i[19]
port 94 nsew signal input
rlabel metal3 s 7200 6400 8000 6520 6 wbs_adr_i[1]
port 95 nsew signal input
rlabel metal3 s 7200 17144 8000 17264 6 wbs_adr_i[20]
port 96 nsew signal input
rlabel metal3 s 7200 17688 8000 17808 6 wbs_adr_i[21]
port 97 nsew signal input
rlabel metal3 s 7200 18368 8000 18488 6 wbs_adr_i[22]
port 98 nsew signal input
rlabel metal3 s 7200 18912 8000 19032 6 wbs_adr_i[23]
port 99 nsew signal input
rlabel metal3 s 7200 19456 8000 19576 6 wbs_adr_i[24]
port 100 nsew signal input
rlabel metal3 s 7200 20000 8000 20120 6 wbs_adr_i[25]
port 101 nsew signal input
rlabel metal3 s 7200 20544 8000 20664 6 wbs_adr_i[26]
port 102 nsew signal input
rlabel metal3 s 7200 21088 8000 21208 6 wbs_adr_i[27]
port 103 nsew signal input
rlabel metal3 s 7200 21768 8000 21888 6 wbs_adr_i[28]
port 104 nsew signal input
rlabel metal3 s 7200 22312 8000 22432 6 wbs_adr_i[29]
port 105 nsew signal input
rlabel metal3 s 7200 6944 8000 7064 6 wbs_adr_i[2]
port 106 nsew signal input
rlabel metal3 s 7200 22856 8000 22976 6 wbs_adr_i[30]
port 107 nsew signal input
rlabel metal3 s 7200 23400 8000 23520 6 wbs_adr_i[31]
port 108 nsew signal input
rlabel metal3 s 7200 7624 8000 7744 6 wbs_adr_i[3]
port 109 nsew signal input
rlabel metal3 s 7200 8168 8000 8288 6 wbs_adr_i[4]
port 110 nsew signal input
rlabel metal3 s 7200 8712 8000 8832 6 wbs_adr_i[5]
port 111 nsew signal input
rlabel metal3 s 7200 9256 8000 9376 6 wbs_adr_i[6]
port 112 nsew signal input
rlabel metal3 s 7200 9800 8000 9920 6 wbs_adr_i[7]
port 113 nsew signal input
rlabel metal3 s 7200 10344 8000 10464 6 wbs_adr_i[8]
port 114 nsew signal input
rlabel metal3 s 7200 11024 8000 11144 6 wbs_adr_i[9]
port 115 nsew signal input
rlabel metal3 s 7200 1912 8000 2032 6 wbs_cyc_i
port 116 nsew signal input
rlabel metal3 s 7200 23944 8000 24064 6 wbs_dat_i[0]
port 117 nsew signal input
rlabel metal3 s 7200 29656 8000 29776 6 wbs_dat_i[10]
port 118 nsew signal input
rlabel metal3 s 7200 30200 8000 30320 6 wbs_dat_i[11]
port 119 nsew signal input
rlabel metal3 s 7200 30744 8000 30864 6 wbs_dat_i[12]
port 120 nsew signal input
rlabel metal3 s 7200 31288 8000 31408 6 wbs_dat_i[13]
port 121 nsew signal input
rlabel metal3 s 7200 31832 8000 31952 6 wbs_dat_i[14]
port 122 nsew signal input
rlabel metal3 s 7200 32512 8000 32632 6 wbs_dat_i[15]
port 123 nsew signal input
rlabel metal3 s 7200 33056 8000 33176 6 wbs_dat_i[16]
port 124 nsew signal input
rlabel metal3 s 7200 33600 8000 33720 6 wbs_dat_i[17]
port 125 nsew signal input
rlabel metal3 s 7200 34144 8000 34264 6 wbs_dat_i[18]
port 126 nsew signal input
rlabel metal3 s 7200 34688 8000 34808 6 wbs_dat_i[19]
port 127 nsew signal input
rlabel metal3 s 7200 24488 8000 24608 6 wbs_dat_i[1]
port 128 nsew signal input
rlabel metal3 s 7200 35232 8000 35352 6 wbs_dat_i[20]
port 129 nsew signal input
rlabel metal3 s 7200 35912 8000 36032 6 wbs_dat_i[21]
port 130 nsew signal input
rlabel metal3 s 7200 36456 8000 36576 6 wbs_dat_i[22]
port 131 nsew signal input
rlabel metal3 s 7200 37000 8000 37120 6 wbs_dat_i[23]
port 132 nsew signal input
rlabel metal3 s 7200 37544 8000 37664 6 wbs_dat_i[24]
port 133 nsew signal input
rlabel metal3 s 7200 38088 8000 38208 6 wbs_dat_i[25]
port 134 nsew signal input
rlabel metal3 s 7200 38632 8000 38752 6 wbs_dat_i[26]
port 135 nsew signal input
rlabel metal3 s 7200 39312 8000 39432 6 wbs_dat_i[27]
port 136 nsew signal input
rlabel metal3 s 7200 39856 8000 39976 6 wbs_dat_i[28]
port 137 nsew signal input
rlabel metal3 s 7200 40400 8000 40520 6 wbs_dat_i[29]
port 138 nsew signal input
rlabel metal3 s 7200 25168 8000 25288 6 wbs_dat_i[2]
port 139 nsew signal input
rlabel metal3 s 7200 40944 8000 41064 6 wbs_dat_i[30]
port 140 nsew signal input
rlabel metal3 s 7200 41488 8000 41608 6 wbs_dat_i[31]
port 141 nsew signal input
rlabel metal3 s 7200 25712 8000 25832 6 wbs_dat_i[3]
port 142 nsew signal input
rlabel metal3 s 7200 26256 8000 26376 6 wbs_dat_i[4]
port 143 nsew signal input
rlabel metal3 s 7200 26800 8000 26920 6 wbs_dat_i[5]
port 144 nsew signal input
rlabel metal3 s 7200 27344 8000 27464 6 wbs_dat_i[6]
port 145 nsew signal input
rlabel metal3 s 7200 27888 8000 28008 6 wbs_dat_i[7]
port 146 nsew signal input
rlabel metal3 s 7200 28568 8000 28688 6 wbs_dat_i[8]
port 147 nsew signal input
rlabel metal3 s 7200 29112 8000 29232 6 wbs_dat_i[9]
port 148 nsew signal input
rlabel metal3 s 7200 42032 8000 42152 6 wbs_dat_o[0]
port 149 nsew signal tristate
rlabel metal3 s 7200 47744 8000 47864 6 wbs_dat_o[10]
port 150 nsew signal tristate
rlabel metal3 s 7200 48288 8000 48408 6 wbs_dat_o[11]
port 151 nsew signal tristate
rlabel metal3 s 7200 48832 8000 48952 6 wbs_dat_o[12]
port 152 nsew signal tristate
rlabel metal3 s 7200 49376 8000 49496 6 wbs_dat_o[13]
port 153 nsew signal tristate
rlabel metal3 s 7200 50056 8000 50176 6 wbs_dat_o[14]
port 154 nsew signal tristate
rlabel metal3 s 7200 50600 8000 50720 6 wbs_dat_o[15]
port 155 nsew signal tristate
rlabel metal3 s 7200 51144 8000 51264 6 wbs_dat_o[16]
port 156 nsew signal tristate
rlabel metal3 s 7200 51688 8000 51808 6 wbs_dat_o[17]
port 157 nsew signal tristate
rlabel metal3 s 7200 52232 8000 52352 6 wbs_dat_o[18]
port 158 nsew signal tristate
rlabel metal3 s 7200 52776 8000 52896 6 wbs_dat_o[19]
port 159 nsew signal tristate
rlabel metal3 s 7200 42712 8000 42832 6 wbs_dat_o[1]
port 160 nsew signal tristate
rlabel metal3 s 7200 53456 8000 53576 6 wbs_dat_o[20]
port 161 nsew signal tristate
rlabel metal3 s 7200 54000 8000 54120 6 wbs_dat_o[21]
port 162 nsew signal tristate
rlabel metal3 s 7200 54544 8000 54664 6 wbs_dat_o[22]
port 163 nsew signal tristate
rlabel metal3 s 7200 55088 8000 55208 6 wbs_dat_o[23]
port 164 nsew signal tristate
rlabel metal3 s 7200 55632 8000 55752 6 wbs_dat_o[24]
port 165 nsew signal tristate
rlabel metal3 s 7200 56176 8000 56296 6 wbs_dat_o[25]
port 166 nsew signal tristate
rlabel metal3 s 7200 56856 8000 56976 6 wbs_dat_o[26]
port 167 nsew signal tristate
rlabel metal3 s 7200 57400 8000 57520 6 wbs_dat_o[27]
port 168 nsew signal tristate
rlabel metal3 s 7200 57944 8000 58064 6 wbs_dat_o[28]
port 169 nsew signal tristate
rlabel metal3 s 7200 58488 8000 58608 6 wbs_dat_o[29]
port 170 nsew signal tristate
rlabel metal3 s 7200 43256 8000 43376 6 wbs_dat_o[2]
port 171 nsew signal tristate
rlabel metal3 s 7200 59032 8000 59152 6 wbs_dat_o[30]
port 172 nsew signal tristate
rlabel metal3 s 7200 59576 8000 59696 6 wbs_dat_o[31]
port 173 nsew signal tristate
rlabel metal3 s 7200 43800 8000 43920 6 wbs_dat_o[3]
port 174 nsew signal tristate
rlabel metal3 s 7200 44344 8000 44464 6 wbs_dat_o[4]
port 175 nsew signal tristate
rlabel metal3 s 7200 44888 8000 45008 6 wbs_dat_o[5]
port 176 nsew signal tristate
rlabel metal3 s 7200 45432 8000 45552 6 wbs_dat_o[6]
port 177 nsew signal tristate
rlabel metal3 s 7200 45976 8000 46096 6 wbs_dat_o[7]
port 178 nsew signal tristate
rlabel metal3 s 7200 46656 8000 46776 6 wbs_dat_o[8]
port 179 nsew signal tristate
rlabel metal3 s 7200 47200 8000 47320 6 wbs_dat_o[9]
port 180 nsew signal tristate
rlabel metal3 s 7200 3544 8000 3664 6 wbs_sel_i[0]
port 181 nsew signal input
rlabel metal3 s 7200 4224 8000 4344 6 wbs_sel_i[1]
port 182 nsew signal input
rlabel metal3 s 7200 4768 8000 4888 6 wbs_sel_i[2]
port 183 nsew signal input
rlabel metal3 s 7200 5312 8000 5432 6 wbs_sel_i[3]
port 184 nsew signal input
rlabel metal3 s 7200 1368 8000 1488 6 wbs_stb_i
port 185 nsew signal input
rlabel metal3 s 7200 2456 8000 2576 6 wbs_we_i
port 186 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 8000 60000
<< end >>
